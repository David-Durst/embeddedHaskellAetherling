module FIFO(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  output [7:0] O_0,
  output [7:0] O_1
);
  reg [7:0] _T__0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg [7:0] _T__1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_1;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_2;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O_0 = _T__0; // @[FIFO.scala 14:7]
  assign O_1 = _T__1; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T__0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T__1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T__0 <= I_0;
    _T__1 <= I_1;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module NestedCounters(
  input   CE,
  output  valid
);
  assign valid = CE; // @[NestedCounters.scala 65:13]
endmodule
module NestedCounters_1(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 53:31]
  wire  NestedCounters_valid; // @[NestedCounters.scala 53:31]
  NestedCounters NestedCounters ( // @[NestedCounters.scala 53:31]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 56:11]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 57:22]
endmodule
module NestedCountersWithNumValid(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 20:44]
  wire  NestedCounters_valid; // @[NestedCounters.scala 20:44]
  NestedCounters_1 NestedCounters ( // @[NestedCounters.scala 20:44]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 22:9]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 21:27]
endmodule
module RAM_ST(
  input        clock,
  input        RE,
  input  [9:0] RADDR,
  output [7:0] RDATA_0,
  output [7:0] RDATA_1,
  input        WE,
  input  [9:0] WADDR,
  input  [7:0] WDATA_0,
  input  [7:0] WDATA_1
);
  wire  write_elem_counter_CE; // @[RAM_ST.scala 20:34]
  wire  write_elem_counter_valid; // @[RAM_ST.scala 20:34]
  wire  read_elem_counter_CE; // @[RAM_ST.scala 21:33]
  wire  read_elem_counter_valid; // @[RAM_ST.scala 21:33]
  reg [15:0] ram [0:959]; // @[RAM_ST.scala 29:24]
  reg [31:0] _RAND_0;
  wire [15:0] ram__T_9_data; // @[RAM_ST.scala 29:24]
  wire [9:0] ram__T_9_addr; // @[RAM_ST.scala 29:24]
  reg [31:0] _RAND_1;
  wire [15:0] ram__T_3_data; // @[RAM_ST.scala 29:24]
  wire [9:0] ram__T_3_addr; // @[RAM_ST.scala 29:24]
  wire  ram__T_3_mask; // @[RAM_ST.scala 29:24]
  wire  ram__T_3_en; // @[RAM_ST.scala 29:24]
  reg  ram__T_9_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [9:0] ram__T_9_addr_pipe_0;
  reg [31:0] _RAND_3;
  wire [9:0] _GEN_1; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_2; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_3; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_4; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_5; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_6; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_7; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_8; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_9; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_10; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_11; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_12; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_13; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_14; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_15; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_16; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_17; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_18; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_19; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_20; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_21; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_22; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_23; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_24; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_25; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_26; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_27; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_28; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_29; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_30; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_31; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_32; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_33; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_34; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_35; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_36; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_37; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_38; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_39; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_40; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_41; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_42; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_43; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_44; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_45; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_46; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_47; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_48; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_49; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_50; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_51; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_52; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_53; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_54; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_55; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_56; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_57; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_58; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_59; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_60; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_61; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_62; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_63; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_64; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_65; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_66; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_67; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_68; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_69; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_70; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_71; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_72; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_73; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_74; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_75; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_76; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_77; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_78; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_79; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_80; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_81; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_82; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_83; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_84; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_85; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_86; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_87; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_88; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_89; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_90; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_91; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_92; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_93; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_94; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_95; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_96; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_97; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_98; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_99; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_100; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_101; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_102; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_103; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_104; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_105; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_106; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_107; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_108; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_109; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_110; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_111; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_112; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_113; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_114; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_115; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_116; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_117; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_118; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_119; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_120; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_121; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_122; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_123; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_124; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_125; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_126; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_127; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_128; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_129; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_130; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_131; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_132; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_133; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_134; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_135; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_136; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_137; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_138; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_139; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_140; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_141; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_142; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_143; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_144; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_145; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_146; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_147; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_148; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_149; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_150; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_151; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_152; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_153; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_154; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_155; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_156; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_157; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_158; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_159; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_160; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_161; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_162; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_163; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_164; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_165; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_166; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_167; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_168; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_169; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_170; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_171; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_172; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_173; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_174; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_175; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_176; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_177; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_178; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_179; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_180; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_181; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_182; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_183; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_184; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_185; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_186; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_187; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_188; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_189; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_190; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_191; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_192; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_193; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_194; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_195; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_196; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_197; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_198; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_199; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_200; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_201; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_202; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_203; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_204; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_205; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_206; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_207; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_208; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_209; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_210; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_211; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_212; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_213; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_214; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_215; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_216; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_217; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_218; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_219; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_220; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_221; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_222; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_223; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_224; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_225; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_226; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_227; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_228; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_229; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_230; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_231; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_232; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_233; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_234; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_235; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_236; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_237; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_238; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_239; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_240; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_241; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_242; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_243; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_244; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_245; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_246; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_247; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_248; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_249; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_250; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_251; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_252; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_253; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_254; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_255; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_256; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_257; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_258; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_259; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_260; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_261; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_262; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_263; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_264; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_265; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_266; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_267; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_268; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_269; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_270; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_271; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_272; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_273; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_274; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_275; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_276; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_277; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_278; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_279; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_280; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_281; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_282; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_283; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_284; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_285; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_286; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_287; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_288; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_289; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_290; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_291; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_292; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_293; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_294; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_295; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_296; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_297; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_298; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_299; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_300; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_301; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_302; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_303; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_304; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_305; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_306; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_307; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_308; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_309; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_310; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_311; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_312; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_313; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_314; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_315; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_316; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_317; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_318; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_319; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_320; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_321; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_322; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_323; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_324; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_325; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_326; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_327; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_328; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_329; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_330; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_331; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_332; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_333; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_334; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_335; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_336; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_337; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_338; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_339; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_340; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_341; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_342; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_343; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_344; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_345; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_346; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_347; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_348; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_349; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_350; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_351; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_352; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_353; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_354; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_355; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_356; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_357; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_358; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_359; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_360; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_361; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_362; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_363; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_364; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_365; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_366; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_367; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_368; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_369; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_370; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_371; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_372; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_373; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_374; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_375; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_376; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_377; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_378; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_379; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_380; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_381; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_382; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_383; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_384; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_385; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_386; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_387; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_388; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_389; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_390; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_391; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_392; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_393; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_394; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_395; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_396; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_397; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_398; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_399; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_400; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_401; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_402; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_403; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_404; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_405; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_406; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_407; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_408; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_409; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_410; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_411; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_412; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_413; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_414; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_415; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_416; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_417; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_418; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_419; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_420; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_421; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_422; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_423; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_424; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_425; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_426; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_427; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_428; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_429; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_430; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_431; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_432; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_433; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_434; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_435; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_436; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_437; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_438; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_439; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_440; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_441; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_442; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_443; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_444; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_445; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_446; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_447; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_448; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_449; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_450; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_451; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_452; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_453; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_454; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_455; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_456; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_457; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_458; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_459; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_460; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_461; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_462; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_463; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_464; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_465; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_466; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_467; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_468; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_469; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_470; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_471; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_472; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_473; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_474; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_475; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_476; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_477; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_478; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_479; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_480; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_481; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_482; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_483; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_484; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_485; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_486; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_487; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_488; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_489; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_490; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_491; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_492; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_493; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_494; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_495; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_496; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_497; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_498; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_499; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_500; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_501; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_502; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_503; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_504; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_505; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_506; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_507; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_508; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_509; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_510; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_511; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_512; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_513; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_514; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_515; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_516; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_517; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_518; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_519; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_520; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_521; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_522; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_523; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_524; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_525; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_526; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_527; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_528; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_529; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_530; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_531; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_532; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_533; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_534; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_535; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_536; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_537; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_538; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_539; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_540; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_541; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_542; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_543; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_544; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_545; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_546; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_547; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_548; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_549; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_550; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_551; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_552; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_553; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_554; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_555; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_556; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_557; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_558; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_559; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_560; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_561; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_562; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_563; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_564; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_565; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_566; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_567; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_568; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_569; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_570; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_571; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_572; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_573; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_574; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_575; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_576; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_577; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_578; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_579; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_580; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_581; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_582; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_583; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_584; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_585; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_586; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_587; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_588; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_589; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_590; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_591; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_592; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_593; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_594; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_595; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_596; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_597; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_598; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_599; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_600; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_601; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_602; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_603; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_604; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_605; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_606; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_607; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_608; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_609; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_610; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_611; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_612; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_613; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_614; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_615; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_616; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_617; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_618; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_619; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_620; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_621; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_622; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_623; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_624; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_625; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_626; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_627; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_628; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_629; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_630; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_631; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_632; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_633; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_634; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_635; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_636; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_637; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_638; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_639; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_640; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_641; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_642; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_643; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_644; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_645; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_646; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_647; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_648; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_649; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_650; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_651; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_652; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_653; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_654; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_655; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_656; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_657; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_658; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_659; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_660; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_661; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_662; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_663; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_664; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_665; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_666; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_667; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_668; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_669; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_670; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_671; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_672; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_673; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_674; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_675; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_676; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_677; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_678; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_679; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_680; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_681; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_682; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_683; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_684; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_685; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_686; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_687; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_688; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_689; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_690; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_691; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_692; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_693; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_694; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_695; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_696; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_697; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_698; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_699; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_700; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_701; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_702; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_703; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_704; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_705; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_706; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_707; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_708; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_709; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_710; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_711; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_712; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_713; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_714; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_715; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_716; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_717; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_718; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_719; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_720; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_721; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_722; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_723; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_724; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_725; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_726; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_727; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_728; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_729; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_730; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_731; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_732; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_733; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_734; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_735; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_736; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_737; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_738; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_739; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_740; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_741; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_742; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_743; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_744; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_745; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_746; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_747; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_748; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_749; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_750; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_751; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_752; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_753; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_754; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_755; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_756; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_757; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_758; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_759; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_760; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_761; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_762; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_763; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_764; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_765; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_766; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_767; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_768; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_769; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_770; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_771; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_772; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_773; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_774; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_775; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_776; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_777; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_778; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_779; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_780; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_781; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_782; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_783; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_784; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_785; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_786; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_787; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_788; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_789; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_790; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_791; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_792; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_793; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_794; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_795; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_796; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_797; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_798; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_799; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_800; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_801; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_802; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_803; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_804; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_805; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_806; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_807; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_808; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_809; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_810; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_811; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_812; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_813; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_814; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_815; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_816; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_817; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_818; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_819; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_820; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_821; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_822; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_823; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_824; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_825; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_826; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_827; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_828; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_829; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_830; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_831; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_832; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_833; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_834; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_835; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_836; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_837; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_838; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_839; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_840; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_841; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_842; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_843; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_844; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_845; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_846; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_847; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_848; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_849; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_850; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_851; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_852; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_853; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_854; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_855; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_856; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_857; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_858; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_859; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_860; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_861; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_862; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_863; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_864; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_865; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_866; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_867; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_868; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_869; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_870; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_871; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_872; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_873; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_874; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_875; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_876; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_877; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_878; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_879; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_880; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_881; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_882; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_883; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_884; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_885; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_886; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_887; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_888; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_889; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_890; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_891; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_892; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_893; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_894; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_895; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_896; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_897; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_898; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_899; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_900; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_901; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_902; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_903; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_904; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_905; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_906; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_907; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_908; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_909; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_910; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_911; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_912; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_913; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_914; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_915; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_916; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_917; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_918; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_919; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_920; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_921; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_922; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_923; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_924; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_925; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_926; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_927; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_928; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_929; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_930; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_931; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_932; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_933; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_934; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_935; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_936; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_937; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_938; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_939; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_940; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_941; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_942; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_943; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_944; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_945; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_946; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_947; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_948; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_949; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_950; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_951; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_952; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_953; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_954; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_955; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_956; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_957; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_958; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_959; // @[RAM_ST.scala 31:71]
  wire [10:0] _T; // @[RAM_ST.scala 31:71]
  wire [9:0] _GEN_966; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_967; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_968; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_969; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_970; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_971; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_972; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_973; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_974; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_975; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_976; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_977; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_978; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_979; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_980; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_981; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_982; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_983; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_984; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_985; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_986; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_987; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_988; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_989; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_990; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_991; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_992; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_993; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_994; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_995; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_996; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_997; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_998; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_999; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1000; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1001; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1002; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1003; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1004; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1005; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1006; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1007; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1008; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1009; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1010; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1011; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1012; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1013; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1014; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1015; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1016; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1017; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1018; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1019; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1020; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1021; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1022; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1023; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1024; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1025; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1026; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1027; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1028; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1029; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1030; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1031; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1032; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1033; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1034; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1035; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1036; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1037; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1038; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1039; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1040; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1041; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1042; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1043; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1044; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1045; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1046; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1047; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1048; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1049; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1050; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1051; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1052; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1053; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1054; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1055; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1056; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1057; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1058; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1059; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1060; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1061; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1062; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1063; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1064; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1065; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1066; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1067; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1068; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1069; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1070; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1071; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1072; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1073; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1074; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1075; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1076; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1077; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1078; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1079; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1080; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1081; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1082; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1083; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1084; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1085; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1086; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1087; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1088; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1089; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1090; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1091; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1092; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1093; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1094; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1095; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1096; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1097; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1098; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1099; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1100; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1101; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1102; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1103; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1104; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1105; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1106; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1107; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1108; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1109; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1110; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1111; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1112; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1113; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1114; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1115; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1116; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1117; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1118; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1119; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1120; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1121; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1122; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1123; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1124; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1125; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1126; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1127; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1128; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1129; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1130; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1131; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1132; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1133; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1134; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1135; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1136; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1137; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1138; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1139; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1140; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1141; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1142; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1143; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1144; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1145; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1146; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1147; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1148; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1149; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1150; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1151; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1152; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1153; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1154; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1155; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1156; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1157; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1158; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1159; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1160; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1161; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1162; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1163; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1164; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1165; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1166; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1167; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1168; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1169; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1170; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1171; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1172; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1173; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1174; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1175; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1176; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1177; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1178; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1179; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1180; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1181; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1182; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1183; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1184; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1185; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1186; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1187; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1188; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1189; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1190; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1191; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1192; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1193; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1194; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1195; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1196; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1197; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1198; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1199; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1200; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1201; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1202; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1203; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1204; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1205; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1206; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1207; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1208; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1209; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1210; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1211; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1212; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1213; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1214; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1215; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1216; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1217; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1218; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1219; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1220; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1221; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1222; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1223; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1224; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1225; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1226; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1227; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1228; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1229; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1230; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1231; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1232; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1233; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1234; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1235; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1236; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1237; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1238; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1239; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1240; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1241; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1242; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1243; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1244; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1245; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1246; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1247; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1248; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1249; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1250; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1251; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1252; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1253; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1254; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1255; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1256; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1257; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1258; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1259; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1260; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1261; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1262; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1263; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1264; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1265; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1266; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1267; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1268; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1269; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1270; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1271; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1272; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1273; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1274; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1275; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1276; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1277; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1278; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1279; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1280; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1281; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1282; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1283; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1284; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1285; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1286; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1287; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1288; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1289; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1290; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1291; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1292; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1293; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1294; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1295; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1296; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1297; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1298; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1299; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1300; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1301; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1302; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1303; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1304; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1305; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1306; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1307; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1308; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1309; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1310; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1311; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1312; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1313; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1314; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1315; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1316; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1317; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1318; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1319; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1320; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1321; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1322; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1323; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1324; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1325; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1326; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1327; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1328; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1329; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1330; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1331; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1332; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1333; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1334; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1335; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1336; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1337; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1338; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1339; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1340; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1341; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1342; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1343; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1344; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1345; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1346; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1347; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1348; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1349; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1350; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1351; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1352; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1353; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1354; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1355; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1356; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1357; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1358; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1359; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1360; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1361; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1362; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1363; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1364; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1365; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1366; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1367; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1368; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1369; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1370; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1371; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1372; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1373; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1374; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1375; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1376; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1377; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1378; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1379; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1380; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1381; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1382; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1383; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1384; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1385; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1386; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1387; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1388; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1389; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1390; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1391; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1392; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1393; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1394; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1395; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1396; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1397; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1398; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1399; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1400; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1401; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1402; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1403; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1404; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1405; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1406; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1407; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1408; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1409; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1410; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1411; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1412; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1413; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1414; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1415; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1416; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1417; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1418; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1419; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1420; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1421; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1422; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1423; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1424; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1425; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1426; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1427; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1428; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1429; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1430; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1431; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1432; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1433; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1434; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1435; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1436; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1437; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1438; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1439; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1440; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1441; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1442; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1443; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1444; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1445; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1446; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1447; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1448; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1449; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1450; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1451; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1452; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1453; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1454; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1455; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1456; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1457; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1458; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1459; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1460; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1461; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1462; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1463; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1464; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1465; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1466; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1467; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1468; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1469; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1470; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1471; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1472; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1473; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1474; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1475; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1476; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1477; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1478; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1479; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1480; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1481; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1482; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1483; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1484; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1485; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1486; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1487; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1488; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1489; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1490; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1491; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1492; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1493; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1494; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1495; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1496; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1497; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1498; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1499; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1500; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1501; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1502; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1503; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1504; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1505; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1506; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1507; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1508; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1509; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1510; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1511; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1512; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1513; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1514; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1515; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1516; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1517; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1518; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1519; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1520; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1521; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1522; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1523; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1524; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1525; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1526; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1527; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1528; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1529; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1530; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1531; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1532; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1533; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1534; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1535; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1536; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1537; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1538; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1539; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1540; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1541; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1542; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1543; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1544; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1545; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1546; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1547; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1548; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1549; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1550; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1551; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1552; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1553; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1554; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1555; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1556; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1557; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1558; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1559; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1560; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1561; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1562; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1563; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1564; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1565; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1566; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1567; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1568; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1569; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1570; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1571; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1572; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1573; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1574; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1575; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1576; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1577; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1578; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1579; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1580; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1581; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1582; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1583; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1584; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1585; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1586; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1587; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1588; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1589; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1590; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1591; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1592; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1593; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1594; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1595; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1596; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1597; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1598; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1599; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1600; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1601; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1602; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1603; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1604; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1605; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1606; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1607; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1608; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1609; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1610; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1611; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1612; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1613; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1614; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1615; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1616; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1617; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1618; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1619; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1620; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1621; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1622; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1623; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1624; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1625; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1626; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1627; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1628; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1629; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1630; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1631; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1632; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1633; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1634; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1635; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1636; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1637; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1638; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1639; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1640; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1641; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1642; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1643; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1644; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1645; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1646; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1647; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1648; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1649; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1650; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1651; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1652; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1653; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1654; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1655; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1656; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1657; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1658; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1659; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1660; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1661; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1662; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1663; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1664; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1665; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1666; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1667; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1668; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1669; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1670; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1671; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1672; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1673; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1674; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1675; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1676; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1677; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1678; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1679; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1680; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1681; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1682; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1683; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1684; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1685; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1686; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1687; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1688; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1689; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1690; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1691; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1692; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1693; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1694; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1695; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1696; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1697; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1698; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1699; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1700; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1701; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1702; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1703; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1704; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1705; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1706; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1707; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1708; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1709; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1710; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1711; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1712; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1713; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1714; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1715; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1716; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1717; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1718; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1719; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1720; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1721; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1722; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1723; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1724; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1725; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1726; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1727; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1728; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1729; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1730; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1731; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1732; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1733; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1734; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1735; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1736; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1737; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1738; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1739; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1740; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1741; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1742; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1743; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1744; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1745; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1746; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1747; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1748; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1749; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1750; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1751; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1752; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1753; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1754; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1755; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1756; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1757; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1758; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1759; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1760; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1761; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1762; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1763; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1764; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1765; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1766; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1767; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1768; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1769; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1770; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1771; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1772; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1773; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1774; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1775; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1776; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1777; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1778; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1779; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1780; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1781; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1782; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1783; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1784; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1785; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1786; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1787; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1788; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1789; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1790; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1791; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1792; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1793; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1794; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1795; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1796; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1797; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1798; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1799; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1800; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1801; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1802; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1803; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1804; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1805; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1806; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1807; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1808; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1809; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1810; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1811; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1812; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1813; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1814; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1815; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1816; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1817; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1818; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1819; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1820; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1821; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1822; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1823; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1824; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1825; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1826; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1827; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1828; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1829; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1830; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1831; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1832; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1833; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1834; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1835; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1836; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1837; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1838; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1839; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1840; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1841; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1842; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1843; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1844; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1845; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1846; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1847; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1848; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1849; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1850; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1851; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1852; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1853; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1854; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1855; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1856; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1857; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1858; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1859; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1860; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1861; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1862; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1863; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1864; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1865; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1866; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1867; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1868; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1869; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1870; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1871; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1872; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1873; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1874; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1875; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1876; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1877; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1878; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1879; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1880; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1881; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1882; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1883; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1884; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1885; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1886; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1887; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1888; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1889; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1890; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1891; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1892; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1893; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1894; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1895; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1896; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1897; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1898; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1899; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1900; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1901; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1902; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1903; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1904; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1905; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1906; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1907; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1908; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1909; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1910; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1911; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1912; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1913; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1914; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1915; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1916; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1917; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1918; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1919; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1920; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1921; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1922; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1923; // @[RAM_ST.scala 32:46]
  wire [9:0] _GEN_1924; // @[RAM_ST.scala 32:46]
  wire [10:0] _T_4; // @[RAM_ST.scala 32:46]
  wire [15:0] _T_11;
  NestedCountersWithNumValid write_elem_counter ( // @[RAM_ST.scala 20:34]
    .CE(write_elem_counter_CE),
    .valid(write_elem_counter_valid)
  );
  NestedCountersWithNumValid read_elem_counter ( // @[RAM_ST.scala 21:33]
    .CE(read_elem_counter_CE),
    .valid(read_elem_counter_valid)
  );
  assign ram__T_9_addr = ram__T_9_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram__T_9_data = ram[ram__T_9_addr]; // @[RAM_ST.scala 29:24]
  `else
  assign ram__T_9_data = ram__T_9_addr >= 10'h3c0 ? _RAND_1[15:0] : ram[ram__T_9_addr]; // @[RAM_ST.scala 29:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram__T_3_data = {WDATA_1,WDATA_0};
  assign ram__T_3_addr = _T[9:0];
  assign ram__T_3_mask = 1'h1;
  assign ram__T_3_en = write_elem_counter_valid;
  assign _GEN_1 = 10'h1 == WADDR ? 10'h1 : 10'h0; // @[RAM_ST.scala 31:71]
  assign _GEN_2 = 10'h2 == WADDR ? 10'h2 : _GEN_1; // @[RAM_ST.scala 31:71]
  assign _GEN_3 = 10'h3 == WADDR ? 10'h3 : _GEN_2; // @[RAM_ST.scala 31:71]
  assign _GEN_4 = 10'h4 == WADDR ? 10'h4 : _GEN_3; // @[RAM_ST.scala 31:71]
  assign _GEN_5 = 10'h5 == WADDR ? 10'h5 : _GEN_4; // @[RAM_ST.scala 31:71]
  assign _GEN_6 = 10'h6 == WADDR ? 10'h6 : _GEN_5; // @[RAM_ST.scala 31:71]
  assign _GEN_7 = 10'h7 == WADDR ? 10'h7 : _GEN_6; // @[RAM_ST.scala 31:71]
  assign _GEN_8 = 10'h8 == WADDR ? 10'h8 : _GEN_7; // @[RAM_ST.scala 31:71]
  assign _GEN_9 = 10'h9 == WADDR ? 10'h9 : _GEN_8; // @[RAM_ST.scala 31:71]
  assign _GEN_10 = 10'ha == WADDR ? 10'ha : _GEN_9; // @[RAM_ST.scala 31:71]
  assign _GEN_11 = 10'hb == WADDR ? 10'hb : _GEN_10; // @[RAM_ST.scala 31:71]
  assign _GEN_12 = 10'hc == WADDR ? 10'hc : _GEN_11; // @[RAM_ST.scala 31:71]
  assign _GEN_13 = 10'hd == WADDR ? 10'hd : _GEN_12; // @[RAM_ST.scala 31:71]
  assign _GEN_14 = 10'he == WADDR ? 10'he : _GEN_13; // @[RAM_ST.scala 31:71]
  assign _GEN_15 = 10'hf == WADDR ? 10'hf : _GEN_14; // @[RAM_ST.scala 31:71]
  assign _GEN_16 = 10'h10 == WADDR ? 10'h10 : _GEN_15; // @[RAM_ST.scala 31:71]
  assign _GEN_17 = 10'h11 == WADDR ? 10'h11 : _GEN_16; // @[RAM_ST.scala 31:71]
  assign _GEN_18 = 10'h12 == WADDR ? 10'h12 : _GEN_17; // @[RAM_ST.scala 31:71]
  assign _GEN_19 = 10'h13 == WADDR ? 10'h13 : _GEN_18; // @[RAM_ST.scala 31:71]
  assign _GEN_20 = 10'h14 == WADDR ? 10'h14 : _GEN_19; // @[RAM_ST.scala 31:71]
  assign _GEN_21 = 10'h15 == WADDR ? 10'h15 : _GEN_20; // @[RAM_ST.scala 31:71]
  assign _GEN_22 = 10'h16 == WADDR ? 10'h16 : _GEN_21; // @[RAM_ST.scala 31:71]
  assign _GEN_23 = 10'h17 == WADDR ? 10'h17 : _GEN_22; // @[RAM_ST.scala 31:71]
  assign _GEN_24 = 10'h18 == WADDR ? 10'h18 : _GEN_23; // @[RAM_ST.scala 31:71]
  assign _GEN_25 = 10'h19 == WADDR ? 10'h19 : _GEN_24; // @[RAM_ST.scala 31:71]
  assign _GEN_26 = 10'h1a == WADDR ? 10'h1a : _GEN_25; // @[RAM_ST.scala 31:71]
  assign _GEN_27 = 10'h1b == WADDR ? 10'h1b : _GEN_26; // @[RAM_ST.scala 31:71]
  assign _GEN_28 = 10'h1c == WADDR ? 10'h1c : _GEN_27; // @[RAM_ST.scala 31:71]
  assign _GEN_29 = 10'h1d == WADDR ? 10'h1d : _GEN_28; // @[RAM_ST.scala 31:71]
  assign _GEN_30 = 10'h1e == WADDR ? 10'h1e : _GEN_29; // @[RAM_ST.scala 31:71]
  assign _GEN_31 = 10'h1f == WADDR ? 10'h1f : _GEN_30; // @[RAM_ST.scala 31:71]
  assign _GEN_32 = 10'h20 == WADDR ? 10'h20 : _GEN_31; // @[RAM_ST.scala 31:71]
  assign _GEN_33 = 10'h21 == WADDR ? 10'h21 : _GEN_32; // @[RAM_ST.scala 31:71]
  assign _GEN_34 = 10'h22 == WADDR ? 10'h22 : _GEN_33; // @[RAM_ST.scala 31:71]
  assign _GEN_35 = 10'h23 == WADDR ? 10'h23 : _GEN_34; // @[RAM_ST.scala 31:71]
  assign _GEN_36 = 10'h24 == WADDR ? 10'h24 : _GEN_35; // @[RAM_ST.scala 31:71]
  assign _GEN_37 = 10'h25 == WADDR ? 10'h25 : _GEN_36; // @[RAM_ST.scala 31:71]
  assign _GEN_38 = 10'h26 == WADDR ? 10'h26 : _GEN_37; // @[RAM_ST.scala 31:71]
  assign _GEN_39 = 10'h27 == WADDR ? 10'h27 : _GEN_38; // @[RAM_ST.scala 31:71]
  assign _GEN_40 = 10'h28 == WADDR ? 10'h28 : _GEN_39; // @[RAM_ST.scala 31:71]
  assign _GEN_41 = 10'h29 == WADDR ? 10'h29 : _GEN_40; // @[RAM_ST.scala 31:71]
  assign _GEN_42 = 10'h2a == WADDR ? 10'h2a : _GEN_41; // @[RAM_ST.scala 31:71]
  assign _GEN_43 = 10'h2b == WADDR ? 10'h2b : _GEN_42; // @[RAM_ST.scala 31:71]
  assign _GEN_44 = 10'h2c == WADDR ? 10'h2c : _GEN_43; // @[RAM_ST.scala 31:71]
  assign _GEN_45 = 10'h2d == WADDR ? 10'h2d : _GEN_44; // @[RAM_ST.scala 31:71]
  assign _GEN_46 = 10'h2e == WADDR ? 10'h2e : _GEN_45; // @[RAM_ST.scala 31:71]
  assign _GEN_47 = 10'h2f == WADDR ? 10'h2f : _GEN_46; // @[RAM_ST.scala 31:71]
  assign _GEN_48 = 10'h30 == WADDR ? 10'h30 : _GEN_47; // @[RAM_ST.scala 31:71]
  assign _GEN_49 = 10'h31 == WADDR ? 10'h31 : _GEN_48; // @[RAM_ST.scala 31:71]
  assign _GEN_50 = 10'h32 == WADDR ? 10'h32 : _GEN_49; // @[RAM_ST.scala 31:71]
  assign _GEN_51 = 10'h33 == WADDR ? 10'h33 : _GEN_50; // @[RAM_ST.scala 31:71]
  assign _GEN_52 = 10'h34 == WADDR ? 10'h34 : _GEN_51; // @[RAM_ST.scala 31:71]
  assign _GEN_53 = 10'h35 == WADDR ? 10'h35 : _GEN_52; // @[RAM_ST.scala 31:71]
  assign _GEN_54 = 10'h36 == WADDR ? 10'h36 : _GEN_53; // @[RAM_ST.scala 31:71]
  assign _GEN_55 = 10'h37 == WADDR ? 10'h37 : _GEN_54; // @[RAM_ST.scala 31:71]
  assign _GEN_56 = 10'h38 == WADDR ? 10'h38 : _GEN_55; // @[RAM_ST.scala 31:71]
  assign _GEN_57 = 10'h39 == WADDR ? 10'h39 : _GEN_56; // @[RAM_ST.scala 31:71]
  assign _GEN_58 = 10'h3a == WADDR ? 10'h3a : _GEN_57; // @[RAM_ST.scala 31:71]
  assign _GEN_59 = 10'h3b == WADDR ? 10'h3b : _GEN_58; // @[RAM_ST.scala 31:71]
  assign _GEN_60 = 10'h3c == WADDR ? 10'h3c : _GEN_59; // @[RAM_ST.scala 31:71]
  assign _GEN_61 = 10'h3d == WADDR ? 10'h3d : _GEN_60; // @[RAM_ST.scala 31:71]
  assign _GEN_62 = 10'h3e == WADDR ? 10'h3e : _GEN_61; // @[RAM_ST.scala 31:71]
  assign _GEN_63 = 10'h3f == WADDR ? 10'h3f : _GEN_62; // @[RAM_ST.scala 31:71]
  assign _GEN_64 = 10'h40 == WADDR ? 10'h40 : _GEN_63; // @[RAM_ST.scala 31:71]
  assign _GEN_65 = 10'h41 == WADDR ? 10'h41 : _GEN_64; // @[RAM_ST.scala 31:71]
  assign _GEN_66 = 10'h42 == WADDR ? 10'h42 : _GEN_65; // @[RAM_ST.scala 31:71]
  assign _GEN_67 = 10'h43 == WADDR ? 10'h43 : _GEN_66; // @[RAM_ST.scala 31:71]
  assign _GEN_68 = 10'h44 == WADDR ? 10'h44 : _GEN_67; // @[RAM_ST.scala 31:71]
  assign _GEN_69 = 10'h45 == WADDR ? 10'h45 : _GEN_68; // @[RAM_ST.scala 31:71]
  assign _GEN_70 = 10'h46 == WADDR ? 10'h46 : _GEN_69; // @[RAM_ST.scala 31:71]
  assign _GEN_71 = 10'h47 == WADDR ? 10'h47 : _GEN_70; // @[RAM_ST.scala 31:71]
  assign _GEN_72 = 10'h48 == WADDR ? 10'h48 : _GEN_71; // @[RAM_ST.scala 31:71]
  assign _GEN_73 = 10'h49 == WADDR ? 10'h49 : _GEN_72; // @[RAM_ST.scala 31:71]
  assign _GEN_74 = 10'h4a == WADDR ? 10'h4a : _GEN_73; // @[RAM_ST.scala 31:71]
  assign _GEN_75 = 10'h4b == WADDR ? 10'h4b : _GEN_74; // @[RAM_ST.scala 31:71]
  assign _GEN_76 = 10'h4c == WADDR ? 10'h4c : _GEN_75; // @[RAM_ST.scala 31:71]
  assign _GEN_77 = 10'h4d == WADDR ? 10'h4d : _GEN_76; // @[RAM_ST.scala 31:71]
  assign _GEN_78 = 10'h4e == WADDR ? 10'h4e : _GEN_77; // @[RAM_ST.scala 31:71]
  assign _GEN_79 = 10'h4f == WADDR ? 10'h4f : _GEN_78; // @[RAM_ST.scala 31:71]
  assign _GEN_80 = 10'h50 == WADDR ? 10'h50 : _GEN_79; // @[RAM_ST.scala 31:71]
  assign _GEN_81 = 10'h51 == WADDR ? 10'h51 : _GEN_80; // @[RAM_ST.scala 31:71]
  assign _GEN_82 = 10'h52 == WADDR ? 10'h52 : _GEN_81; // @[RAM_ST.scala 31:71]
  assign _GEN_83 = 10'h53 == WADDR ? 10'h53 : _GEN_82; // @[RAM_ST.scala 31:71]
  assign _GEN_84 = 10'h54 == WADDR ? 10'h54 : _GEN_83; // @[RAM_ST.scala 31:71]
  assign _GEN_85 = 10'h55 == WADDR ? 10'h55 : _GEN_84; // @[RAM_ST.scala 31:71]
  assign _GEN_86 = 10'h56 == WADDR ? 10'h56 : _GEN_85; // @[RAM_ST.scala 31:71]
  assign _GEN_87 = 10'h57 == WADDR ? 10'h57 : _GEN_86; // @[RAM_ST.scala 31:71]
  assign _GEN_88 = 10'h58 == WADDR ? 10'h58 : _GEN_87; // @[RAM_ST.scala 31:71]
  assign _GEN_89 = 10'h59 == WADDR ? 10'h59 : _GEN_88; // @[RAM_ST.scala 31:71]
  assign _GEN_90 = 10'h5a == WADDR ? 10'h5a : _GEN_89; // @[RAM_ST.scala 31:71]
  assign _GEN_91 = 10'h5b == WADDR ? 10'h5b : _GEN_90; // @[RAM_ST.scala 31:71]
  assign _GEN_92 = 10'h5c == WADDR ? 10'h5c : _GEN_91; // @[RAM_ST.scala 31:71]
  assign _GEN_93 = 10'h5d == WADDR ? 10'h5d : _GEN_92; // @[RAM_ST.scala 31:71]
  assign _GEN_94 = 10'h5e == WADDR ? 10'h5e : _GEN_93; // @[RAM_ST.scala 31:71]
  assign _GEN_95 = 10'h5f == WADDR ? 10'h5f : _GEN_94; // @[RAM_ST.scala 31:71]
  assign _GEN_96 = 10'h60 == WADDR ? 10'h60 : _GEN_95; // @[RAM_ST.scala 31:71]
  assign _GEN_97 = 10'h61 == WADDR ? 10'h61 : _GEN_96; // @[RAM_ST.scala 31:71]
  assign _GEN_98 = 10'h62 == WADDR ? 10'h62 : _GEN_97; // @[RAM_ST.scala 31:71]
  assign _GEN_99 = 10'h63 == WADDR ? 10'h63 : _GEN_98; // @[RAM_ST.scala 31:71]
  assign _GEN_100 = 10'h64 == WADDR ? 10'h64 : _GEN_99; // @[RAM_ST.scala 31:71]
  assign _GEN_101 = 10'h65 == WADDR ? 10'h65 : _GEN_100; // @[RAM_ST.scala 31:71]
  assign _GEN_102 = 10'h66 == WADDR ? 10'h66 : _GEN_101; // @[RAM_ST.scala 31:71]
  assign _GEN_103 = 10'h67 == WADDR ? 10'h67 : _GEN_102; // @[RAM_ST.scala 31:71]
  assign _GEN_104 = 10'h68 == WADDR ? 10'h68 : _GEN_103; // @[RAM_ST.scala 31:71]
  assign _GEN_105 = 10'h69 == WADDR ? 10'h69 : _GEN_104; // @[RAM_ST.scala 31:71]
  assign _GEN_106 = 10'h6a == WADDR ? 10'h6a : _GEN_105; // @[RAM_ST.scala 31:71]
  assign _GEN_107 = 10'h6b == WADDR ? 10'h6b : _GEN_106; // @[RAM_ST.scala 31:71]
  assign _GEN_108 = 10'h6c == WADDR ? 10'h6c : _GEN_107; // @[RAM_ST.scala 31:71]
  assign _GEN_109 = 10'h6d == WADDR ? 10'h6d : _GEN_108; // @[RAM_ST.scala 31:71]
  assign _GEN_110 = 10'h6e == WADDR ? 10'h6e : _GEN_109; // @[RAM_ST.scala 31:71]
  assign _GEN_111 = 10'h6f == WADDR ? 10'h6f : _GEN_110; // @[RAM_ST.scala 31:71]
  assign _GEN_112 = 10'h70 == WADDR ? 10'h70 : _GEN_111; // @[RAM_ST.scala 31:71]
  assign _GEN_113 = 10'h71 == WADDR ? 10'h71 : _GEN_112; // @[RAM_ST.scala 31:71]
  assign _GEN_114 = 10'h72 == WADDR ? 10'h72 : _GEN_113; // @[RAM_ST.scala 31:71]
  assign _GEN_115 = 10'h73 == WADDR ? 10'h73 : _GEN_114; // @[RAM_ST.scala 31:71]
  assign _GEN_116 = 10'h74 == WADDR ? 10'h74 : _GEN_115; // @[RAM_ST.scala 31:71]
  assign _GEN_117 = 10'h75 == WADDR ? 10'h75 : _GEN_116; // @[RAM_ST.scala 31:71]
  assign _GEN_118 = 10'h76 == WADDR ? 10'h76 : _GEN_117; // @[RAM_ST.scala 31:71]
  assign _GEN_119 = 10'h77 == WADDR ? 10'h77 : _GEN_118; // @[RAM_ST.scala 31:71]
  assign _GEN_120 = 10'h78 == WADDR ? 10'h78 : _GEN_119; // @[RAM_ST.scala 31:71]
  assign _GEN_121 = 10'h79 == WADDR ? 10'h79 : _GEN_120; // @[RAM_ST.scala 31:71]
  assign _GEN_122 = 10'h7a == WADDR ? 10'h7a : _GEN_121; // @[RAM_ST.scala 31:71]
  assign _GEN_123 = 10'h7b == WADDR ? 10'h7b : _GEN_122; // @[RAM_ST.scala 31:71]
  assign _GEN_124 = 10'h7c == WADDR ? 10'h7c : _GEN_123; // @[RAM_ST.scala 31:71]
  assign _GEN_125 = 10'h7d == WADDR ? 10'h7d : _GEN_124; // @[RAM_ST.scala 31:71]
  assign _GEN_126 = 10'h7e == WADDR ? 10'h7e : _GEN_125; // @[RAM_ST.scala 31:71]
  assign _GEN_127 = 10'h7f == WADDR ? 10'h7f : _GEN_126; // @[RAM_ST.scala 31:71]
  assign _GEN_128 = 10'h80 == WADDR ? 10'h80 : _GEN_127; // @[RAM_ST.scala 31:71]
  assign _GEN_129 = 10'h81 == WADDR ? 10'h81 : _GEN_128; // @[RAM_ST.scala 31:71]
  assign _GEN_130 = 10'h82 == WADDR ? 10'h82 : _GEN_129; // @[RAM_ST.scala 31:71]
  assign _GEN_131 = 10'h83 == WADDR ? 10'h83 : _GEN_130; // @[RAM_ST.scala 31:71]
  assign _GEN_132 = 10'h84 == WADDR ? 10'h84 : _GEN_131; // @[RAM_ST.scala 31:71]
  assign _GEN_133 = 10'h85 == WADDR ? 10'h85 : _GEN_132; // @[RAM_ST.scala 31:71]
  assign _GEN_134 = 10'h86 == WADDR ? 10'h86 : _GEN_133; // @[RAM_ST.scala 31:71]
  assign _GEN_135 = 10'h87 == WADDR ? 10'h87 : _GEN_134; // @[RAM_ST.scala 31:71]
  assign _GEN_136 = 10'h88 == WADDR ? 10'h88 : _GEN_135; // @[RAM_ST.scala 31:71]
  assign _GEN_137 = 10'h89 == WADDR ? 10'h89 : _GEN_136; // @[RAM_ST.scala 31:71]
  assign _GEN_138 = 10'h8a == WADDR ? 10'h8a : _GEN_137; // @[RAM_ST.scala 31:71]
  assign _GEN_139 = 10'h8b == WADDR ? 10'h8b : _GEN_138; // @[RAM_ST.scala 31:71]
  assign _GEN_140 = 10'h8c == WADDR ? 10'h8c : _GEN_139; // @[RAM_ST.scala 31:71]
  assign _GEN_141 = 10'h8d == WADDR ? 10'h8d : _GEN_140; // @[RAM_ST.scala 31:71]
  assign _GEN_142 = 10'h8e == WADDR ? 10'h8e : _GEN_141; // @[RAM_ST.scala 31:71]
  assign _GEN_143 = 10'h8f == WADDR ? 10'h8f : _GEN_142; // @[RAM_ST.scala 31:71]
  assign _GEN_144 = 10'h90 == WADDR ? 10'h90 : _GEN_143; // @[RAM_ST.scala 31:71]
  assign _GEN_145 = 10'h91 == WADDR ? 10'h91 : _GEN_144; // @[RAM_ST.scala 31:71]
  assign _GEN_146 = 10'h92 == WADDR ? 10'h92 : _GEN_145; // @[RAM_ST.scala 31:71]
  assign _GEN_147 = 10'h93 == WADDR ? 10'h93 : _GEN_146; // @[RAM_ST.scala 31:71]
  assign _GEN_148 = 10'h94 == WADDR ? 10'h94 : _GEN_147; // @[RAM_ST.scala 31:71]
  assign _GEN_149 = 10'h95 == WADDR ? 10'h95 : _GEN_148; // @[RAM_ST.scala 31:71]
  assign _GEN_150 = 10'h96 == WADDR ? 10'h96 : _GEN_149; // @[RAM_ST.scala 31:71]
  assign _GEN_151 = 10'h97 == WADDR ? 10'h97 : _GEN_150; // @[RAM_ST.scala 31:71]
  assign _GEN_152 = 10'h98 == WADDR ? 10'h98 : _GEN_151; // @[RAM_ST.scala 31:71]
  assign _GEN_153 = 10'h99 == WADDR ? 10'h99 : _GEN_152; // @[RAM_ST.scala 31:71]
  assign _GEN_154 = 10'h9a == WADDR ? 10'h9a : _GEN_153; // @[RAM_ST.scala 31:71]
  assign _GEN_155 = 10'h9b == WADDR ? 10'h9b : _GEN_154; // @[RAM_ST.scala 31:71]
  assign _GEN_156 = 10'h9c == WADDR ? 10'h9c : _GEN_155; // @[RAM_ST.scala 31:71]
  assign _GEN_157 = 10'h9d == WADDR ? 10'h9d : _GEN_156; // @[RAM_ST.scala 31:71]
  assign _GEN_158 = 10'h9e == WADDR ? 10'h9e : _GEN_157; // @[RAM_ST.scala 31:71]
  assign _GEN_159 = 10'h9f == WADDR ? 10'h9f : _GEN_158; // @[RAM_ST.scala 31:71]
  assign _GEN_160 = 10'ha0 == WADDR ? 10'ha0 : _GEN_159; // @[RAM_ST.scala 31:71]
  assign _GEN_161 = 10'ha1 == WADDR ? 10'ha1 : _GEN_160; // @[RAM_ST.scala 31:71]
  assign _GEN_162 = 10'ha2 == WADDR ? 10'ha2 : _GEN_161; // @[RAM_ST.scala 31:71]
  assign _GEN_163 = 10'ha3 == WADDR ? 10'ha3 : _GEN_162; // @[RAM_ST.scala 31:71]
  assign _GEN_164 = 10'ha4 == WADDR ? 10'ha4 : _GEN_163; // @[RAM_ST.scala 31:71]
  assign _GEN_165 = 10'ha5 == WADDR ? 10'ha5 : _GEN_164; // @[RAM_ST.scala 31:71]
  assign _GEN_166 = 10'ha6 == WADDR ? 10'ha6 : _GEN_165; // @[RAM_ST.scala 31:71]
  assign _GEN_167 = 10'ha7 == WADDR ? 10'ha7 : _GEN_166; // @[RAM_ST.scala 31:71]
  assign _GEN_168 = 10'ha8 == WADDR ? 10'ha8 : _GEN_167; // @[RAM_ST.scala 31:71]
  assign _GEN_169 = 10'ha9 == WADDR ? 10'ha9 : _GEN_168; // @[RAM_ST.scala 31:71]
  assign _GEN_170 = 10'haa == WADDR ? 10'haa : _GEN_169; // @[RAM_ST.scala 31:71]
  assign _GEN_171 = 10'hab == WADDR ? 10'hab : _GEN_170; // @[RAM_ST.scala 31:71]
  assign _GEN_172 = 10'hac == WADDR ? 10'hac : _GEN_171; // @[RAM_ST.scala 31:71]
  assign _GEN_173 = 10'had == WADDR ? 10'had : _GEN_172; // @[RAM_ST.scala 31:71]
  assign _GEN_174 = 10'hae == WADDR ? 10'hae : _GEN_173; // @[RAM_ST.scala 31:71]
  assign _GEN_175 = 10'haf == WADDR ? 10'haf : _GEN_174; // @[RAM_ST.scala 31:71]
  assign _GEN_176 = 10'hb0 == WADDR ? 10'hb0 : _GEN_175; // @[RAM_ST.scala 31:71]
  assign _GEN_177 = 10'hb1 == WADDR ? 10'hb1 : _GEN_176; // @[RAM_ST.scala 31:71]
  assign _GEN_178 = 10'hb2 == WADDR ? 10'hb2 : _GEN_177; // @[RAM_ST.scala 31:71]
  assign _GEN_179 = 10'hb3 == WADDR ? 10'hb3 : _GEN_178; // @[RAM_ST.scala 31:71]
  assign _GEN_180 = 10'hb4 == WADDR ? 10'hb4 : _GEN_179; // @[RAM_ST.scala 31:71]
  assign _GEN_181 = 10'hb5 == WADDR ? 10'hb5 : _GEN_180; // @[RAM_ST.scala 31:71]
  assign _GEN_182 = 10'hb6 == WADDR ? 10'hb6 : _GEN_181; // @[RAM_ST.scala 31:71]
  assign _GEN_183 = 10'hb7 == WADDR ? 10'hb7 : _GEN_182; // @[RAM_ST.scala 31:71]
  assign _GEN_184 = 10'hb8 == WADDR ? 10'hb8 : _GEN_183; // @[RAM_ST.scala 31:71]
  assign _GEN_185 = 10'hb9 == WADDR ? 10'hb9 : _GEN_184; // @[RAM_ST.scala 31:71]
  assign _GEN_186 = 10'hba == WADDR ? 10'hba : _GEN_185; // @[RAM_ST.scala 31:71]
  assign _GEN_187 = 10'hbb == WADDR ? 10'hbb : _GEN_186; // @[RAM_ST.scala 31:71]
  assign _GEN_188 = 10'hbc == WADDR ? 10'hbc : _GEN_187; // @[RAM_ST.scala 31:71]
  assign _GEN_189 = 10'hbd == WADDR ? 10'hbd : _GEN_188; // @[RAM_ST.scala 31:71]
  assign _GEN_190 = 10'hbe == WADDR ? 10'hbe : _GEN_189; // @[RAM_ST.scala 31:71]
  assign _GEN_191 = 10'hbf == WADDR ? 10'hbf : _GEN_190; // @[RAM_ST.scala 31:71]
  assign _GEN_192 = 10'hc0 == WADDR ? 10'hc0 : _GEN_191; // @[RAM_ST.scala 31:71]
  assign _GEN_193 = 10'hc1 == WADDR ? 10'hc1 : _GEN_192; // @[RAM_ST.scala 31:71]
  assign _GEN_194 = 10'hc2 == WADDR ? 10'hc2 : _GEN_193; // @[RAM_ST.scala 31:71]
  assign _GEN_195 = 10'hc3 == WADDR ? 10'hc3 : _GEN_194; // @[RAM_ST.scala 31:71]
  assign _GEN_196 = 10'hc4 == WADDR ? 10'hc4 : _GEN_195; // @[RAM_ST.scala 31:71]
  assign _GEN_197 = 10'hc5 == WADDR ? 10'hc5 : _GEN_196; // @[RAM_ST.scala 31:71]
  assign _GEN_198 = 10'hc6 == WADDR ? 10'hc6 : _GEN_197; // @[RAM_ST.scala 31:71]
  assign _GEN_199 = 10'hc7 == WADDR ? 10'hc7 : _GEN_198; // @[RAM_ST.scala 31:71]
  assign _GEN_200 = 10'hc8 == WADDR ? 10'hc8 : _GEN_199; // @[RAM_ST.scala 31:71]
  assign _GEN_201 = 10'hc9 == WADDR ? 10'hc9 : _GEN_200; // @[RAM_ST.scala 31:71]
  assign _GEN_202 = 10'hca == WADDR ? 10'hca : _GEN_201; // @[RAM_ST.scala 31:71]
  assign _GEN_203 = 10'hcb == WADDR ? 10'hcb : _GEN_202; // @[RAM_ST.scala 31:71]
  assign _GEN_204 = 10'hcc == WADDR ? 10'hcc : _GEN_203; // @[RAM_ST.scala 31:71]
  assign _GEN_205 = 10'hcd == WADDR ? 10'hcd : _GEN_204; // @[RAM_ST.scala 31:71]
  assign _GEN_206 = 10'hce == WADDR ? 10'hce : _GEN_205; // @[RAM_ST.scala 31:71]
  assign _GEN_207 = 10'hcf == WADDR ? 10'hcf : _GEN_206; // @[RAM_ST.scala 31:71]
  assign _GEN_208 = 10'hd0 == WADDR ? 10'hd0 : _GEN_207; // @[RAM_ST.scala 31:71]
  assign _GEN_209 = 10'hd1 == WADDR ? 10'hd1 : _GEN_208; // @[RAM_ST.scala 31:71]
  assign _GEN_210 = 10'hd2 == WADDR ? 10'hd2 : _GEN_209; // @[RAM_ST.scala 31:71]
  assign _GEN_211 = 10'hd3 == WADDR ? 10'hd3 : _GEN_210; // @[RAM_ST.scala 31:71]
  assign _GEN_212 = 10'hd4 == WADDR ? 10'hd4 : _GEN_211; // @[RAM_ST.scala 31:71]
  assign _GEN_213 = 10'hd5 == WADDR ? 10'hd5 : _GEN_212; // @[RAM_ST.scala 31:71]
  assign _GEN_214 = 10'hd6 == WADDR ? 10'hd6 : _GEN_213; // @[RAM_ST.scala 31:71]
  assign _GEN_215 = 10'hd7 == WADDR ? 10'hd7 : _GEN_214; // @[RAM_ST.scala 31:71]
  assign _GEN_216 = 10'hd8 == WADDR ? 10'hd8 : _GEN_215; // @[RAM_ST.scala 31:71]
  assign _GEN_217 = 10'hd9 == WADDR ? 10'hd9 : _GEN_216; // @[RAM_ST.scala 31:71]
  assign _GEN_218 = 10'hda == WADDR ? 10'hda : _GEN_217; // @[RAM_ST.scala 31:71]
  assign _GEN_219 = 10'hdb == WADDR ? 10'hdb : _GEN_218; // @[RAM_ST.scala 31:71]
  assign _GEN_220 = 10'hdc == WADDR ? 10'hdc : _GEN_219; // @[RAM_ST.scala 31:71]
  assign _GEN_221 = 10'hdd == WADDR ? 10'hdd : _GEN_220; // @[RAM_ST.scala 31:71]
  assign _GEN_222 = 10'hde == WADDR ? 10'hde : _GEN_221; // @[RAM_ST.scala 31:71]
  assign _GEN_223 = 10'hdf == WADDR ? 10'hdf : _GEN_222; // @[RAM_ST.scala 31:71]
  assign _GEN_224 = 10'he0 == WADDR ? 10'he0 : _GEN_223; // @[RAM_ST.scala 31:71]
  assign _GEN_225 = 10'he1 == WADDR ? 10'he1 : _GEN_224; // @[RAM_ST.scala 31:71]
  assign _GEN_226 = 10'he2 == WADDR ? 10'he2 : _GEN_225; // @[RAM_ST.scala 31:71]
  assign _GEN_227 = 10'he3 == WADDR ? 10'he3 : _GEN_226; // @[RAM_ST.scala 31:71]
  assign _GEN_228 = 10'he4 == WADDR ? 10'he4 : _GEN_227; // @[RAM_ST.scala 31:71]
  assign _GEN_229 = 10'he5 == WADDR ? 10'he5 : _GEN_228; // @[RAM_ST.scala 31:71]
  assign _GEN_230 = 10'he6 == WADDR ? 10'he6 : _GEN_229; // @[RAM_ST.scala 31:71]
  assign _GEN_231 = 10'he7 == WADDR ? 10'he7 : _GEN_230; // @[RAM_ST.scala 31:71]
  assign _GEN_232 = 10'he8 == WADDR ? 10'he8 : _GEN_231; // @[RAM_ST.scala 31:71]
  assign _GEN_233 = 10'he9 == WADDR ? 10'he9 : _GEN_232; // @[RAM_ST.scala 31:71]
  assign _GEN_234 = 10'hea == WADDR ? 10'hea : _GEN_233; // @[RAM_ST.scala 31:71]
  assign _GEN_235 = 10'heb == WADDR ? 10'heb : _GEN_234; // @[RAM_ST.scala 31:71]
  assign _GEN_236 = 10'hec == WADDR ? 10'hec : _GEN_235; // @[RAM_ST.scala 31:71]
  assign _GEN_237 = 10'hed == WADDR ? 10'hed : _GEN_236; // @[RAM_ST.scala 31:71]
  assign _GEN_238 = 10'hee == WADDR ? 10'hee : _GEN_237; // @[RAM_ST.scala 31:71]
  assign _GEN_239 = 10'hef == WADDR ? 10'hef : _GEN_238; // @[RAM_ST.scala 31:71]
  assign _GEN_240 = 10'hf0 == WADDR ? 10'hf0 : _GEN_239; // @[RAM_ST.scala 31:71]
  assign _GEN_241 = 10'hf1 == WADDR ? 10'hf1 : _GEN_240; // @[RAM_ST.scala 31:71]
  assign _GEN_242 = 10'hf2 == WADDR ? 10'hf2 : _GEN_241; // @[RAM_ST.scala 31:71]
  assign _GEN_243 = 10'hf3 == WADDR ? 10'hf3 : _GEN_242; // @[RAM_ST.scala 31:71]
  assign _GEN_244 = 10'hf4 == WADDR ? 10'hf4 : _GEN_243; // @[RAM_ST.scala 31:71]
  assign _GEN_245 = 10'hf5 == WADDR ? 10'hf5 : _GEN_244; // @[RAM_ST.scala 31:71]
  assign _GEN_246 = 10'hf6 == WADDR ? 10'hf6 : _GEN_245; // @[RAM_ST.scala 31:71]
  assign _GEN_247 = 10'hf7 == WADDR ? 10'hf7 : _GEN_246; // @[RAM_ST.scala 31:71]
  assign _GEN_248 = 10'hf8 == WADDR ? 10'hf8 : _GEN_247; // @[RAM_ST.scala 31:71]
  assign _GEN_249 = 10'hf9 == WADDR ? 10'hf9 : _GEN_248; // @[RAM_ST.scala 31:71]
  assign _GEN_250 = 10'hfa == WADDR ? 10'hfa : _GEN_249; // @[RAM_ST.scala 31:71]
  assign _GEN_251 = 10'hfb == WADDR ? 10'hfb : _GEN_250; // @[RAM_ST.scala 31:71]
  assign _GEN_252 = 10'hfc == WADDR ? 10'hfc : _GEN_251; // @[RAM_ST.scala 31:71]
  assign _GEN_253 = 10'hfd == WADDR ? 10'hfd : _GEN_252; // @[RAM_ST.scala 31:71]
  assign _GEN_254 = 10'hfe == WADDR ? 10'hfe : _GEN_253; // @[RAM_ST.scala 31:71]
  assign _GEN_255 = 10'hff == WADDR ? 10'hff : _GEN_254; // @[RAM_ST.scala 31:71]
  assign _GEN_256 = 10'h100 == WADDR ? 10'h100 : _GEN_255; // @[RAM_ST.scala 31:71]
  assign _GEN_257 = 10'h101 == WADDR ? 10'h101 : _GEN_256; // @[RAM_ST.scala 31:71]
  assign _GEN_258 = 10'h102 == WADDR ? 10'h102 : _GEN_257; // @[RAM_ST.scala 31:71]
  assign _GEN_259 = 10'h103 == WADDR ? 10'h103 : _GEN_258; // @[RAM_ST.scala 31:71]
  assign _GEN_260 = 10'h104 == WADDR ? 10'h104 : _GEN_259; // @[RAM_ST.scala 31:71]
  assign _GEN_261 = 10'h105 == WADDR ? 10'h105 : _GEN_260; // @[RAM_ST.scala 31:71]
  assign _GEN_262 = 10'h106 == WADDR ? 10'h106 : _GEN_261; // @[RAM_ST.scala 31:71]
  assign _GEN_263 = 10'h107 == WADDR ? 10'h107 : _GEN_262; // @[RAM_ST.scala 31:71]
  assign _GEN_264 = 10'h108 == WADDR ? 10'h108 : _GEN_263; // @[RAM_ST.scala 31:71]
  assign _GEN_265 = 10'h109 == WADDR ? 10'h109 : _GEN_264; // @[RAM_ST.scala 31:71]
  assign _GEN_266 = 10'h10a == WADDR ? 10'h10a : _GEN_265; // @[RAM_ST.scala 31:71]
  assign _GEN_267 = 10'h10b == WADDR ? 10'h10b : _GEN_266; // @[RAM_ST.scala 31:71]
  assign _GEN_268 = 10'h10c == WADDR ? 10'h10c : _GEN_267; // @[RAM_ST.scala 31:71]
  assign _GEN_269 = 10'h10d == WADDR ? 10'h10d : _GEN_268; // @[RAM_ST.scala 31:71]
  assign _GEN_270 = 10'h10e == WADDR ? 10'h10e : _GEN_269; // @[RAM_ST.scala 31:71]
  assign _GEN_271 = 10'h10f == WADDR ? 10'h10f : _GEN_270; // @[RAM_ST.scala 31:71]
  assign _GEN_272 = 10'h110 == WADDR ? 10'h110 : _GEN_271; // @[RAM_ST.scala 31:71]
  assign _GEN_273 = 10'h111 == WADDR ? 10'h111 : _GEN_272; // @[RAM_ST.scala 31:71]
  assign _GEN_274 = 10'h112 == WADDR ? 10'h112 : _GEN_273; // @[RAM_ST.scala 31:71]
  assign _GEN_275 = 10'h113 == WADDR ? 10'h113 : _GEN_274; // @[RAM_ST.scala 31:71]
  assign _GEN_276 = 10'h114 == WADDR ? 10'h114 : _GEN_275; // @[RAM_ST.scala 31:71]
  assign _GEN_277 = 10'h115 == WADDR ? 10'h115 : _GEN_276; // @[RAM_ST.scala 31:71]
  assign _GEN_278 = 10'h116 == WADDR ? 10'h116 : _GEN_277; // @[RAM_ST.scala 31:71]
  assign _GEN_279 = 10'h117 == WADDR ? 10'h117 : _GEN_278; // @[RAM_ST.scala 31:71]
  assign _GEN_280 = 10'h118 == WADDR ? 10'h118 : _GEN_279; // @[RAM_ST.scala 31:71]
  assign _GEN_281 = 10'h119 == WADDR ? 10'h119 : _GEN_280; // @[RAM_ST.scala 31:71]
  assign _GEN_282 = 10'h11a == WADDR ? 10'h11a : _GEN_281; // @[RAM_ST.scala 31:71]
  assign _GEN_283 = 10'h11b == WADDR ? 10'h11b : _GEN_282; // @[RAM_ST.scala 31:71]
  assign _GEN_284 = 10'h11c == WADDR ? 10'h11c : _GEN_283; // @[RAM_ST.scala 31:71]
  assign _GEN_285 = 10'h11d == WADDR ? 10'h11d : _GEN_284; // @[RAM_ST.scala 31:71]
  assign _GEN_286 = 10'h11e == WADDR ? 10'h11e : _GEN_285; // @[RAM_ST.scala 31:71]
  assign _GEN_287 = 10'h11f == WADDR ? 10'h11f : _GEN_286; // @[RAM_ST.scala 31:71]
  assign _GEN_288 = 10'h120 == WADDR ? 10'h120 : _GEN_287; // @[RAM_ST.scala 31:71]
  assign _GEN_289 = 10'h121 == WADDR ? 10'h121 : _GEN_288; // @[RAM_ST.scala 31:71]
  assign _GEN_290 = 10'h122 == WADDR ? 10'h122 : _GEN_289; // @[RAM_ST.scala 31:71]
  assign _GEN_291 = 10'h123 == WADDR ? 10'h123 : _GEN_290; // @[RAM_ST.scala 31:71]
  assign _GEN_292 = 10'h124 == WADDR ? 10'h124 : _GEN_291; // @[RAM_ST.scala 31:71]
  assign _GEN_293 = 10'h125 == WADDR ? 10'h125 : _GEN_292; // @[RAM_ST.scala 31:71]
  assign _GEN_294 = 10'h126 == WADDR ? 10'h126 : _GEN_293; // @[RAM_ST.scala 31:71]
  assign _GEN_295 = 10'h127 == WADDR ? 10'h127 : _GEN_294; // @[RAM_ST.scala 31:71]
  assign _GEN_296 = 10'h128 == WADDR ? 10'h128 : _GEN_295; // @[RAM_ST.scala 31:71]
  assign _GEN_297 = 10'h129 == WADDR ? 10'h129 : _GEN_296; // @[RAM_ST.scala 31:71]
  assign _GEN_298 = 10'h12a == WADDR ? 10'h12a : _GEN_297; // @[RAM_ST.scala 31:71]
  assign _GEN_299 = 10'h12b == WADDR ? 10'h12b : _GEN_298; // @[RAM_ST.scala 31:71]
  assign _GEN_300 = 10'h12c == WADDR ? 10'h12c : _GEN_299; // @[RAM_ST.scala 31:71]
  assign _GEN_301 = 10'h12d == WADDR ? 10'h12d : _GEN_300; // @[RAM_ST.scala 31:71]
  assign _GEN_302 = 10'h12e == WADDR ? 10'h12e : _GEN_301; // @[RAM_ST.scala 31:71]
  assign _GEN_303 = 10'h12f == WADDR ? 10'h12f : _GEN_302; // @[RAM_ST.scala 31:71]
  assign _GEN_304 = 10'h130 == WADDR ? 10'h130 : _GEN_303; // @[RAM_ST.scala 31:71]
  assign _GEN_305 = 10'h131 == WADDR ? 10'h131 : _GEN_304; // @[RAM_ST.scala 31:71]
  assign _GEN_306 = 10'h132 == WADDR ? 10'h132 : _GEN_305; // @[RAM_ST.scala 31:71]
  assign _GEN_307 = 10'h133 == WADDR ? 10'h133 : _GEN_306; // @[RAM_ST.scala 31:71]
  assign _GEN_308 = 10'h134 == WADDR ? 10'h134 : _GEN_307; // @[RAM_ST.scala 31:71]
  assign _GEN_309 = 10'h135 == WADDR ? 10'h135 : _GEN_308; // @[RAM_ST.scala 31:71]
  assign _GEN_310 = 10'h136 == WADDR ? 10'h136 : _GEN_309; // @[RAM_ST.scala 31:71]
  assign _GEN_311 = 10'h137 == WADDR ? 10'h137 : _GEN_310; // @[RAM_ST.scala 31:71]
  assign _GEN_312 = 10'h138 == WADDR ? 10'h138 : _GEN_311; // @[RAM_ST.scala 31:71]
  assign _GEN_313 = 10'h139 == WADDR ? 10'h139 : _GEN_312; // @[RAM_ST.scala 31:71]
  assign _GEN_314 = 10'h13a == WADDR ? 10'h13a : _GEN_313; // @[RAM_ST.scala 31:71]
  assign _GEN_315 = 10'h13b == WADDR ? 10'h13b : _GEN_314; // @[RAM_ST.scala 31:71]
  assign _GEN_316 = 10'h13c == WADDR ? 10'h13c : _GEN_315; // @[RAM_ST.scala 31:71]
  assign _GEN_317 = 10'h13d == WADDR ? 10'h13d : _GEN_316; // @[RAM_ST.scala 31:71]
  assign _GEN_318 = 10'h13e == WADDR ? 10'h13e : _GEN_317; // @[RAM_ST.scala 31:71]
  assign _GEN_319 = 10'h13f == WADDR ? 10'h13f : _GEN_318; // @[RAM_ST.scala 31:71]
  assign _GEN_320 = 10'h140 == WADDR ? 10'h140 : _GEN_319; // @[RAM_ST.scala 31:71]
  assign _GEN_321 = 10'h141 == WADDR ? 10'h141 : _GEN_320; // @[RAM_ST.scala 31:71]
  assign _GEN_322 = 10'h142 == WADDR ? 10'h142 : _GEN_321; // @[RAM_ST.scala 31:71]
  assign _GEN_323 = 10'h143 == WADDR ? 10'h143 : _GEN_322; // @[RAM_ST.scala 31:71]
  assign _GEN_324 = 10'h144 == WADDR ? 10'h144 : _GEN_323; // @[RAM_ST.scala 31:71]
  assign _GEN_325 = 10'h145 == WADDR ? 10'h145 : _GEN_324; // @[RAM_ST.scala 31:71]
  assign _GEN_326 = 10'h146 == WADDR ? 10'h146 : _GEN_325; // @[RAM_ST.scala 31:71]
  assign _GEN_327 = 10'h147 == WADDR ? 10'h147 : _GEN_326; // @[RAM_ST.scala 31:71]
  assign _GEN_328 = 10'h148 == WADDR ? 10'h148 : _GEN_327; // @[RAM_ST.scala 31:71]
  assign _GEN_329 = 10'h149 == WADDR ? 10'h149 : _GEN_328; // @[RAM_ST.scala 31:71]
  assign _GEN_330 = 10'h14a == WADDR ? 10'h14a : _GEN_329; // @[RAM_ST.scala 31:71]
  assign _GEN_331 = 10'h14b == WADDR ? 10'h14b : _GEN_330; // @[RAM_ST.scala 31:71]
  assign _GEN_332 = 10'h14c == WADDR ? 10'h14c : _GEN_331; // @[RAM_ST.scala 31:71]
  assign _GEN_333 = 10'h14d == WADDR ? 10'h14d : _GEN_332; // @[RAM_ST.scala 31:71]
  assign _GEN_334 = 10'h14e == WADDR ? 10'h14e : _GEN_333; // @[RAM_ST.scala 31:71]
  assign _GEN_335 = 10'h14f == WADDR ? 10'h14f : _GEN_334; // @[RAM_ST.scala 31:71]
  assign _GEN_336 = 10'h150 == WADDR ? 10'h150 : _GEN_335; // @[RAM_ST.scala 31:71]
  assign _GEN_337 = 10'h151 == WADDR ? 10'h151 : _GEN_336; // @[RAM_ST.scala 31:71]
  assign _GEN_338 = 10'h152 == WADDR ? 10'h152 : _GEN_337; // @[RAM_ST.scala 31:71]
  assign _GEN_339 = 10'h153 == WADDR ? 10'h153 : _GEN_338; // @[RAM_ST.scala 31:71]
  assign _GEN_340 = 10'h154 == WADDR ? 10'h154 : _GEN_339; // @[RAM_ST.scala 31:71]
  assign _GEN_341 = 10'h155 == WADDR ? 10'h155 : _GEN_340; // @[RAM_ST.scala 31:71]
  assign _GEN_342 = 10'h156 == WADDR ? 10'h156 : _GEN_341; // @[RAM_ST.scala 31:71]
  assign _GEN_343 = 10'h157 == WADDR ? 10'h157 : _GEN_342; // @[RAM_ST.scala 31:71]
  assign _GEN_344 = 10'h158 == WADDR ? 10'h158 : _GEN_343; // @[RAM_ST.scala 31:71]
  assign _GEN_345 = 10'h159 == WADDR ? 10'h159 : _GEN_344; // @[RAM_ST.scala 31:71]
  assign _GEN_346 = 10'h15a == WADDR ? 10'h15a : _GEN_345; // @[RAM_ST.scala 31:71]
  assign _GEN_347 = 10'h15b == WADDR ? 10'h15b : _GEN_346; // @[RAM_ST.scala 31:71]
  assign _GEN_348 = 10'h15c == WADDR ? 10'h15c : _GEN_347; // @[RAM_ST.scala 31:71]
  assign _GEN_349 = 10'h15d == WADDR ? 10'h15d : _GEN_348; // @[RAM_ST.scala 31:71]
  assign _GEN_350 = 10'h15e == WADDR ? 10'h15e : _GEN_349; // @[RAM_ST.scala 31:71]
  assign _GEN_351 = 10'h15f == WADDR ? 10'h15f : _GEN_350; // @[RAM_ST.scala 31:71]
  assign _GEN_352 = 10'h160 == WADDR ? 10'h160 : _GEN_351; // @[RAM_ST.scala 31:71]
  assign _GEN_353 = 10'h161 == WADDR ? 10'h161 : _GEN_352; // @[RAM_ST.scala 31:71]
  assign _GEN_354 = 10'h162 == WADDR ? 10'h162 : _GEN_353; // @[RAM_ST.scala 31:71]
  assign _GEN_355 = 10'h163 == WADDR ? 10'h163 : _GEN_354; // @[RAM_ST.scala 31:71]
  assign _GEN_356 = 10'h164 == WADDR ? 10'h164 : _GEN_355; // @[RAM_ST.scala 31:71]
  assign _GEN_357 = 10'h165 == WADDR ? 10'h165 : _GEN_356; // @[RAM_ST.scala 31:71]
  assign _GEN_358 = 10'h166 == WADDR ? 10'h166 : _GEN_357; // @[RAM_ST.scala 31:71]
  assign _GEN_359 = 10'h167 == WADDR ? 10'h167 : _GEN_358; // @[RAM_ST.scala 31:71]
  assign _GEN_360 = 10'h168 == WADDR ? 10'h168 : _GEN_359; // @[RAM_ST.scala 31:71]
  assign _GEN_361 = 10'h169 == WADDR ? 10'h169 : _GEN_360; // @[RAM_ST.scala 31:71]
  assign _GEN_362 = 10'h16a == WADDR ? 10'h16a : _GEN_361; // @[RAM_ST.scala 31:71]
  assign _GEN_363 = 10'h16b == WADDR ? 10'h16b : _GEN_362; // @[RAM_ST.scala 31:71]
  assign _GEN_364 = 10'h16c == WADDR ? 10'h16c : _GEN_363; // @[RAM_ST.scala 31:71]
  assign _GEN_365 = 10'h16d == WADDR ? 10'h16d : _GEN_364; // @[RAM_ST.scala 31:71]
  assign _GEN_366 = 10'h16e == WADDR ? 10'h16e : _GEN_365; // @[RAM_ST.scala 31:71]
  assign _GEN_367 = 10'h16f == WADDR ? 10'h16f : _GEN_366; // @[RAM_ST.scala 31:71]
  assign _GEN_368 = 10'h170 == WADDR ? 10'h170 : _GEN_367; // @[RAM_ST.scala 31:71]
  assign _GEN_369 = 10'h171 == WADDR ? 10'h171 : _GEN_368; // @[RAM_ST.scala 31:71]
  assign _GEN_370 = 10'h172 == WADDR ? 10'h172 : _GEN_369; // @[RAM_ST.scala 31:71]
  assign _GEN_371 = 10'h173 == WADDR ? 10'h173 : _GEN_370; // @[RAM_ST.scala 31:71]
  assign _GEN_372 = 10'h174 == WADDR ? 10'h174 : _GEN_371; // @[RAM_ST.scala 31:71]
  assign _GEN_373 = 10'h175 == WADDR ? 10'h175 : _GEN_372; // @[RAM_ST.scala 31:71]
  assign _GEN_374 = 10'h176 == WADDR ? 10'h176 : _GEN_373; // @[RAM_ST.scala 31:71]
  assign _GEN_375 = 10'h177 == WADDR ? 10'h177 : _GEN_374; // @[RAM_ST.scala 31:71]
  assign _GEN_376 = 10'h178 == WADDR ? 10'h178 : _GEN_375; // @[RAM_ST.scala 31:71]
  assign _GEN_377 = 10'h179 == WADDR ? 10'h179 : _GEN_376; // @[RAM_ST.scala 31:71]
  assign _GEN_378 = 10'h17a == WADDR ? 10'h17a : _GEN_377; // @[RAM_ST.scala 31:71]
  assign _GEN_379 = 10'h17b == WADDR ? 10'h17b : _GEN_378; // @[RAM_ST.scala 31:71]
  assign _GEN_380 = 10'h17c == WADDR ? 10'h17c : _GEN_379; // @[RAM_ST.scala 31:71]
  assign _GEN_381 = 10'h17d == WADDR ? 10'h17d : _GEN_380; // @[RAM_ST.scala 31:71]
  assign _GEN_382 = 10'h17e == WADDR ? 10'h17e : _GEN_381; // @[RAM_ST.scala 31:71]
  assign _GEN_383 = 10'h17f == WADDR ? 10'h17f : _GEN_382; // @[RAM_ST.scala 31:71]
  assign _GEN_384 = 10'h180 == WADDR ? 10'h180 : _GEN_383; // @[RAM_ST.scala 31:71]
  assign _GEN_385 = 10'h181 == WADDR ? 10'h181 : _GEN_384; // @[RAM_ST.scala 31:71]
  assign _GEN_386 = 10'h182 == WADDR ? 10'h182 : _GEN_385; // @[RAM_ST.scala 31:71]
  assign _GEN_387 = 10'h183 == WADDR ? 10'h183 : _GEN_386; // @[RAM_ST.scala 31:71]
  assign _GEN_388 = 10'h184 == WADDR ? 10'h184 : _GEN_387; // @[RAM_ST.scala 31:71]
  assign _GEN_389 = 10'h185 == WADDR ? 10'h185 : _GEN_388; // @[RAM_ST.scala 31:71]
  assign _GEN_390 = 10'h186 == WADDR ? 10'h186 : _GEN_389; // @[RAM_ST.scala 31:71]
  assign _GEN_391 = 10'h187 == WADDR ? 10'h187 : _GEN_390; // @[RAM_ST.scala 31:71]
  assign _GEN_392 = 10'h188 == WADDR ? 10'h188 : _GEN_391; // @[RAM_ST.scala 31:71]
  assign _GEN_393 = 10'h189 == WADDR ? 10'h189 : _GEN_392; // @[RAM_ST.scala 31:71]
  assign _GEN_394 = 10'h18a == WADDR ? 10'h18a : _GEN_393; // @[RAM_ST.scala 31:71]
  assign _GEN_395 = 10'h18b == WADDR ? 10'h18b : _GEN_394; // @[RAM_ST.scala 31:71]
  assign _GEN_396 = 10'h18c == WADDR ? 10'h18c : _GEN_395; // @[RAM_ST.scala 31:71]
  assign _GEN_397 = 10'h18d == WADDR ? 10'h18d : _GEN_396; // @[RAM_ST.scala 31:71]
  assign _GEN_398 = 10'h18e == WADDR ? 10'h18e : _GEN_397; // @[RAM_ST.scala 31:71]
  assign _GEN_399 = 10'h18f == WADDR ? 10'h18f : _GEN_398; // @[RAM_ST.scala 31:71]
  assign _GEN_400 = 10'h190 == WADDR ? 10'h190 : _GEN_399; // @[RAM_ST.scala 31:71]
  assign _GEN_401 = 10'h191 == WADDR ? 10'h191 : _GEN_400; // @[RAM_ST.scala 31:71]
  assign _GEN_402 = 10'h192 == WADDR ? 10'h192 : _GEN_401; // @[RAM_ST.scala 31:71]
  assign _GEN_403 = 10'h193 == WADDR ? 10'h193 : _GEN_402; // @[RAM_ST.scala 31:71]
  assign _GEN_404 = 10'h194 == WADDR ? 10'h194 : _GEN_403; // @[RAM_ST.scala 31:71]
  assign _GEN_405 = 10'h195 == WADDR ? 10'h195 : _GEN_404; // @[RAM_ST.scala 31:71]
  assign _GEN_406 = 10'h196 == WADDR ? 10'h196 : _GEN_405; // @[RAM_ST.scala 31:71]
  assign _GEN_407 = 10'h197 == WADDR ? 10'h197 : _GEN_406; // @[RAM_ST.scala 31:71]
  assign _GEN_408 = 10'h198 == WADDR ? 10'h198 : _GEN_407; // @[RAM_ST.scala 31:71]
  assign _GEN_409 = 10'h199 == WADDR ? 10'h199 : _GEN_408; // @[RAM_ST.scala 31:71]
  assign _GEN_410 = 10'h19a == WADDR ? 10'h19a : _GEN_409; // @[RAM_ST.scala 31:71]
  assign _GEN_411 = 10'h19b == WADDR ? 10'h19b : _GEN_410; // @[RAM_ST.scala 31:71]
  assign _GEN_412 = 10'h19c == WADDR ? 10'h19c : _GEN_411; // @[RAM_ST.scala 31:71]
  assign _GEN_413 = 10'h19d == WADDR ? 10'h19d : _GEN_412; // @[RAM_ST.scala 31:71]
  assign _GEN_414 = 10'h19e == WADDR ? 10'h19e : _GEN_413; // @[RAM_ST.scala 31:71]
  assign _GEN_415 = 10'h19f == WADDR ? 10'h19f : _GEN_414; // @[RAM_ST.scala 31:71]
  assign _GEN_416 = 10'h1a0 == WADDR ? 10'h1a0 : _GEN_415; // @[RAM_ST.scala 31:71]
  assign _GEN_417 = 10'h1a1 == WADDR ? 10'h1a1 : _GEN_416; // @[RAM_ST.scala 31:71]
  assign _GEN_418 = 10'h1a2 == WADDR ? 10'h1a2 : _GEN_417; // @[RAM_ST.scala 31:71]
  assign _GEN_419 = 10'h1a3 == WADDR ? 10'h1a3 : _GEN_418; // @[RAM_ST.scala 31:71]
  assign _GEN_420 = 10'h1a4 == WADDR ? 10'h1a4 : _GEN_419; // @[RAM_ST.scala 31:71]
  assign _GEN_421 = 10'h1a5 == WADDR ? 10'h1a5 : _GEN_420; // @[RAM_ST.scala 31:71]
  assign _GEN_422 = 10'h1a6 == WADDR ? 10'h1a6 : _GEN_421; // @[RAM_ST.scala 31:71]
  assign _GEN_423 = 10'h1a7 == WADDR ? 10'h1a7 : _GEN_422; // @[RAM_ST.scala 31:71]
  assign _GEN_424 = 10'h1a8 == WADDR ? 10'h1a8 : _GEN_423; // @[RAM_ST.scala 31:71]
  assign _GEN_425 = 10'h1a9 == WADDR ? 10'h1a9 : _GEN_424; // @[RAM_ST.scala 31:71]
  assign _GEN_426 = 10'h1aa == WADDR ? 10'h1aa : _GEN_425; // @[RAM_ST.scala 31:71]
  assign _GEN_427 = 10'h1ab == WADDR ? 10'h1ab : _GEN_426; // @[RAM_ST.scala 31:71]
  assign _GEN_428 = 10'h1ac == WADDR ? 10'h1ac : _GEN_427; // @[RAM_ST.scala 31:71]
  assign _GEN_429 = 10'h1ad == WADDR ? 10'h1ad : _GEN_428; // @[RAM_ST.scala 31:71]
  assign _GEN_430 = 10'h1ae == WADDR ? 10'h1ae : _GEN_429; // @[RAM_ST.scala 31:71]
  assign _GEN_431 = 10'h1af == WADDR ? 10'h1af : _GEN_430; // @[RAM_ST.scala 31:71]
  assign _GEN_432 = 10'h1b0 == WADDR ? 10'h1b0 : _GEN_431; // @[RAM_ST.scala 31:71]
  assign _GEN_433 = 10'h1b1 == WADDR ? 10'h1b1 : _GEN_432; // @[RAM_ST.scala 31:71]
  assign _GEN_434 = 10'h1b2 == WADDR ? 10'h1b2 : _GEN_433; // @[RAM_ST.scala 31:71]
  assign _GEN_435 = 10'h1b3 == WADDR ? 10'h1b3 : _GEN_434; // @[RAM_ST.scala 31:71]
  assign _GEN_436 = 10'h1b4 == WADDR ? 10'h1b4 : _GEN_435; // @[RAM_ST.scala 31:71]
  assign _GEN_437 = 10'h1b5 == WADDR ? 10'h1b5 : _GEN_436; // @[RAM_ST.scala 31:71]
  assign _GEN_438 = 10'h1b6 == WADDR ? 10'h1b6 : _GEN_437; // @[RAM_ST.scala 31:71]
  assign _GEN_439 = 10'h1b7 == WADDR ? 10'h1b7 : _GEN_438; // @[RAM_ST.scala 31:71]
  assign _GEN_440 = 10'h1b8 == WADDR ? 10'h1b8 : _GEN_439; // @[RAM_ST.scala 31:71]
  assign _GEN_441 = 10'h1b9 == WADDR ? 10'h1b9 : _GEN_440; // @[RAM_ST.scala 31:71]
  assign _GEN_442 = 10'h1ba == WADDR ? 10'h1ba : _GEN_441; // @[RAM_ST.scala 31:71]
  assign _GEN_443 = 10'h1bb == WADDR ? 10'h1bb : _GEN_442; // @[RAM_ST.scala 31:71]
  assign _GEN_444 = 10'h1bc == WADDR ? 10'h1bc : _GEN_443; // @[RAM_ST.scala 31:71]
  assign _GEN_445 = 10'h1bd == WADDR ? 10'h1bd : _GEN_444; // @[RAM_ST.scala 31:71]
  assign _GEN_446 = 10'h1be == WADDR ? 10'h1be : _GEN_445; // @[RAM_ST.scala 31:71]
  assign _GEN_447 = 10'h1bf == WADDR ? 10'h1bf : _GEN_446; // @[RAM_ST.scala 31:71]
  assign _GEN_448 = 10'h1c0 == WADDR ? 10'h1c0 : _GEN_447; // @[RAM_ST.scala 31:71]
  assign _GEN_449 = 10'h1c1 == WADDR ? 10'h1c1 : _GEN_448; // @[RAM_ST.scala 31:71]
  assign _GEN_450 = 10'h1c2 == WADDR ? 10'h1c2 : _GEN_449; // @[RAM_ST.scala 31:71]
  assign _GEN_451 = 10'h1c3 == WADDR ? 10'h1c3 : _GEN_450; // @[RAM_ST.scala 31:71]
  assign _GEN_452 = 10'h1c4 == WADDR ? 10'h1c4 : _GEN_451; // @[RAM_ST.scala 31:71]
  assign _GEN_453 = 10'h1c5 == WADDR ? 10'h1c5 : _GEN_452; // @[RAM_ST.scala 31:71]
  assign _GEN_454 = 10'h1c6 == WADDR ? 10'h1c6 : _GEN_453; // @[RAM_ST.scala 31:71]
  assign _GEN_455 = 10'h1c7 == WADDR ? 10'h1c7 : _GEN_454; // @[RAM_ST.scala 31:71]
  assign _GEN_456 = 10'h1c8 == WADDR ? 10'h1c8 : _GEN_455; // @[RAM_ST.scala 31:71]
  assign _GEN_457 = 10'h1c9 == WADDR ? 10'h1c9 : _GEN_456; // @[RAM_ST.scala 31:71]
  assign _GEN_458 = 10'h1ca == WADDR ? 10'h1ca : _GEN_457; // @[RAM_ST.scala 31:71]
  assign _GEN_459 = 10'h1cb == WADDR ? 10'h1cb : _GEN_458; // @[RAM_ST.scala 31:71]
  assign _GEN_460 = 10'h1cc == WADDR ? 10'h1cc : _GEN_459; // @[RAM_ST.scala 31:71]
  assign _GEN_461 = 10'h1cd == WADDR ? 10'h1cd : _GEN_460; // @[RAM_ST.scala 31:71]
  assign _GEN_462 = 10'h1ce == WADDR ? 10'h1ce : _GEN_461; // @[RAM_ST.scala 31:71]
  assign _GEN_463 = 10'h1cf == WADDR ? 10'h1cf : _GEN_462; // @[RAM_ST.scala 31:71]
  assign _GEN_464 = 10'h1d0 == WADDR ? 10'h1d0 : _GEN_463; // @[RAM_ST.scala 31:71]
  assign _GEN_465 = 10'h1d1 == WADDR ? 10'h1d1 : _GEN_464; // @[RAM_ST.scala 31:71]
  assign _GEN_466 = 10'h1d2 == WADDR ? 10'h1d2 : _GEN_465; // @[RAM_ST.scala 31:71]
  assign _GEN_467 = 10'h1d3 == WADDR ? 10'h1d3 : _GEN_466; // @[RAM_ST.scala 31:71]
  assign _GEN_468 = 10'h1d4 == WADDR ? 10'h1d4 : _GEN_467; // @[RAM_ST.scala 31:71]
  assign _GEN_469 = 10'h1d5 == WADDR ? 10'h1d5 : _GEN_468; // @[RAM_ST.scala 31:71]
  assign _GEN_470 = 10'h1d6 == WADDR ? 10'h1d6 : _GEN_469; // @[RAM_ST.scala 31:71]
  assign _GEN_471 = 10'h1d7 == WADDR ? 10'h1d7 : _GEN_470; // @[RAM_ST.scala 31:71]
  assign _GEN_472 = 10'h1d8 == WADDR ? 10'h1d8 : _GEN_471; // @[RAM_ST.scala 31:71]
  assign _GEN_473 = 10'h1d9 == WADDR ? 10'h1d9 : _GEN_472; // @[RAM_ST.scala 31:71]
  assign _GEN_474 = 10'h1da == WADDR ? 10'h1da : _GEN_473; // @[RAM_ST.scala 31:71]
  assign _GEN_475 = 10'h1db == WADDR ? 10'h1db : _GEN_474; // @[RAM_ST.scala 31:71]
  assign _GEN_476 = 10'h1dc == WADDR ? 10'h1dc : _GEN_475; // @[RAM_ST.scala 31:71]
  assign _GEN_477 = 10'h1dd == WADDR ? 10'h1dd : _GEN_476; // @[RAM_ST.scala 31:71]
  assign _GEN_478 = 10'h1de == WADDR ? 10'h1de : _GEN_477; // @[RAM_ST.scala 31:71]
  assign _GEN_479 = 10'h1df == WADDR ? 10'h1df : _GEN_478; // @[RAM_ST.scala 31:71]
  assign _GEN_480 = 10'h1e0 == WADDR ? 10'h1e0 : _GEN_479; // @[RAM_ST.scala 31:71]
  assign _GEN_481 = 10'h1e1 == WADDR ? 10'h1e1 : _GEN_480; // @[RAM_ST.scala 31:71]
  assign _GEN_482 = 10'h1e2 == WADDR ? 10'h1e2 : _GEN_481; // @[RAM_ST.scala 31:71]
  assign _GEN_483 = 10'h1e3 == WADDR ? 10'h1e3 : _GEN_482; // @[RAM_ST.scala 31:71]
  assign _GEN_484 = 10'h1e4 == WADDR ? 10'h1e4 : _GEN_483; // @[RAM_ST.scala 31:71]
  assign _GEN_485 = 10'h1e5 == WADDR ? 10'h1e5 : _GEN_484; // @[RAM_ST.scala 31:71]
  assign _GEN_486 = 10'h1e6 == WADDR ? 10'h1e6 : _GEN_485; // @[RAM_ST.scala 31:71]
  assign _GEN_487 = 10'h1e7 == WADDR ? 10'h1e7 : _GEN_486; // @[RAM_ST.scala 31:71]
  assign _GEN_488 = 10'h1e8 == WADDR ? 10'h1e8 : _GEN_487; // @[RAM_ST.scala 31:71]
  assign _GEN_489 = 10'h1e9 == WADDR ? 10'h1e9 : _GEN_488; // @[RAM_ST.scala 31:71]
  assign _GEN_490 = 10'h1ea == WADDR ? 10'h1ea : _GEN_489; // @[RAM_ST.scala 31:71]
  assign _GEN_491 = 10'h1eb == WADDR ? 10'h1eb : _GEN_490; // @[RAM_ST.scala 31:71]
  assign _GEN_492 = 10'h1ec == WADDR ? 10'h1ec : _GEN_491; // @[RAM_ST.scala 31:71]
  assign _GEN_493 = 10'h1ed == WADDR ? 10'h1ed : _GEN_492; // @[RAM_ST.scala 31:71]
  assign _GEN_494 = 10'h1ee == WADDR ? 10'h1ee : _GEN_493; // @[RAM_ST.scala 31:71]
  assign _GEN_495 = 10'h1ef == WADDR ? 10'h1ef : _GEN_494; // @[RAM_ST.scala 31:71]
  assign _GEN_496 = 10'h1f0 == WADDR ? 10'h1f0 : _GEN_495; // @[RAM_ST.scala 31:71]
  assign _GEN_497 = 10'h1f1 == WADDR ? 10'h1f1 : _GEN_496; // @[RAM_ST.scala 31:71]
  assign _GEN_498 = 10'h1f2 == WADDR ? 10'h1f2 : _GEN_497; // @[RAM_ST.scala 31:71]
  assign _GEN_499 = 10'h1f3 == WADDR ? 10'h1f3 : _GEN_498; // @[RAM_ST.scala 31:71]
  assign _GEN_500 = 10'h1f4 == WADDR ? 10'h1f4 : _GEN_499; // @[RAM_ST.scala 31:71]
  assign _GEN_501 = 10'h1f5 == WADDR ? 10'h1f5 : _GEN_500; // @[RAM_ST.scala 31:71]
  assign _GEN_502 = 10'h1f6 == WADDR ? 10'h1f6 : _GEN_501; // @[RAM_ST.scala 31:71]
  assign _GEN_503 = 10'h1f7 == WADDR ? 10'h1f7 : _GEN_502; // @[RAM_ST.scala 31:71]
  assign _GEN_504 = 10'h1f8 == WADDR ? 10'h1f8 : _GEN_503; // @[RAM_ST.scala 31:71]
  assign _GEN_505 = 10'h1f9 == WADDR ? 10'h1f9 : _GEN_504; // @[RAM_ST.scala 31:71]
  assign _GEN_506 = 10'h1fa == WADDR ? 10'h1fa : _GEN_505; // @[RAM_ST.scala 31:71]
  assign _GEN_507 = 10'h1fb == WADDR ? 10'h1fb : _GEN_506; // @[RAM_ST.scala 31:71]
  assign _GEN_508 = 10'h1fc == WADDR ? 10'h1fc : _GEN_507; // @[RAM_ST.scala 31:71]
  assign _GEN_509 = 10'h1fd == WADDR ? 10'h1fd : _GEN_508; // @[RAM_ST.scala 31:71]
  assign _GEN_510 = 10'h1fe == WADDR ? 10'h1fe : _GEN_509; // @[RAM_ST.scala 31:71]
  assign _GEN_511 = 10'h1ff == WADDR ? 10'h1ff : _GEN_510; // @[RAM_ST.scala 31:71]
  assign _GEN_512 = 10'h200 == WADDR ? 10'h200 : _GEN_511; // @[RAM_ST.scala 31:71]
  assign _GEN_513 = 10'h201 == WADDR ? 10'h201 : _GEN_512; // @[RAM_ST.scala 31:71]
  assign _GEN_514 = 10'h202 == WADDR ? 10'h202 : _GEN_513; // @[RAM_ST.scala 31:71]
  assign _GEN_515 = 10'h203 == WADDR ? 10'h203 : _GEN_514; // @[RAM_ST.scala 31:71]
  assign _GEN_516 = 10'h204 == WADDR ? 10'h204 : _GEN_515; // @[RAM_ST.scala 31:71]
  assign _GEN_517 = 10'h205 == WADDR ? 10'h205 : _GEN_516; // @[RAM_ST.scala 31:71]
  assign _GEN_518 = 10'h206 == WADDR ? 10'h206 : _GEN_517; // @[RAM_ST.scala 31:71]
  assign _GEN_519 = 10'h207 == WADDR ? 10'h207 : _GEN_518; // @[RAM_ST.scala 31:71]
  assign _GEN_520 = 10'h208 == WADDR ? 10'h208 : _GEN_519; // @[RAM_ST.scala 31:71]
  assign _GEN_521 = 10'h209 == WADDR ? 10'h209 : _GEN_520; // @[RAM_ST.scala 31:71]
  assign _GEN_522 = 10'h20a == WADDR ? 10'h20a : _GEN_521; // @[RAM_ST.scala 31:71]
  assign _GEN_523 = 10'h20b == WADDR ? 10'h20b : _GEN_522; // @[RAM_ST.scala 31:71]
  assign _GEN_524 = 10'h20c == WADDR ? 10'h20c : _GEN_523; // @[RAM_ST.scala 31:71]
  assign _GEN_525 = 10'h20d == WADDR ? 10'h20d : _GEN_524; // @[RAM_ST.scala 31:71]
  assign _GEN_526 = 10'h20e == WADDR ? 10'h20e : _GEN_525; // @[RAM_ST.scala 31:71]
  assign _GEN_527 = 10'h20f == WADDR ? 10'h20f : _GEN_526; // @[RAM_ST.scala 31:71]
  assign _GEN_528 = 10'h210 == WADDR ? 10'h210 : _GEN_527; // @[RAM_ST.scala 31:71]
  assign _GEN_529 = 10'h211 == WADDR ? 10'h211 : _GEN_528; // @[RAM_ST.scala 31:71]
  assign _GEN_530 = 10'h212 == WADDR ? 10'h212 : _GEN_529; // @[RAM_ST.scala 31:71]
  assign _GEN_531 = 10'h213 == WADDR ? 10'h213 : _GEN_530; // @[RAM_ST.scala 31:71]
  assign _GEN_532 = 10'h214 == WADDR ? 10'h214 : _GEN_531; // @[RAM_ST.scala 31:71]
  assign _GEN_533 = 10'h215 == WADDR ? 10'h215 : _GEN_532; // @[RAM_ST.scala 31:71]
  assign _GEN_534 = 10'h216 == WADDR ? 10'h216 : _GEN_533; // @[RAM_ST.scala 31:71]
  assign _GEN_535 = 10'h217 == WADDR ? 10'h217 : _GEN_534; // @[RAM_ST.scala 31:71]
  assign _GEN_536 = 10'h218 == WADDR ? 10'h218 : _GEN_535; // @[RAM_ST.scala 31:71]
  assign _GEN_537 = 10'h219 == WADDR ? 10'h219 : _GEN_536; // @[RAM_ST.scala 31:71]
  assign _GEN_538 = 10'h21a == WADDR ? 10'h21a : _GEN_537; // @[RAM_ST.scala 31:71]
  assign _GEN_539 = 10'h21b == WADDR ? 10'h21b : _GEN_538; // @[RAM_ST.scala 31:71]
  assign _GEN_540 = 10'h21c == WADDR ? 10'h21c : _GEN_539; // @[RAM_ST.scala 31:71]
  assign _GEN_541 = 10'h21d == WADDR ? 10'h21d : _GEN_540; // @[RAM_ST.scala 31:71]
  assign _GEN_542 = 10'h21e == WADDR ? 10'h21e : _GEN_541; // @[RAM_ST.scala 31:71]
  assign _GEN_543 = 10'h21f == WADDR ? 10'h21f : _GEN_542; // @[RAM_ST.scala 31:71]
  assign _GEN_544 = 10'h220 == WADDR ? 10'h220 : _GEN_543; // @[RAM_ST.scala 31:71]
  assign _GEN_545 = 10'h221 == WADDR ? 10'h221 : _GEN_544; // @[RAM_ST.scala 31:71]
  assign _GEN_546 = 10'h222 == WADDR ? 10'h222 : _GEN_545; // @[RAM_ST.scala 31:71]
  assign _GEN_547 = 10'h223 == WADDR ? 10'h223 : _GEN_546; // @[RAM_ST.scala 31:71]
  assign _GEN_548 = 10'h224 == WADDR ? 10'h224 : _GEN_547; // @[RAM_ST.scala 31:71]
  assign _GEN_549 = 10'h225 == WADDR ? 10'h225 : _GEN_548; // @[RAM_ST.scala 31:71]
  assign _GEN_550 = 10'h226 == WADDR ? 10'h226 : _GEN_549; // @[RAM_ST.scala 31:71]
  assign _GEN_551 = 10'h227 == WADDR ? 10'h227 : _GEN_550; // @[RAM_ST.scala 31:71]
  assign _GEN_552 = 10'h228 == WADDR ? 10'h228 : _GEN_551; // @[RAM_ST.scala 31:71]
  assign _GEN_553 = 10'h229 == WADDR ? 10'h229 : _GEN_552; // @[RAM_ST.scala 31:71]
  assign _GEN_554 = 10'h22a == WADDR ? 10'h22a : _GEN_553; // @[RAM_ST.scala 31:71]
  assign _GEN_555 = 10'h22b == WADDR ? 10'h22b : _GEN_554; // @[RAM_ST.scala 31:71]
  assign _GEN_556 = 10'h22c == WADDR ? 10'h22c : _GEN_555; // @[RAM_ST.scala 31:71]
  assign _GEN_557 = 10'h22d == WADDR ? 10'h22d : _GEN_556; // @[RAM_ST.scala 31:71]
  assign _GEN_558 = 10'h22e == WADDR ? 10'h22e : _GEN_557; // @[RAM_ST.scala 31:71]
  assign _GEN_559 = 10'h22f == WADDR ? 10'h22f : _GEN_558; // @[RAM_ST.scala 31:71]
  assign _GEN_560 = 10'h230 == WADDR ? 10'h230 : _GEN_559; // @[RAM_ST.scala 31:71]
  assign _GEN_561 = 10'h231 == WADDR ? 10'h231 : _GEN_560; // @[RAM_ST.scala 31:71]
  assign _GEN_562 = 10'h232 == WADDR ? 10'h232 : _GEN_561; // @[RAM_ST.scala 31:71]
  assign _GEN_563 = 10'h233 == WADDR ? 10'h233 : _GEN_562; // @[RAM_ST.scala 31:71]
  assign _GEN_564 = 10'h234 == WADDR ? 10'h234 : _GEN_563; // @[RAM_ST.scala 31:71]
  assign _GEN_565 = 10'h235 == WADDR ? 10'h235 : _GEN_564; // @[RAM_ST.scala 31:71]
  assign _GEN_566 = 10'h236 == WADDR ? 10'h236 : _GEN_565; // @[RAM_ST.scala 31:71]
  assign _GEN_567 = 10'h237 == WADDR ? 10'h237 : _GEN_566; // @[RAM_ST.scala 31:71]
  assign _GEN_568 = 10'h238 == WADDR ? 10'h238 : _GEN_567; // @[RAM_ST.scala 31:71]
  assign _GEN_569 = 10'h239 == WADDR ? 10'h239 : _GEN_568; // @[RAM_ST.scala 31:71]
  assign _GEN_570 = 10'h23a == WADDR ? 10'h23a : _GEN_569; // @[RAM_ST.scala 31:71]
  assign _GEN_571 = 10'h23b == WADDR ? 10'h23b : _GEN_570; // @[RAM_ST.scala 31:71]
  assign _GEN_572 = 10'h23c == WADDR ? 10'h23c : _GEN_571; // @[RAM_ST.scala 31:71]
  assign _GEN_573 = 10'h23d == WADDR ? 10'h23d : _GEN_572; // @[RAM_ST.scala 31:71]
  assign _GEN_574 = 10'h23e == WADDR ? 10'h23e : _GEN_573; // @[RAM_ST.scala 31:71]
  assign _GEN_575 = 10'h23f == WADDR ? 10'h23f : _GEN_574; // @[RAM_ST.scala 31:71]
  assign _GEN_576 = 10'h240 == WADDR ? 10'h240 : _GEN_575; // @[RAM_ST.scala 31:71]
  assign _GEN_577 = 10'h241 == WADDR ? 10'h241 : _GEN_576; // @[RAM_ST.scala 31:71]
  assign _GEN_578 = 10'h242 == WADDR ? 10'h242 : _GEN_577; // @[RAM_ST.scala 31:71]
  assign _GEN_579 = 10'h243 == WADDR ? 10'h243 : _GEN_578; // @[RAM_ST.scala 31:71]
  assign _GEN_580 = 10'h244 == WADDR ? 10'h244 : _GEN_579; // @[RAM_ST.scala 31:71]
  assign _GEN_581 = 10'h245 == WADDR ? 10'h245 : _GEN_580; // @[RAM_ST.scala 31:71]
  assign _GEN_582 = 10'h246 == WADDR ? 10'h246 : _GEN_581; // @[RAM_ST.scala 31:71]
  assign _GEN_583 = 10'h247 == WADDR ? 10'h247 : _GEN_582; // @[RAM_ST.scala 31:71]
  assign _GEN_584 = 10'h248 == WADDR ? 10'h248 : _GEN_583; // @[RAM_ST.scala 31:71]
  assign _GEN_585 = 10'h249 == WADDR ? 10'h249 : _GEN_584; // @[RAM_ST.scala 31:71]
  assign _GEN_586 = 10'h24a == WADDR ? 10'h24a : _GEN_585; // @[RAM_ST.scala 31:71]
  assign _GEN_587 = 10'h24b == WADDR ? 10'h24b : _GEN_586; // @[RAM_ST.scala 31:71]
  assign _GEN_588 = 10'h24c == WADDR ? 10'h24c : _GEN_587; // @[RAM_ST.scala 31:71]
  assign _GEN_589 = 10'h24d == WADDR ? 10'h24d : _GEN_588; // @[RAM_ST.scala 31:71]
  assign _GEN_590 = 10'h24e == WADDR ? 10'h24e : _GEN_589; // @[RAM_ST.scala 31:71]
  assign _GEN_591 = 10'h24f == WADDR ? 10'h24f : _GEN_590; // @[RAM_ST.scala 31:71]
  assign _GEN_592 = 10'h250 == WADDR ? 10'h250 : _GEN_591; // @[RAM_ST.scala 31:71]
  assign _GEN_593 = 10'h251 == WADDR ? 10'h251 : _GEN_592; // @[RAM_ST.scala 31:71]
  assign _GEN_594 = 10'h252 == WADDR ? 10'h252 : _GEN_593; // @[RAM_ST.scala 31:71]
  assign _GEN_595 = 10'h253 == WADDR ? 10'h253 : _GEN_594; // @[RAM_ST.scala 31:71]
  assign _GEN_596 = 10'h254 == WADDR ? 10'h254 : _GEN_595; // @[RAM_ST.scala 31:71]
  assign _GEN_597 = 10'h255 == WADDR ? 10'h255 : _GEN_596; // @[RAM_ST.scala 31:71]
  assign _GEN_598 = 10'h256 == WADDR ? 10'h256 : _GEN_597; // @[RAM_ST.scala 31:71]
  assign _GEN_599 = 10'h257 == WADDR ? 10'h257 : _GEN_598; // @[RAM_ST.scala 31:71]
  assign _GEN_600 = 10'h258 == WADDR ? 10'h258 : _GEN_599; // @[RAM_ST.scala 31:71]
  assign _GEN_601 = 10'h259 == WADDR ? 10'h259 : _GEN_600; // @[RAM_ST.scala 31:71]
  assign _GEN_602 = 10'h25a == WADDR ? 10'h25a : _GEN_601; // @[RAM_ST.scala 31:71]
  assign _GEN_603 = 10'h25b == WADDR ? 10'h25b : _GEN_602; // @[RAM_ST.scala 31:71]
  assign _GEN_604 = 10'h25c == WADDR ? 10'h25c : _GEN_603; // @[RAM_ST.scala 31:71]
  assign _GEN_605 = 10'h25d == WADDR ? 10'h25d : _GEN_604; // @[RAM_ST.scala 31:71]
  assign _GEN_606 = 10'h25e == WADDR ? 10'h25e : _GEN_605; // @[RAM_ST.scala 31:71]
  assign _GEN_607 = 10'h25f == WADDR ? 10'h25f : _GEN_606; // @[RAM_ST.scala 31:71]
  assign _GEN_608 = 10'h260 == WADDR ? 10'h260 : _GEN_607; // @[RAM_ST.scala 31:71]
  assign _GEN_609 = 10'h261 == WADDR ? 10'h261 : _GEN_608; // @[RAM_ST.scala 31:71]
  assign _GEN_610 = 10'h262 == WADDR ? 10'h262 : _GEN_609; // @[RAM_ST.scala 31:71]
  assign _GEN_611 = 10'h263 == WADDR ? 10'h263 : _GEN_610; // @[RAM_ST.scala 31:71]
  assign _GEN_612 = 10'h264 == WADDR ? 10'h264 : _GEN_611; // @[RAM_ST.scala 31:71]
  assign _GEN_613 = 10'h265 == WADDR ? 10'h265 : _GEN_612; // @[RAM_ST.scala 31:71]
  assign _GEN_614 = 10'h266 == WADDR ? 10'h266 : _GEN_613; // @[RAM_ST.scala 31:71]
  assign _GEN_615 = 10'h267 == WADDR ? 10'h267 : _GEN_614; // @[RAM_ST.scala 31:71]
  assign _GEN_616 = 10'h268 == WADDR ? 10'h268 : _GEN_615; // @[RAM_ST.scala 31:71]
  assign _GEN_617 = 10'h269 == WADDR ? 10'h269 : _GEN_616; // @[RAM_ST.scala 31:71]
  assign _GEN_618 = 10'h26a == WADDR ? 10'h26a : _GEN_617; // @[RAM_ST.scala 31:71]
  assign _GEN_619 = 10'h26b == WADDR ? 10'h26b : _GEN_618; // @[RAM_ST.scala 31:71]
  assign _GEN_620 = 10'h26c == WADDR ? 10'h26c : _GEN_619; // @[RAM_ST.scala 31:71]
  assign _GEN_621 = 10'h26d == WADDR ? 10'h26d : _GEN_620; // @[RAM_ST.scala 31:71]
  assign _GEN_622 = 10'h26e == WADDR ? 10'h26e : _GEN_621; // @[RAM_ST.scala 31:71]
  assign _GEN_623 = 10'h26f == WADDR ? 10'h26f : _GEN_622; // @[RAM_ST.scala 31:71]
  assign _GEN_624 = 10'h270 == WADDR ? 10'h270 : _GEN_623; // @[RAM_ST.scala 31:71]
  assign _GEN_625 = 10'h271 == WADDR ? 10'h271 : _GEN_624; // @[RAM_ST.scala 31:71]
  assign _GEN_626 = 10'h272 == WADDR ? 10'h272 : _GEN_625; // @[RAM_ST.scala 31:71]
  assign _GEN_627 = 10'h273 == WADDR ? 10'h273 : _GEN_626; // @[RAM_ST.scala 31:71]
  assign _GEN_628 = 10'h274 == WADDR ? 10'h274 : _GEN_627; // @[RAM_ST.scala 31:71]
  assign _GEN_629 = 10'h275 == WADDR ? 10'h275 : _GEN_628; // @[RAM_ST.scala 31:71]
  assign _GEN_630 = 10'h276 == WADDR ? 10'h276 : _GEN_629; // @[RAM_ST.scala 31:71]
  assign _GEN_631 = 10'h277 == WADDR ? 10'h277 : _GEN_630; // @[RAM_ST.scala 31:71]
  assign _GEN_632 = 10'h278 == WADDR ? 10'h278 : _GEN_631; // @[RAM_ST.scala 31:71]
  assign _GEN_633 = 10'h279 == WADDR ? 10'h279 : _GEN_632; // @[RAM_ST.scala 31:71]
  assign _GEN_634 = 10'h27a == WADDR ? 10'h27a : _GEN_633; // @[RAM_ST.scala 31:71]
  assign _GEN_635 = 10'h27b == WADDR ? 10'h27b : _GEN_634; // @[RAM_ST.scala 31:71]
  assign _GEN_636 = 10'h27c == WADDR ? 10'h27c : _GEN_635; // @[RAM_ST.scala 31:71]
  assign _GEN_637 = 10'h27d == WADDR ? 10'h27d : _GEN_636; // @[RAM_ST.scala 31:71]
  assign _GEN_638 = 10'h27e == WADDR ? 10'h27e : _GEN_637; // @[RAM_ST.scala 31:71]
  assign _GEN_639 = 10'h27f == WADDR ? 10'h27f : _GEN_638; // @[RAM_ST.scala 31:71]
  assign _GEN_640 = 10'h280 == WADDR ? 10'h280 : _GEN_639; // @[RAM_ST.scala 31:71]
  assign _GEN_641 = 10'h281 == WADDR ? 10'h281 : _GEN_640; // @[RAM_ST.scala 31:71]
  assign _GEN_642 = 10'h282 == WADDR ? 10'h282 : _GEN_641; // @[RAM_ST.scala 31:71]
  assign _GEN_643 = 10'h283 == WADDR ? 10'h283 : _GEN_642; // @[RAM_ST.scala 31:71]
  assign _GEN_644 = 10'h284 == WADDR ? 10'h284 : _GEN_643; // @[RAM_ST.scala 31:71]
  assign _GEN_645 = 10'h285 == WADDR ? 10'h285 : _GEN_644; // @[RAM_ST.scala 31:71]
  assign _GEN_646 = 10'h286 == WADDR ? 10'h286 : _GEN_645; // @[RAM_ST.scala 31:71]
  assign _GEN_647 = 10'h287 == WADDR ? 10'h287 : _GEN_646; // @[RAM_ST.scala 31:71]
  assign _GEN_648 = 10'h288 == WADDR ? 10'h288 : _GEN_647; // @[RAM_ST.scala 31:71]
  assign _GEN_649 = 10'h289 == WADDR ? 10'h289 : _GEN_648; // @[RAM_ST.scala 31:71]
  assign _GEN_650 = 10'h28a == WADDR ? 10'h28a : _GEN_649; // @[RAM_ST.scala 31:71]
  assign _GEN_651 = 10'h28b == WADDR ? 10'h28b : _GEN_650; // @[RAM_ST.scala 31:71]
  assign _GEN_652 = 10'h28c == WADDR ? 10'h28c : _GEN_651; // @[RAM_ST.scala 31:71]
  assign _GEN_653 = 10'h28d == WADDR ? 10'h28d : _GEN_652; // @[RAM_ST.scala 31:71]
  assign _GEN_654 = 10'h28e == WADDR ? 10'h28e : _GEN_653; // @[RAM_ST.scala 31:71]
  assign _GEN_655 = 10'h28f == WADDR ? 10'h28f : _GEN_654; // @[RAM_ST.scala 31:71]
  assign _GEN_656 = 10'h290 == WADDR ? 10'h290 : _GEN_655; // @[RAM_ST.scala 31:71]
  assign _GEN_657 = 10'h291 == WADDR ? 10'h291 : _GEN_656; // @[RAM_ST.scala 31:71]
  assign _GEN_658 = 10'h292 == WADDR ? 10'h292 : _GEN_657; // @[RAM_ST.scala 31:71]
  assign _GEN_659 = 10'h293 == WADDR ? 10'h293 : _GEN_658; // @[RAM_ST.scala 31:71]
  assign _GEN_660 = 10'h294 == WADDR ? 10'h294 : _GEN_659; // @[RAM_ST.scala 31:71]
  assign _GEN_661 = 10'h295 == WADDR ? 10'h295 : _GEN_660; // @[RAM_ST.scala 31:71]
  assign _GEN_662 = 10'h296 == WADDR ? 10'h296 : _GEN_661; // @[RAM_ST.scala 31:71]
  assign _GEN_663 = 10'h297 == WADDR ? 10'h297 : _GEN_662; // @[RAM_ST.scala 31:71]
  assign _GEN_664 = 10'h298 == WADDR ? 10'h298 : _GEN_663; // @[RAM_ST.scala 31:71]
  assign _GEN_665 = 10'h299 == WADDR ? 10'h299 : _GEN_664; // @[RAM_ST.scala 31:71]
  assign _GEN_666 = 10'h29a == WADDR ? 10'h29a : _GEN_665; // @[RAM_ST.scala 31:71]
  assign _GEN_667 = 10'h29b == WADDR ? 10'h29b : _GEN_666; // @[RAM_ST.scala 31:71]
  assign _GEN_668 = 10'h29c == WADDR ? 10'h29c : _GEN_667; // @[RAM_ST.scala 31:71]
  assign _GEN_669 = 10'h29d == WADDR ? 10'h29d : _GEN_668; // @[RAM_ST.scala 31:71]
  assign _GEN_670 = 10'h29e == WADDR ? 10'h29e : _GEN_669; // @[RAM_ST.scala 31:71]
  assign _GEN_671 = 10'h29f == WADDR ? 10'h29f : _GEN_670; // @[RAM_ST.scala 31:71]
  assign _GEN_672 = 10'h2a0 == WADDR ? 10'h2a0 : _GEN_671; // @[RAM_ST.scala 31:71]
  assign _GEN_673 = 10'h2a1 == WADDR ? 10'h2a1 : _GEN_672; // @[RAM_ST.scala 31:71]
  assign _GEN_674 = 10'h2a2 == WADDR ? 10'h2a2 : _GEN_673; // @[RAM_ST.scala 31:71]
  assign _GEN_675 = 10'h2a3 == WADDR ? 10'h2a3 : _GEN_674; // @[RAM_ST.scala 31:71]
  assign _GEN_676 = 10'h2a4 == WADDR ? 10'h2a4 : _GEN_675; // @[RAM_ST.scala 31:71]
  assign _GEN_677 = 10'h2a5 == WADDR ? 10'h2a5 : _GEN_676; // @[RAM_ST.scala 31:71]
  assign _GEN_678 = 10'h2a6 == WADDR ? 10'h2a6 : _GEN_677; // @[RAM_ST.scala 31:71]
  assign _GEN_679 = 10'h2a7 == WADDR ? 10'h2a7 : _GEN_678; // @[RAM_ST.scala 31:71]
  assign _GEN_680 = 10'h2a8 == WADDR ? 10'h2a8 : _GEN_679; // @[RAM_ST.scala 31:71]
  assign _GEN_681 = 10'h2a9 == WADDR ? 10'h2a9 : _GEN_680; // @[RAM_ST.scala 31:71]
  assign _GEN_682 = 10'h2aa == WADDR ? 10'h2aa : _GEN_681; // @[RAM_ST.scala 31:71]
  assign _GEN_683 = 10'h2ab == WADDR ? 10'h2ab : _GEN_682; // @[RAM_ST.scala 31:71]
  assign _GEN_684 = 10'h2ac == WADDR ? 10'h2ac : _GEN_683; // @[RAM_ST.scala 31:71]
  assign _GEN_685 = 10'h2ad == WADDR ? 10'h2ad : _GEN_684; // @[RAM_ST.scala 31:71]
  assign _GEN_686 = 10'h2ae == WADDR ? 10'h2ae : _GEN_685; // @[RAM_ST.scala 31:71]
  assign _GEN_687 = 10'h2af == WADDR ? 10'h2af : _GEN_686; // @[RAM_ST.scala 31:71]
  assign _GEN_688 = 10'h2b0 == WADDR ? 10'h2b0 : _GEN_687; // @[RAM_ST.scala 31:71]
  assign _GEN_689 = 10'h2b1 == WADDR ? 10'h2b1 : _GEN_688; // @[RAM_ST.scala 31:71]
  assign _GEN_690 = 10'h2b2 == WADDR ? 10'h2b2 : _GEN_689; // @[RAM_ST.scala 31:71]
  assign _GEN_691 = 10'h2b3 == WADDR ? 10'h2b3 : _GEN_690; // @[RAM_ST.scala 31:71]
  assign _GEN_692 = 10'h2b4 == WADDR ? 10'h2b4 : _GEN_691; // @[RAM_ST.scala 31:71]
  assign _GEN_693 = 10'h2b5 == WADDR ? 10'h2b5 : _GEN_692; // @[RAM_ST.scala 31:71]
  assign _GEN_694 = 10'h2b6 == WADDR ? 10'h2b6 : _GEN_693; // @[RAM_ST.scala 31:71]
  assign _GEN_695 = 10'h2b7 == WADDR ? 10'h2b7 : _GEN_694; // @[RAM_ST.scala 31:71]
  assign _GEN_696 = 10'h2b8 == WADDR ? 10'h2b8 : _GEN_695; // @[RAM_ST.scala 31:71]
  assign _GEN_697 = 10'h2b9 == WADDR ? 10'h2b9 : _GEN_696; // @[RAM_ST.scala 31:71]
  assign _GEN_698 = 10'h2ba == WADDR ? 10'h2ba : _GEN_697; // @[RAM_ST.scala 31:71]
  assign _GEN_699 = 10'h2bb == WADDR ? 10'h2bb : _GEN_698; // @[RAM_ST.scala 31:71]
  assign _GEN_700 = 10'h2bc == WADDR ? 10'h2bc : _GEN_699; // @[RAM_ST.scala 31:71]
  assign _GEN_701 = 10'h2bd == WADDR ? 10'h2bd : _GEN_700; // @[RAM_ST.scala 31:71]
  assign _GEN_702 = 10'h2be == WADDR ? 10'h2be : _GEN_701; // @[RAM_ST.scala 31:71]
  assign _GEN_703 = 10'h2bf == WADDR ? 10'h2bf : _GEN_702; // @[RAM_ST.scala 31:71]
  assign _GEN_704 = 10'h2c0 == WADDR ? 10'h2c0 : _GEN_703; // @[RAM_ST.scala 31:71]
  assign _GEN_705 = 10'h2c1 == WADDR ? 10'h2c1 : _GEN_704; // @[RAM_ST.scala 31:71]
  assign _GEN_706 = 10'h2c2 == WADDR ? 10'h2c2 : _GEN_705; // @[RAM_ST.scala 31:71]
  assign _GEN_707 = 10'h2c3 == WADDR ? 10'h2c3 : _GEN_706; // @[RAM_ST.scala 31:71]
  assign _GEN_708 = 10'h2c4 == WADDR ? 10'h2c4 : _GEN_707; // @[RAM_ST.scala 31:71]
  assign _GEN_709 = 10'h2c5 == WADDR ? 10'h2c5 : _GEN_708; // @[RAM_ST.scala 31:71]
  assign _GEN_710 = 10'h2c6 == WADDR ? 10'h2c6 : _GEN_709; // @[RAM_ST.scala 31:71]
  assign _GEN_711 = 10'h2c7 == WADDR ? 10'h2c7 : _GEN_710; // @[RAM_ST.scala 31:71]
  assign _GEN_712 = 10'h2c8 == WADDR ? 10'h2c8 : _GEN_711; // @[RAM_ST.scala 31:71]
  assign _GEN_713 = 10'h2c9 == WADDR ? 10'h2c9 : _GEN_712; // @[RAM_ST.scala 31:71]
  assign _GEN_714 = 10'h2ca == WADDR ? 10'h2ca : _GEN_713; // @[RAM_ST.scala 31:71]
  assign _GEN_715 = 10'h2cb == WADDR ? 10'h2cb : _GEN_714; // @[RAM_ST.scala 31:71]
  assign _GEN_716 = 10'h2cc == WADDR ? 10'h2cc : _GEN_715; // @[RAM_ST.scala 31:71]
  assign _GEN_717 = 10'h2cd == WADDR ? 10'h2cd : _GEN_716; // @[RAM_ST.scala 31:71]
  assign _GEN_718 = 10'h2ce == WADDR ? 10'h2ce : _GEN_717; // @[RAM_ST.scala 31:71]
  assign _GEN_719 = 10'h2cf == WADDR ? 10'h2cf : _GEN_718; // @[RAM_ST.scala 31:71]
  assign _GEN_720 = 10'h2d0 == WADDR ? 10'h2d0 : _GEN_719; // @[RAM_ST.scala 31:71]
  assign _GEN_721 = 10'h2d1 == WADDR ? 10'h2d1 : _GEN_720; // @[RAM_ST.scala 31:71]
  assign _GEN_722 = 10'h2d2 == WADDR ? 10'h2d2 : _GEN_721; // @[RAM_ST.scala 31:71]
  assign _GEN_723 = 10'h2d3 == WADDR ? 10'h2d3 : _GEN_722; // @[RAM_ST.scala 31:71]
  assign _GEN_724 = 10'h2d4 == WADDR ? 10'h2d4 : _GEN_723; // @[RAM_ST.scala 31:71]
  assign _GEN_725 = 10'h2d5 == WADDR ? 10'h2d5 : _GEN_724; // @[RAM_ST.scala 31:71]
  assign _GEN_726 = 10'h2d6 == WADDR ? 10'h2d6 : _GEN_725; // @[RAM_ST.scala 31:71]
  assign _GEN_727 = 10'h2d7 == WADDR ? 10'h2d7 : _GEN_726; // @[RAM_ST.scala 31:71]
  assign _GEN_728 = 10'h2d8 == WADDR ? 10'h2d8 : _GEN_727; // @[RAM_ST.scala 31:71]
  assign _GEN_729 = 10'h2d9 == WADDR ? 10'h2d9 : _GEN_728; // @[RAM_ST.scala 31:71]
  assign _GEN_730 = 10'h2da == WADDR ? 10'h2da : _GEN_729; // @[RAM_ST.scala 31:71]
  assign _GEN_731 = 10'h2db == WADDR ? 10'h2db : _GEN_730; // @[RAM_ST.scala 31:71]
  assign _GEN_732 = 10'h2dc == WADDR ? 10'h2dc : _GEN_731; // @[RAM_ST.scala 31:71]
  assign _GEN_733 = 10'h2dd == WADDR ? 10'h2dd : _GEN_732; // @[RAM_ST.scala 31:71]
  assign _GEN_734 = 10'h2de == WADDR ? 10'h2de : _GEN_733; // @[RAM_ST.scala 31:71]
  assign _GEN_735 = 10'h2df == WADDR ? 10'h2df : _GEN_734; // @[RAM_ST.scala 31:71]
  assign _GEN_736 = 10'h2e0 == WADDR ? 10'h2e0 : _GEN_735; // @[RAM_ST.scala 31:71]
  assign _GEN_737 = 10'h2e1 == WADDR ? 10'h2e1 : _GEN_736; // @[RAM_ST.scala 31:71]
  assign _GEN_738 = 10'h2e2 == WADDR ? 10'h2e2 : _GEN_737; // @[RAM_ST.scala 31:71]
  assign _GEN_739 = 10'h2e3 == WADDR ? 10'h2e3 : _GEN_738; // @[RAM_ST.scala 31:71]
  assign _GEN_740 = 10'h2e4 == WADDR ? 10'h2e4 : _GEN_739; // @[RAM_ST.scala 31:71]
  assign _GEN_741 = 10'h2e5 == WADDR ? 10'h2e5 : _GEN_740; // @[RAM_ST.scala 31:71]
  assign _GEN_742 = 10'h2e6 == WADDR ? 10'h2e6 : _GEN_741; // @[RAM_ST.scala 31:71]
  assign _GEN_743 = 10'h2e7 == WADDR ? 10'h2e7 : _GEN_742; // @[RAM_ST.scala 31:71]
  assign _GEN_744 = 10'h2e8 == WADDR ? 10'h2e8 : _GEN_743; // @[RAM_ST.scala 31:71]
  assign _GEN_745 = 10'h2e9 == WADDR ? 10'h2e9 : _GEN_744; // @[RAM_ST.scala 31:71]
  assign _GEN_746 = 10'h2ea == WADDR ? 10'h2ea : _GEN_745; // @[RAM_ST.scala 31:71]
  assign _GEN_747 = 10'h2eb == WADDR ? 10'h2eb : _GEN_746; // @[RAM_ST.scala 31:71]
  assign _GEN_748 = 10'h2ec == WADDR ? 10'h2ec : _GEN_747; // @[RAM_ST.scala 31:71]
  assign _GEN_749 = 10'h2ed == WADDR ? 10'h2ed : _GEN_748; // @[RAM_ST.scala 31:71]
  assign _GEN_750 = 10'h2ee == WADDR ? 10'h2ee : _GEN_749; // @[RAM_ST.scala 31:71]
  assign _GEN_751 = 10'h2ef == WADDR ? 10'h2ef : _GEN_750; // @[RAM_ST.scala 31:71]
  assign _GEN_752 = 10'h2f0 == WADDR ? 10'h2f0 : _GEN_751; // @[RAM_ST.scala 31:71]
  assign _GEN_753 = 10'h2f1 == WADDR ? 10'h2f1 : _GEN_752; // @[RAM_ST.scala 31:71]
  assign _GEN_754 = 10'h2f2 == WADDR ? 10'h2f2 : _GEN_753; // @[RAM_ST.scala 31:71]
  assign _GEN_755 = 10'h2f3 == WADDR ? 10'h2f3 : _GEN_754; // @[RAM_ST.scala 31:71]
  assign _GEN_756 = 10'h2f4 == WADDR ? 10'h2f4 : _GEN_755; // @[RAM_ST.scala 31:71]
  assign _GEN_757 = 10'h2f5 == WADDR ? 10'h2f5 : _GEN_756; // @[RAM_ST.scala 31:71]
  assign _GEN_758 = 10'h2f6 == WADDR ? 10'h2f6 : _GEN_757; // @[RAM_ST.scala 31:71]
  assign _GEN_759 = 10'h2f7 == WADDR ? 10'h2f7 : _GEN_758; // @[RAM_ST.scala 31:71]
  assign _GEN_760 = 10'h2f8 == WADDR ? 10'h2f8 : _GEN_759; // @[RAM_ST.scala 31:71]
  assign _GEN_761 = 10'h2f9 == WADDR ? 10'h2f9 : _GEN_760; // @[RAM_ST.scala 31:71]
  assign _GEN_762 = 10'h2fa == WADDR ? 10'h2fa : _GEN_761; // @[RAM_ST.scala 31:71]
  assign _GEN_763 = 10'h2fb == WADDR ? 10'h2fb : _GEN_762; // @[RAM_ST.scala 31:71]
  assign _GEN_764 = 10'h2fc == WADDR ? 10'h2fc : _GEN_763; // @[RAM_ST.scala 31:71]
  assign _GEN_765 = 10'h2fd == WADDR ? 10'h2fd : _GEN_764; // @[RAM_ST.scala 31:71]
  assign _GEN_766 = 10'h2fe == WADDR ? 10'h2fe : _GEN_765; // @[RAM_ST.scala 31:71]
  assign _GEN_767 = 10'h2ff == WADDR ? 10'h2ff : _GEN_766; // @[RAM_ST.scala 31:71]
  assign _GEN_768 = 10'h300 == WADDR ? 10'h300 : _GEN_767; // @[RAM_ST.scala 31:71]
  assign _GEN_769 = 10'h301 == WADDR ? 10'h301 : _GEN_768; // @[RAM_ST.scala 31:71]
  assign _GEN_770 = 10'h302 == WADDR ? 10'h302 : _GEN_769; // @[RAM_ST.scala 31:71]
  assign _GEN_771 = 10'h303 == WADDR ? 10'h303 : _GEN_770; // @[RAM_ST.scala 31:71]
  assign _GEN_772 = 10'h304 == WADDR ? 10'h304 : _GEN_771; // @[RAM_ST.scala 31:71]
  assign _GEN_773 = 10'h305 == WADDR ? 10'h305 : _GEN_772; // @[RAM_ST.scala 31:71]
  assign _GEN_774 = 10'h306 == WADDR ? 10'h306 : _GEN_773; // @[RAM_ST.scala 31:71]
  assign _GEN_775 = 10'h307 == WADDR ? 10'h307 : _GEN_774; // @[RAM_ST.scala 31:71]
  assign _GEN_776 = 10'h308 == WADDR ? 10'h308 : _GEN_775; // @[RAM_ST.scala 31:71]
  assign _GEN_777 = 10'h309 == WADDR ? 10'h309 : _GEN_776; // @[RAM_ST.scala 31:71]
  assign _GEN_778 = 10'h30a == WADDR ? 10'h30a : _GEN_777; // @[RAM_ST.scala 31:71]
  assign _GEN_779 = 10'h30b == WADDR ? 10'h30b : _GEN_778; // @[RAM_ST.scala 31:71]
  assign _GEN_780 = 10'h30c == WADDR ? 10'h30c : _GEN_779; // @[RAM_ST.scala 31:71]
  assign _GEN_781 = 10'h30d == WADDR ? 10'h30d : _GEN_780; // @[RAM_ST.scala 31:71]
  assign _GEN_782 = 10'h30e == WADDR ? 10'h30e : _GEN_781; // @[RAM_ST.scala 31:71]
  assign _GEN_783 = 10'h30f == WADDR ? 10'h30f : _GEN_782; // @[RAM_ST.scala 31:71]
  assign _GEN_784 = 10'h310 == WADDR ? 10'h310 : _GEN_783; // @[RAM_ST.scala 31:71]
  assign _GEN_785 = 10'h311 == WADDR ? 10'h311 : _GEN_784; // @[RAM_ST.scala 31:71]
  assign _GEN_786 = 10'h312 == WADDR ? 10'h312 : _GEN_785; // @[RAM_ST.scala 31:71]
  assign _GEN_787 = 10'h313 == WADDR ? 10'h313 : _GEN_786; // @[RAM_ST.scala 31:71]
  assign _GEN_788 = 10'h314 == WADDR ? 10'h314 : _GEN_787; // @[RAM_ST.scala 31:71]
  assign _GEN_789 = 10'h315 == WADDR ? 10'h315 : _GEN_788; // @[RAM_ST.scala 31:71]
  assign _GEN_790 = 10'h316 == WADDR ? 10'h316 : _GEN_789; // @[RAM_ST.scala 31:71]
  assign _GEN_791 = 10'h317 == WADDR ? 10'h317 : _GEN_790; // @[RAM_ST.scala 31:71]
  assign _GEN_792 = 10'h318 == WADDR ? 10'h318 : _GEN_791; // @[RAM_ST.scala 31:71]
  assign _GEN_793 = 10'h319 == WADDR ? 10'h319 : _GEN_792; // @[RAM_ST.scala 31:71]
  assign _GEN_794 = 10'h31a == WADDR ? 10'h31a : _GEN_793; // @[RAM_ST.scala 31:71]
  assign _GEN_795 = 10'h31b == WADDR ? 10'h31b : _GEN_794; // @[RAM_ST.scala 31:71]
  assign _GEN_796 = 10'h31c == WADDR ? 10'h31c : _GEN_795; // @[RAM_ST.scala 31:71]
  assign _GEN_797 = 10'h31d == WADDR ? 10'h31d : _GEN_796; // @[RAM_ST.scala 31:71]
  assign _GEN_798 = 10'h31e == WADDR ? 10'h31e : _GEN_797; // @[RAM_ST.scala 31:71]
  assign _GEN_799 = 10'h31f == WADDR ? 10'h31f : _GEN_798; // @[RAM_ST.scala 31:71]
  assign _GEN_800 = 10'h320 == WADDR ? 10'h320 : _GEN_799; // @[RAM_ST.scala 31:71]
  assign _GEN_801 = 10'h321 == WADDR ? 10'h321 : _GEN_800; // @[RAM_ST.scala 31:71]
  assign _GEN_802 = 10'h322 == WADDR ? 10'h322 : _GEN_801; // @[RAM_ST.scala 31:71]
  assign _GEN_803 = 10'h323 == WADDR ? 10'h323 : _GEN_802; // @[RAM_ST.scala 31:71]
  assign _GEN_804 = 10'h324 == WADDR ? 10'h324 : _GEN_803; // @[RAM_ST.scala 31:71]
  assign _GEN_805 = 10'h325 == WADDR ? 10'h325 : _GEN_804; // @[RAM_ST.scala 31:71]
  assign _GEN_806 = 10'h326 == WADDR ? 10'h326 : _GEN_805; // @[RAM_ST.scala 31:71]
  assign _GEN_807 = 10'h327 == WADDR ? 10'h327 : _GEN_806; // @[RAM_ST.scala 31:71]
  assign _GEN_808 = 10'h328 == WADDR ? 10'h328 : _GEN_807; // @[RAM_ST.scala 31:71]
  assign _GEN_809 = 10'h329 == WADDR ? 10'h329 : _GEN_808; // @[RAM_ST.scala 31:71]
  assign _GEN_810 = 10'h32a == WADDR ? 10'h32a : _GEN_809; // @[RAM_ST.scala 31:71]
  assign _GEN_811 = 10'h32b == WADDR ? 10'h32b : _GEN_810; // @[RAM_ST.scala 31:71]
  assign _GEN_812 = 10'h32c == WADDR ? 10'h32c : _GEN_811; // @[RAM_ST.scala 31:71]
  assign _GEN_813 = 10'h32d == WADDR ? 10'h32d : _GEN_812; // @[RAM_ST.scala 31:71]
  assign _GEN_814 = 10'h32e == WADDR ? 10'h32e : _GEN_813; // @[RAM_ST.scala 31:71]
  assign _GEN_815 = 10'h32f == WADDR ? 10'h32f : _GEN_814; // @[RAM_ST.scala 31:71]
  assign _GEN_816 = 10'h330 == WADDR ? 10'h330 : _GEN_815; // @[RAM_ST.scala 31:71]
  assign _GEN_817 = 10'h331 == WADDR ? 10'h331 : _GEN_816; // @[RAM_ST.scala 31:71]
  assign _GEN_818 = 10'h332 == WADDR ? 10'h332 : _GEN_817; // @[RAM_ST.scala 31:71]
  assign _GEN_819 = 10'h333 == WADDR ? 10'h333 : _GEN_818; // @[RAM_ST.scala 31:71]
  assign _GEN_820 = 10'h334 == WADDR ? 10'h334 : _GEN_819; // @[RAM_ST.scala 31:71]
  assign _GEN_821 = 10'h335 == WADDR ? 10'h335 : _GEN_820; // @[RAM_ST.scala 31:71]
  assign _GEN_822 = 10'h336 == WADDR ? 10'h336 : _GEN_821; // @[RAM_ST.scala 31:71]
  assign _GEN_823 = 10'h337 == WADDR ? 10'h337 : _GEN_822; // @[RAM_ST.scala 31:71]
  assign _GEN_824 = 10'h338 == WADDR ? 10'h338 : _GEN_823; // @[RAM_ST.scala 31:71]
  assign _GEN_825 = 10'h339 == WADDR ? 10'h339 : _GEN_824; // @[RAM_ST.scala 31:71]
  assign _GEN_826 = 10'h33a == WADDR ? 10'h33a : _GEN_825; // @[RAM_ST.scala 31:71]
  assign _GEN_827 = 10'h33b == WADDR ? 10'h33b : _GEN_826; // @[RAM_ST.scala 31:71]
  assign _GEN_828 = 10'h33c == WADDR ? 10'h33c : _GEN_827; // @[RAM_ST.scala 31:71]
  assign _GEN_829 = 10'h33d == WADDR ? 10'h33d : _GEN_828; // @[RAM_ST.scala 31:71]
  assign _GEN_830 = 10'h33e == WADDR ? 10'h33e : _GEN_829; // @[RAM_ST.scala 31:71]
  assign _GEN_831 = 10'h33f == WADDR ? 10'h33f : _GEN_830; // @[RAM_ST.scala 31:71]
  assign _GEN_832 = 10'h340 == WADDR ? 10'h340 : _GEN_831; // @[RAM_ST.scala 31:71]
  assign _GEN_833 = 10'h341 == WADDR ? 10'h341 : _GEN_832; // @[RAM_ST.scala 31:71]
  assign _GEN_834 = 10'h342 == WADDR ? 10'h342 : _GEN_833; // @[RAM_ST.scala 31:71]
  assign _GEN_835 = 10'h343 == WADDR ? 10'h343 : _GEN_834; // @[RAM_ST.scala 31:71]
  assign _GEN_836 = 10'h344 == WADDR ? 10'h344 : _GEN_835; // @[RAM_ST.scala 31:71]
  assign _GEN_837 = 10'h345 == WADDR ? 10'h345 : _GEN_836; // @[RAM_ST.scala 31:71]
  assign _GEN_838 = 10'h346 == WADDR ? 10'h346 : _GEN_837; // @[RAM_ST.scala 31:71]
  assign _GEN_839 = 10'h347 == WADDR ? 10'h347 : _GEN_838; // @[RAM_ST.scala 31:71]
  assign _GEN_840 = 10'h348 == WADDR ? 10'h348 : _GEN_839; // @[RAM_ST.scala 31:71]
  assign _GEN_841 = 10'h349 == WADDR ? 10'h349 : _GEN_840; // @[RAM_ST.scala 31:71]
  assign _GEN_842 = 10'h34a == WADDR ? 10'h34a : _GEN_841; // @[RAM_ST.scala 31:71]
  assign _GEN_843 = 10'h34b == WADDR ? 10'h34b : _GEN_842; // @[RAM_ST.scala 31:71]
  assign _GEN_844 = 10'h34c == WADDR ? 10'h34c : _GEN_843; // @[RAM_ST.scala 31:71]
  assign _GEN_845 = 10'h34d == WADDR ? 10'h34d : _GEN_844; // @[RAM_ST.scala 31:71]
  assign _GEN_846 = 10'h34e == WADDR ? 10'h34e : _GEN_845; // @[RAM_ST.scala 31:71]
  assign _GEN_847 = 10'h34f == WADDR ? 10'h34f : _GEN_846; // @[RAM_ST.scala 31:71]
  assign _GEN_848 = 10'h350 == WADDR ? 10'h350 : _GEN_847; // @[RAM_ST.scala 31:71]
  assign _GEN_849 = 10'h351 == WADDR ? 10'h351 : _GEN_848; // @[RAM_ST.scala 31:71]
  assign _GEN_850 = 10'h352 == WADDR ? 10'h352 : _GEN_849; // @[RAM_ST.scala 31:71]
  assign _GEN_851 = 10'h353 == WADDR ? 10'h353 : _GEN_850; // @[RAM_ST.scala 31:71]
  assign _GEN_852 = 10'h354 == WADDR ? 10'h354 : _GEN_851; // @[RAM_ST.scala 31:71]
  assign _GEN_853 = 10'h355 == WADDR ? 10'h355 : _GEN_852; // @[RAM_ST.scala 31:71]
  assign _GEN_854 = 10'h356 == WADDR ? 10'h356 : _GEN_853; // @[RAM_ST.scala 31:71]
  assign _GEN_855 = 10'h357 == WADDR ? 10'h357 : _GEN_854; // @[RAM_ST.scala 31:71]
  assign _GEN_856 = 10'h358 == WADDR ? 10'h358 : _GEN_855; // @[RAM_ST.scala 31:71]
  assign _GEN_857 = 10'h359 == WADDR ? 10'h359 : _GEN_856; // @[RAM_ST.scala 31:71]
  assign _GEN_858 = 10'h35a == WADDR ? 10'h35a : _GEN_857; // @[RAM_ST.scala 31:71]
  assign _GEN_859 = 10'h35b == WADDR ? 10'h35b : _GEN_858; // @[RAM_ST.scala 31:71]
  assign _GEN_860 = 10'h35c == WADDR ? 10'h35c : _GEN_859; // @[RAM_ST.scala 31:71]
  assign _GEN_861 = 10'h35d == WADDR ? 10'h35d : _GEN_860; // @[RAM_ST.scala 31:71]
  assign _GEN_862 = 10'h35e == WADDR ? 10'h35e : _GEN_861; // @[RAM_ST.scala 31:71]
  assign _GEN_863 = 10'h35f == WADDR ? 10'h35f : _GEN_862; // @[RAM_ST.scala 31:71]
  assign _GEN_864 = 10'h360 == WADDR ? 10'h360 : _GEN_863; // @[RAM_ST.scala 31:71]
  assign _GEN_865 = 10'h361 == WADDR ? 10'h361 : _GEN_864; // @[RAM_ST.scala 31:71]
  assign _GEN_866 = 10'h362 == WADDR ? 10'h362 : _GEN_865; // @[RAM_ST.scala 31:71]
  assign _GEN_867 = 10'h363 == WADDR ? 10'h363 : _GEN_866; // @[RAM_ST.scala 31:71]
  assign _GEN_868 = 10'h364 == WADDR ? 10'h364 : _GEN_867; // @[RAM_ST.scala 31:71]
  assign _GEN_869 = 10'h365 == WADDR ? 10'h365 : _GEN_868; // @[RAM_ST.scala 31:71]
  assign _GEN_870 = 10'h366 == WADDR ? 10'h366 : _GEN_869; // @[RAM_ST.scala 31:71]
  assign _GEN_871 = 10'h367 == WADDR ? 10'h367 : _GEN_870; // @[RAM_ST.scala 31:71]
  assign _GEN_872 = 10'h368 == WADDR ? 10'h368 : _GEN_871; // @[RAM_ST.scala 31:71]
  assign _GEN_873 = 10'h369 == WADDR ? 10'h369 : _GEN_872; // @[RAM_ST.scala 31:71]
  assign _GEN_874 = 10'h36a == WADDR ? 10'h36a : _GEN_873; // @[RAM_ST.scala 31:71]
  assign _GEN_875 = 10'h36b == WADDR ? 10'h36b : _GEN_874; // @[RAM_ST.scala 31:71]
  assign _GEN_876 = 10'h36c == WADDR ? 10'h36c : _GEN_875; // @[RAM_ST.scala 31:71]
  assign _GEN_877 = 10'h36d == WADDR ? 10'h36d : _GEN_876; // @[RAM_ST.scala 31:71]
  assign _GEN_878 = 10'h36e == WADDR ? 10'h36e : _GEN_877; // @[RAM_ST.scala 31:71]
  assign _GEN_879 = 10'h36f == WADDR ? 10'h36f : _GEN_878; // @[RAM_ST.scala 31:71]
  assign _GEN_880 = 10'h370 == WADDR ? 10'h370 : _GEN_879; // @[RAM_ST.scala 31:71]
  assign _GEN_881 = 10'h371 == WADDR ? 10'h371 : _GEN_880; // @[RAM_ST.scala 31:71]
  assign _GEN_882 = 10'h372 == WADDR ? 10'h372 : _GEN_881; // @[RAM_ST.scala 31:71]
  assign _GEN_883 = 10'h373 == WADDR ? 10'h373 : _GEN_882; // @[RAM_ST.scala 31:71]
  assign _GEN_884 = 10'h374 == WADDR ? 10'h374 : _GEN_883; // @[RAM_ST.scala 31:71]
  assign _GEN_885 = 10'h375 == WADDR ? 10'h375 : _GEN_884; // @[RAM_ST.scala 31:71]
  assign _GEN_886 = 10'h376 == WADDR ? 10'h376 : _GEN_885; // @[RAM_ST.scala 31:71]
  assign _GEN_887 = 10'h377 == WADDR ? 10'h377 : _GEN_886; // @[RAM_ST.scala 31:71]
  assign _GEN_888 = 10'h378 == WADDR ? 10'h378 : _GEN_887; // @[RAM_ST.scala 31:71]
  assign _GEN_889 = 10'h379 == WADDR ? 10'h379 : _GEN_888; // @[RAM_ST.scala 31:71]
  assign _GEN_890 = 10'h37a == WADDR ? 10'h37a : _GEN_889; // @[RAM_ST.scala 31:71]
  assign _GEN_891 = 10'h37b == WADDR ? 10'h37b : _GEN_890; // @[RAM_ST.scala 31:71]
  assign _GEN_892 = 10'h37c == WADDR ? 10'h37c : _GEN_891; // @[RAM_ST.scala 31:71]
  assign _GEN_893 = 10'h37d == WADDR ? 10'h37d : _GEN_892; // @[RAM_ST.scala 31:71]
  assign _GEN_894 = 10'h37e == WADDR ? 10'h37e : _GEN_893; // @[RAM_ST.scala 31:71]
  assign _GEN_895 = 10'h37f == WADDR ? 10'h37f : _GEN_894; // @[RAM_ST.scala 31:71]
  assign _GEN_896 = 10'h380 == WADDR ? 10'h380 : _GEN_895; // @[RAM_ST.scala 31:71]
  assign _GEN_897 = 10'h381 == WADDR ? 10'h381 : _GEN_896; // @[RAM_ST.scala 31:71]
  assign _GEN_898 = 10'h382 == WADDR ? 10'h382 : _GEN_897; // @[RAM_ST.scala 31:71]
  assign _GEN_899 = 10'h383 == WADDR ? 10'h383 : _GEN_898; // @[RAM_ST.scala 31:71]
  assign _GEN_900 = 10'h384 == WADDR ? 10'h384 : _GEN_899; // @[RAM_ST.scala 31:71]
  assign _GEN_901 = 10'h385 == WADDR ? 10'h385 : _GEN_900; // @[RAM_ST.scala 31:71]
  assign _GEN_902 = 10'h386 == WADDR ? 10'h386 : _GEN_901; // @[RAM_ST.scala 31:71]
  assign _GEN_903 = 10'h387 == WADDR ? 10'h387 : _GEN_902; // @[RAM_ST.scala 31:71]
  assign _GEN_904 = 10'h388 == WADDR ? 10'h388 : _GEN_903; // @[RAM_ST.scala 31:71]
  assign _GEN_905 = 10'h389 == WADDR ? 10'h389 : _GEN_904; // @[RAM_ST.scala 31:71]
  assign _GEN_906 = 10'h38a == WADDR ? 10'h38a : _GEN_905; // @[RAM_ST.scala 31:71]
  assign _GEN_907 = 10'h38b == WADDR ? 10'h38b : _GEN_906; // @[RAM_ST.scala 31:71]
  assign _GEN_908 = 10'h38c == WADDR ? 10'h38c : _GEN_907; // @[RAM_ST.scala 31:71]
  assign _GEN_909 = 10'h38d == WADDR ? 10'h38d : _GEN_908; // @[RAM_ST.scala 31:71]
  assign _GEN_910 = 10'h38e == WADDR ? 10'h38e : _GEN_909; // @[RAM_ST.scala 31:71]
  assign _GEN_911 = 10'h38f == WADDR ? 10'h38f : _GEN_910; // @[RAM_ST.scala 31:71]
  assign _GEN_912 = 10'h390 == WADDR ? 10'h390 : _GEN_911; // @[RAM_ST.scala 31:71]
  assign _GEN_913 = 10'h391 == WADDR ? 10'h391 : _GEN_912; // @[RAM_ST.scala 31:71]
  assign _GEN_914 = 10'h392 == WADDR ? 10'h392 : _GEN_913; // @[RAM_ST.scala 31:71]
  assign _GEN_915 = 10'h393 == WADDR ? 10'h393 : _GEN_914; // @[RAM_ST.scala 31:71]
  assign _GEN_916 = 10'h394 == WADDR ? 10'h394 : _GEN_915; // @[RAM_ST.scala 31:71]
  assign _GEN_917 = 10'h395 == WADDR ? 10'h395 : _GEN_916; // @[RAM_ST.scala 31:71]
  assign _GEN_918 = 10'h396 == WADDR ? 10'h396 : _GEN_917; // @[RAM_ST.scala 31:71]
  assign _GEN_919 = 10'h397 == WADDR ? 10'h397 : _GEN_918; // @[RAM_ST.scala 31:71]
  assign _GEN_920 = 10'h398 == WADDR ? 10'h398 : _GEN_919; // @[RAM_ST.scala 31:71]
  assign _GEN_921 = 10'h399 == WADDR ? 10'h399 : _GEN_920; // @[RAM_ST.scala 31:71]
  assign _GEN_922 = 10'h39a == WADDR ? 10'h39a : _GEN_921; // @[RAM_ST.scala 31:71]
  assign _GEN_923 = 10'h39b == WADDR ? 10'h39b : _GEN_922; // @[RAM_ST.scala 31:71]
  assign _GEN_924 = 10'h39c == WADDR ? 10'h39c : _GEN_923; // @[RAM_ST.scala 31:71]
  assign _GEN_925 = 10'h39d == WADDR ? 10'h39d : _GEN_924; // @[RAM_ST.scala 31:71]
  assign _GEN_926 = 10'h39e == WADDR ? 10'h39e : _GEN_925; // @[RAM_ST.scala 31:71]
  assign _GEN_927 = 10'h39f == WADDR ? 10'h39f : _GEN_926; // @[RAM_ST.scala 31:71]
  assign _GEN_928 = 10'h3a0 == WADDR ? 10'h3a0 : _GEN_927; // @[RAM_ST.scala 31:71]
  assign _GEN_929 = 10'h3a1 == WADDR ? 10'h3a1 : _GEN_928; // @[RAM_ST.scala 31:71]
  assign _GEN_930 = 10'h3a2 == WADDR ? 10'h3a2 : _GEN_929; // @[RAM_ST.scala 31:71]
  assign _GEN_931 = 10'h3a3 == WADDR ? 10'h3a3 : _GEN_930; // @[RAM_ST.scala 31:71]
  assign _GEN_932 = 10'h3a4 == WADDR ? 10'h3a4 : _GEN_931; // @[RAM_ST.scala 31:71]
  assign _GEN_933 = 10'h3a5 == WADDR ? 10'h3a5 : _GEN_932; // @[RAM_ST.scala 31:71]
  assign _GEN_934 = 10'h3a6 == WADDR ? 10'h3a6 : _GEN_933; // @[RAM_ST.scala 31:71]
  assign _GEN_935 = 10'h3a7 == WADDR ? 10'h3a7 : _GEN_934; // @[RAM_ST.scala 31:71]
  assign _GEN_936 = 10'h3a8 == WADDR ? 10'h3a8 : _GEN_935; // @[RAM_ST.scala 31:71]
  assign _GEN_937 = 10'h3a9 == WADDR ? 10'h3a9 : _GEN_936; // @[RAM_ST.scala 31:71]
  assign _GEN_938 = 10'h3aa == WADDR ? 10'h3aa : _GEN_937; // @[RAM_ST.scala 31:71]
  assign _GEN_939 = 10'h3ab == WADDR ? 10'h3ab : _GEN_938; // @[RAM_ST.scala 31:71]
  assign _GEN_940 = 10'h3ac == WADDR ? 10'h3ac : _GEN_939; // @[RAM_ST.scala 31:71]
  assign _GEN_941 = 10'h3ad == WADDR ? 10'h3ad : _GEN_940; // @[RAM_ST.scala 31:71]
  assign _GEN_942 = 10'h3ae == WADDR ? 10'h3ae : _GEN_941; // @[RAM_ST.scala 31:71]
  assign _GEN_943 = 10'h3af == WADDR ? 10'h3af : _GEN_942; // @[RAM_ST.scala 31:71]
  assign _GEN_944 = 10'h3b0 == WADDR ? 10'h3b0 : _GEN_943; // @[RAM_ST.scala 31:71]
  assign _GEN_945 = 10'h3b1 == WADDR ? 10'h3b1 : _GEN_944; // @[RAM_ST.scala 31:71]
  assign _GEN_946 = 10'h3b2 == WADDR ? 10'h3b2 : _GEN_945; // @[RAM_ST.scala 31:71]
  assign _GEN_947 = 10'h3b3 == WADDR ? 10'h3b3 : _GEN_946; // @[RAM_ST.scala 31:71]
  assign _GEN_948 = 10'h3b4 == WADDR ? 10'h3b4 : _GEN_947; // @[RAM_ST.scala 31:71]
  assign _GEN_949 = 10'h3b5 == WADDR ? 10'h3b5 : _GEN_948; // @[RAM_ST.scala 31:71]
  assign _GEN_950 = 10'h3b6 == WADDR ? 10'h3b6 : _GEN_949; // @[RAM_ST.scala 31:71]
  assign _GEN_951 = 10'h3b7 == WADDR ? 10'h3b7 : _GEN_950; // @[RAM_ST.scala 31:71]
  assign _GEN_952 = 10'h3b8 == WADDR ? 10'h3b8 : _GEN_951; // @[RAM_ST.scala 31:71]
  assign _GEN_953 = 10'h3b9 == WADDR ? 10'h3b9 : _GEN_952; // @[RAM_ST.scala 31:71]
  assign _GEN_954 = 10'h3ba == WADDR ? 10'h3ba : _GEN_953; // @[RAM_ST.scala 31:71]
  assign _GEN_955 = 10'h3bb == WADDR ? 10'h3bb : _GEN_954; // @[RAM_ST.scala 31:71]
  assign _GEN_956 = 10'h3bc == WADDR ? 10'h3bc : _GEN_955; // @[RAM_ST.scala 31:71]
  assign _GEN_957 = 10'h3bd == WADDR ? 10'h3bd : _GEN_956; // @[RAM_ST.scala 31:71]
  assign _GEN_958 = 10'h3be == WADDR ? 10'h3be : _GEN_957; // @[RAM_ST.scala 31:71]
  assign _GEN_959 = 10'h3bf == WADDR ? 10'h3bf : _GEN_958; // @[RAM_ST.scala 31:71]
  assign _T = {{1'd0}, _GEN_959}; // @[RAM_ST.scala 31:71]
  assign _GEN_966 = 10'h1 == RADDR ? 10'h1 : 10'h0; // @[RAM_ST.scala 32:46]
  assign _GEN_967 = 10'h2 == RADDR ? 10'h2 : _GEN_966; // @[RAM_ST.scala 32:46]
  assign _GEN_968 = 10'h3 == RADDR ? 10'h3 : _GEN_967; // @[RAM_ST.scala 32:46]
  assign _GEN_969 = 10'h4 == RADDR ? 10'h4 : _GEN_968; // @[RAM_ST.scala 32:46]
  assign _GEN_970 = 10'h5 == RADDR ? 10'h5 : _GEN_969; // @[RAM_ST.scala 32:46]
  assign _GEN_971 = 10'h6 == RADDR ? 10'h6 : _GEN_970; // @[RAM_ST.scala 32:46]
  assign _GEN_972 = 10'h7 == RADDR ? 10'h7 : _GEN_971; // @[RAM_ST.scala 32:46]
  assign _GEN_973 = 10'h8 == RADDR ? 10'h8 : _GEN_972; // @[RAM_ST.scala 32:46]
  assign _GEN_974 = 10'h9 == RADDR ? 10'h9 : _GEN_973; // @[RAM_ST.scala 32:46]
  assign _GEN_975 = 10'ha == RADDR ? 10'ha : _GEN_974; // @[RAM_ST.scala 32:46]
  assign _GEN_976 = 10'hb == RADDR ? 10'hb : _GEN_975; // @[RAM_ST.scala 32:46]
  assign _GEN_977 = 10'hc == RADDR ? 10'hc : _GEN_976; // @[RAM_ST.scala 32:46]
  assign _GEN_978 = 10'hd == RADDR ? 10'hd : _GEN_977; // @[RAM_ST.scala 32:46]
  assign _GEN_979 = 10'he == RADDR ? 10'he : _GEN_978; // @[RAM_ST.scala 32:46]
  assign _GEN_980 = 10'hf == RADDR ? 10'hf : _GEN_979; // @[RAM_ST.scala 32:46]
  assign _GEN_981 = 10'h10 == RADDR ? 10'h10 : _GEN_980; // @[RAM_ST.scala 32:46]
  assign _GEN_982 = 10'h11 == RADDR ? 10'h11 : _GEN_981; // @[RAM_ST.scala 32:46]
  assign _GEN_983 = 10'h12 == RADDR ? 10'h12 : _GEN_982; // @[RAM_ST.scala 32:46]
  assign _GEN_984 = 10'h13 == RADDR ? 10'h13 : _GEN_983; // @[RAM_ST.scala 32:46]
  assign _GEN_985 = 10'h14 == RADDR ? 10'h14 : _GEN_984; // @[RAM_ST.scala 32:46]
  assign _GEN_986 = 10'h15 == RADDR ? 10'h15 : _GEN_985; // @[RAM_ST.scala 32:46]
  assign _GEN_987 = 10'h16 == RADDR ? 10'h16 : _GEN_986; // @[RAM_ST.scala 32:46]
  assign _GEN_988 = 10'h17 == RADDR ? 10'h17 : _GEN_987; // @[RAM_ST.scala 32:46]
  assign _GEN_989 = 10'h18 == RADDR ? 10'h18 : _GEN_988; // @[RAM_ST.scala 32:46]
  assign _GEN_990 = 10'h19 == RADDR ? 10'h19 : _GEN_989; // @[RAM_ST.scala 32:46]
  assign _GEN_991 = 10'h1a == RADDR ? 10'h1a : _GEN_990; // @[RAM_ST.scala 32:46]
  assign _GEN_992 = 10'h1b == RADDR ? 10'h1b : _GEN_991; // @[RAM_ST.scala 32:46]
  assign _GEN_993 = 10'h1c == RADDR ? 10'h1c : _GEN_992; // @[RAM_ST.scala 32:46]
  assign _GEN_994 = 10'h1d == RADDR ? 10'h1d : _GEN_993; // @[RAM_ST.scala 32:46]
  assign _GEN_995 = 10'h1e == RADDR ? 10'h1e : _GEN_994; // @[RAM_ST.scala 32:46]
  assign _GEN_996 = 10'h1f == RADDR ? 10'h1f : _GEN_995; // @[RAM_ST.scala 32:46]
  assign _GEN_997 = 10'h20 == RADDR ? 10'h20 : _GEN_996; // @[RAM_ST.scala 32:46]
  assign _GEN_998 = 10'h21 == RADDR ? 10'h21 : _GEN_997; // @[RAM_ST.scala 32:46]
  assign _GEN_999 = 10'h22 == RADDR ? 10'h22 : _GEN_998; // @[RAM_ST.scala 32:46]
  assign _GEN_1000 = 10'h23 == RADDR ? 10'h23 : _GEN_999; // @[RAM_ST.scala 32:46]
  assign _GEN_1001 = 10'h24 == RADDR ? 10'h24 : _GEN_1000; // @[RAM_ST.scala 32:46]
  assign _GEN_1002 = 10'h25 == RADDR ? 10'h25 : _GEN_1001; // @[RAM_ST.scala 32:46]
  assign _GEN_1003 = 10'h26 == RADDR ? 10'h26 : _GEN_1002; // @[RAM_ST.scala 32:46]
  assign _GEN_1004 = 10'h27 == RADDR ? 10'h27 : _GEN_1003; // @[RAM_ST.scala 32:46]
  assign _GEN_1005 = 10'h28 == RADDR ? 10'h28 : _GEN_1004; // @[RAM_ST.scala 32:46]
  assign _GEN_1006 = 10'h29 == RADDR ? 10'h29 : _GEN_1005; // @[RAM_ST.scala 32:46]
  assign _GEN_1007 = 10'h2a == RADDR ? 10'h2a : _GEN_1006; // @[RAM_ST.scala 32:46]
  assign _GEN_1008 = 10'h2b == RADDR ? 10'h2b : _GEN_1007; // @[RAM_ST.scala 32:46]
  assign _GEN_1009 = 10'h2c == RADDR ? 10'h2c : _GEN_1008; // @[RAM_ST.scala 32:46]
  assign _GEN_1010 = 10'h2d == RADDR ? 10'h2d : _GEN_1009; // @[RAM_ST.scala 32:46]
  assign _GEN_1011 = 10'h2e == RADDR ? 10'h2e : _GEN_1010; // @[RAM_ST.scala 32:46]
  assign _GEN_1012 = 10'h2f == RADDR ? 10'h2f : _GEN_1011; // @[RAM_ST.scala 32:46]
  assign _GEN_1013 = 10'h30 == RADDR ? 10'h30 : _GEN_1012; // @[RAM_ST.scala 32:46]
  assign _GEN_1014 = 10'h31 == RADDR ? 10'h31 : _GEN_1013; // @[RAM_ST.scala 32:46]
  assign _GEN_1015 = 10'h32 == RADDR ? 10'h32 : _GEN_1014; // @[RAM_ST.scala 32:46]
  assign _GEN_1016 = 10'h33 == RADDR ? 10'h33 : _GEN_1015; // @[RAM_ST.scala 32:46]
  assign _GEN_1017 = 10'h34 == RADDR ? 10'h34 : _GEN_1016; // @[RAM_ST.scala 32:46]
  assign _GEN_1018 = 10'h35 == RADDR ? 10'h35 : _GEN_1017; // @[RAM_ST.scala 32:46]
  assign _GEN_1019 = 10'h36 == RADDR ? 10'h36 : _GEN_1018; // @[RAM_ST.scala 32:46]
  assign _GEN_1020 = 10'h37 == RADDR ? 10'h37 : _GEN_1019; // @[RAM_ST.scala 32:46]
  assign _GEN_1021 = 10'h38 == RADDR ? 10'h38 : _GEN_1020; // @[RAM_ST.scala 32:46]
  assign _GEN_1022 = 10'h39 == RADDR ? 10'h39 : _GEN_1021; // @[RAM_ST.scala 32:46]
  assign _GEN_1023 = 10'h3a == RADDR ? 10'h3a : _GEN_1022; // @[RAM_ST.scala 32:46]
  assign _GEN_1024 = 10'h3b == RADDR ? 10'h3b : _GEN_1023; // @[RAM_ST.scala 32:46]
  assign _GEN_1025 = 10'h3c == RADDR ? 10'h3c : _GEN_1024; // @[RAM_ST.scala 32:46]
  assign _GEN_1026 = 10'h3d == RADDR ? 10'h3d : _GEN_1025; // @[RAM_ST.scala 32:46]
  assign _GEN_1027 = 10'h3e == RADDR ? 10'h3e : _GEN_1026; // @[RAM_ST.scala 32:46]
  assign _GEN_1028 = 10'h3f == RADDR ? 10'h3f : _GEN_1027; // @[RAM_ST.scala 32:46]
  assign _GEN_1029 = 10'h40 == RADDR ? 10'h40 : _GEN_1028; // @[RAM_ST.scala 32:46]
  assign _GEN_1030 = 10'h41 == RADDR ? 10'h41 : _GEN_1029; // @[RAM_ST.scala 32:46]
  assign _GEN_1031 = 10'h42 == RADDR ? 10'h42 : _GEN_1030; // @[RAM_ST.scala 32:46]
  assign _GEN_1032 = 10'h43 == RADDR ? 10'h43 : _GEN_1031; // @[RAM_ST.scala 32:46]
  assign _GEN_1033 = 10'h44 == RADDR ? 10'h44 : _GEN_1032; // @[RAM_ST.scala 32:46]
  assign _GEN_1034 = 10'h45 == RADDR ? 10'h45 : _GEN_1033; // @[RAM_ST.scala 32:46]
  assign _GEN_1035 = 10'h46 == RADDR ? 10'h46 : _GEN_1034; // @[RAM_ST.scala 32:46]
  assign _GEN_1036 = 10'h47 == RADDR ? 10'h47 : _GEN_1035; // @[RAM_ST.scala 32:46]
  assign _GEN_1037 = 10'h48 == RADDR ? 10'h48 : _GEN_1036; // @[RAM_ST.scala 32:46]
  assign _GEN_1038 = 10'h49 == RADDR ? 10'h49 : _GEN_1037; // @[RAM_ST.scala 32:46]
  assign _GEN_1039 = 10'h4a == RADDR ? 10'h4a : _GEN_1038; // @[RAM_ST.scala 32:46]
  assign _GEN_1040 = 10'h4b == RADDR ? 10'h4b : _GEN_1039; // @[RAM_ST.scala 32:46]
  assign _GEN_1041 = 10'h4c == RADDR ? 10'h4c : _GEN_1040; // @[RAM_ST.scala 32:46]
  assign _GEN_1042 = 10'h4d == RADDR ? 10'h4d : _GEN_1041; // @[RAM_ST.scala 32:46]
  assign _GEN_1043 = 10'h4e == RADDR ? 10'h4e : _GEN_1042; // @[RAM_ST.scala 32:46]
  assign _GEN_1044 = 10'h4f == RADDR ? 10'h4f : _GEN_1043; // @[RAM_ST.scala 32:46]
  assign _GEN_1045 = 10'h50 == RADDR ? 10'h50 : _GEN_1044; // @[RAM_ST.scala 32:46]
  assign _GEN_1046 = 10'h51 == RADDR ? 10'h51 : _GEN_1045; // @[RAM_ST.scala 32:46]
  assign _GEN_1047 = 10'h52 == RADDR ? 10'h52 : _GEN_1046; // @[RAM_ST.scala 32:46]
  assign _GEN_1048 = 10'h53 == RADDR ? 10'h53 : _GEN_1047; // @[RAM_ST.scala 32:46]
  assign _GEN_1049 = 10'h54 == RADDR ? 10'h54 : _GEN_1048; // @[RAM_ST.scala 32:46]
  assign _GEN_1050 = 10'h55 == RADDR ? 10'h55 : _GEN_1049; // @[RAM_ST.scala 32:46]
  assign _GEN_1051 = 10'h56 == RADDR ? 10'h56 : _GEN_1050; // @[RAM_ST.scala 32:46]
  assign _GEN_1052 = 10'h57 == RADDR ? 10'h57 : _GEN_1051; // @[RAM_ST.scala 32:46]
  assign _GEN_1053 = 10'h58 == RADDR ? 10'h58 : _GEN_1052; // @[RAM_ST.scala 32:46]
  assign _GEN_1054 = 10'h59 == RADDR ? 10'h59 : _GEN_1053; // @[RAM_ST.scala 32:46]
  assign _GEN_1055 = 10'h5a == RADDR ? 10'h5a : _GEN_1054; // @[RAM_ST.scala 32:46]
  assign _GEN_1056 = 10'h5b == RADDR ? 10'h5b : _GEN_1055; // @[RAM_ST.scala 32:46]
  assign _GEN_1057 = 10'h5c == RADDR ? 10'h5c : _GEN_1056; // @[RAM_ST.scala 32:46]
  assign _GEN_1058 = 10'h5d == RADDR ? 10'h5d : _GEN_1057; // @[RAM_ST.scala 32:46]
  assign _GEN_1059 = 10'h5e == RADDR ? 10'h5e : _GEN_1058; // @[RAM_ST.scala 32:46]
  assign _GEN_1060 = 10'h5f == RADDR ? 10'h5f : _GEN_1059; // @[RAM_ST.scala 32:46]
  assign _GEN_1061 = 10'h60 == RADDR ? 10'h60 : _GEN_1060; // @[RAM_ST.scala 32:46]
  assign _GEN_1062 = 10'h61 == RADDR ? 10'h61 : _GEN_1061; // @[RAM_ST.scala 32:46]
  assign _GEN_1063 = 10'h62 == RADDR ? 10'h62 : _GEN_1062; // @[RAM_ST.scala 32:46]
  assign _GEN_1064 = 10'h63 == RADDR ? 10'h63 : _GEN_1063; // @[RAM_ST.scala 32:46]
  assign _GEN_1065 = 10'h64 == RADDR ? 10'h64 : _GEN_1064; // @[RAM_ST.scala 32:46]
  assign _GEN_1066 = 10'h65 == RADDR ? 10'h65 : _GEN_1065; // @[RAM_ST.scala 32:46]
  assign _GEN_1067 = 10'h66 == RADDR ? 10'h66 : _GEN_1066; // @[RAM_ST.scala 32:46]
  assign _GEN_1068 = 10'h67 == RADDR ? 10'h67 : _GEN_1067; // @[RAM_ST.scala 32:46]
  assign _GEN_1069 = 10'h68 == RADDR ? 10'h68 : _GEN_1068; // @[RAM_ST.scala 32:46]
  assign _GEN_1070 = 10'h69 == RADDR ? 10'h69 : _GEN_1069; // @[RAM_ST.scala 32:46]
  assign _GEN_1071 = 10'h6a == RADDR ? 10'h6a : _GEN_1070; // @[RAM_ST.scala 32:46]
  assign _GEN_1072 = 10'h6b == RADDR ? 10'h6b : _GEN_1071; // @[RAM_ST.scala 32:46]
  assign _GEN_1073 = 10'h6c == RADDR ? 10'h6c : _GEN_1072; // @[RAM_ST.scala 32:46]
  assign _GEN_1074 = 10'h6d == RADDR ? 10'h6d : _GEN_1073; // @[RAM_ST.scala 32:46]
  assign _GEN_1075 = 10'h6e == RADDR ? 10'h6e : _GEN_1074; // @[RAM_ST.scala 32:46]
  assign _GEN_1076 = 10'h6f == RADDR ? 10'h6f : _GEN_1075; // @[RAM_ST.scala 32:46]
  assign _GEN_1077 = 10'h70 == RADDR ? 10'h70 : _GEN_1076; // @[RAM_ST.scala 32:46]
  assign _GEN_1078 = 10'h71 == RADDR ? 10'h71 : _GEN_1077; // @[RAM_ST.scala 32:46]
  assign _GEN_1079 = 10'h72 == RADDR ? 10'h72 : _GEN_1078; // @[RAM_ST.scala 32:46]
  assign _GEN_1080 = 10'h73 == RADDR ? 10'h73 : _GEN_1079; // @[RAM_ST.scala 32:46]
  assign _GEN_1081 = 10'h74 == RADDR ? 10'h74 : _GEN_1080; // @[RAM_ST.scala 32:46]
  assign _GEN_1082 = 10'h75 == RADDR ? 10'h75 : _GEN_1081; // @[RAM_ST.scala 32:46]
  assign _GEN_1083 = 10'h76 == RADDR ? 10'h76 : _GEN_1082; // @[RAM_ST.scala 32:46]
  assign _GEN_1084 = 10'h77 == RADDR ? 10'h77 : _GEN_1083; // @[RAM_ST.scala 32:46]
  assign _GEN_1085 = 10'h78 == RADDR ? 10'h78 : _GEN_1084; // @[RAM_ST.scala 32:46]
  assign _GEN_1086 = 10'h79 == RADDR ? 10'h79 : _GEN_1085; // @[RAM_ST.scala 32:46]
  assign _GEN_1087 = 10'h7a == RADDR ? 10'h7a : _GEN_1086; // @[RAM_ST.scala 32:46]
  assign _GEN_1088 = 10'h7b == RADDR ? 10'h7b : _GEN_1087; // @[RAM_ST.scala 32:46]
  assign _GEN_1089 = 10'h7c == RADDR ? 10'h7c : _GEN_1088; // @[RAM_ST.scala 32:46]
  assign _GEN_1090 = 10'h7d == RADDR ? 10'h7d : _GEN_1089; // @[RAM_ST.scala 32:46]
  assign _GEN_1091 = 10'h7e == RADDR ? 10'h7e : _GEN_1090; // @[RAM_ST.scala 32:46]
  assign _GEN_1092 = 10'h7f == RADDR ? 10'h7f : _GEN_1091; // @[RAM_ST.scala 32:46]
  assign _GEN_1093 = 10'h80 == RADDR ? 10'h80 : _GEN_1092; // @[RAM_ST.scala 32:46]
  assign _GEN_1094 = 10'h81 == RADDR ? 10'h81 : _GEN_1093; // @[RAM_ST.scala 32:46]
  assign _GEN_1095 = 10'h82 == RADDR ? 10'h82 : _GEN_1094; // @[RAM_ST.scala 32:46]
  assign _GEN_1096 = 10'h83 == RADDR ? 10'h83 : _GEN_1095; // @[RAM_ST.scala 32:46]
  assign _GEN_1097 = 10'h84 == RADDR ? 10'h84 : _GEN_1096; // @[RAM_ST.scala 32:46]
  assign _GEN_1098 = 10'h85 == RADDR ? 10'h85 : _GEN_1097; // @[RAM_ST.scala 32:46]
  assign _GEN_1099 = 10'h86 == RADDR ? 10'h86 : _GEN_1098; // @[RAM_ST.scala 32:46]
  assign _GEN_1100 = 10'h87 == RADDR ? 10'h87 : _GEN_1099; // @[RAM_ST.scala 32:46]
  assign _GEN_1101 = 10'h88 == RADDR ? 10'h88 : _GEN_1100; // @[RAM_ST.scala 32:46]
  assign _GEN_1102 = 10'h89 == RADDR ? 10'h89 : _GEN_1101; // @[RAM_ST.scala 32:46]
  assign _GEN_1103 = 10'h8a == RADDR ? 10'h8a : _GEN_1102; // @[RAM_ST.scala 32:46]
  assign _GEN_1104 = 10'h8b == RADDR ? 10'h8b : _GEN_1103; // @[RAM_ST.scala 32:46]
  assign _GEN_1105 = 10'h8c == RADDR ? 10'h8c : _GEN_1104; // @[RAM_ST.scala 32:46]
  assign _GEN_1106 = 10'h8d == RADDR ? 10'h8d : _GEN_1105; // @[RAM_ST.scala 32:46]
  assign _GEN_1107 = 10'h8e == RADDR ? 10'h8e : _GEN_1106; // @[RAM_ST.scala 32:46]
  assign _GEN_1108 = 10'h8f == RADDR ? 10'h8f : _GEN_1107; // @[RAM_ST.scala 32:46]
  assign _GEN_1109 = 10'h90 == RADDR ? 10'h90 : _GEN_1108; // @[RAM_ST.scala 32:46]
  assign _GEN_1110 = 10'h91 == RADDR ? 10'h91 : _GEN_1109; // @[RAM_ST.scala 32:46]
  assign _GEN_1111 = 10'h92 == RADDR ? 10'h92 : _GEN_1110; // @[RAM_ST.scala 32:46]
  assign _GEN_1112 = 10'h93 == RADDR ? 10'h93 : _GEN_1111; // @[RAM_ST.scala 32:46]
  assign _GEN_1113 = 10'h94 == RADDR ? 10'h94 : _GEN_1112; // @[RAM_ST.scala 32:46]
  assign _GEN_1114 = 10'h95 == RADDR ? 10'h95 : _GEN_1113; // @[RAM_ST.scala 32:46]
  assign _GEN_1115 = 10'h96 == RADDR ? 10'h96 : _GEN_1114; // @[RAM_ST.scala 32:46]
  assign _GEN_1116 = 10'h97 == RADDR ? 10'h97 : _GEN_1115; // @[RAM_ST.scala 32:46]
  assign _GEN_1117 = 10'h98 == RADDR ? 10'h98 : _GEN_1116; // @[RAM_ST.scala 32:46]
  assign _GEN_1118 = 10'h99 == RADDR ? 10'h99 : _GEN_1117; // @[RAM_ST.scala 32:46]
  assign _GEN_1119 = 10'h9a == RADDR ? 10'h9a : _GEN_1118; // @[RAM_ST.scala 32:46]
  assign _GEN_1120 = 10'h9b == RADDR ? 10'h9b : _GEN_1119; // @[RAM_ST.scala 32:46]
  assign _GEN_1121 = 10'h9c == RADDR ? 10'h9c : _GEN_1120; // @[RAM_ST.scala 32:46]
  assign _GEN_1122 = 10'h9d == RADDR ? 10'h9d : _GEN_1121; // @[RAM_ST.scala 32:46]
  assign _GEN_1123 = 10'h9e == RADDR ? 10'h9e : _GEN_1122; // @[RAM_ST.scala 32:46]
  assign _GEN_1124 = 10'h9f == RADDR ? 10'h9f : _GEN_1123; // @[RAM_ST.scala 32:46]
  assign _GEN_1125 = 10'ha0 == RADDR ? 10'ha0 : _GEN_1124; // @[RAM_ST.scala 32:46]
  assign _GEN_1126 = 10'ha1 == RADDR ? 10'ha1 : _GEN_1125; // @[RAM_ST.scala 32:46]
  assign _GEN_1127 = 10'ha2 == RADDR ? 10'ha2 : _GEN_1126; // @[RAM_ST.scala 32:46]
  assign _GEN_1128 = 10'ha3 == RADDR ? 10'ha3 : _GEN_1127; // @[RAM_ST.scala 32:46]
  assign _GEN_1129 = 10'ha4 == RADDR ? 10'ha4 : _GEN_1128; // @[RAM_ST.scala 32:46]
  assign _GEN_1130 = 10'ha5 == RADDR ? 10'ha5 : _GEN_1129; // @[RAM_ST.scala 32:46]
  assign _GEN_1131 = 10'ha6 == RADDR ? 10'ha6 : _GEN_1130; // @[RAM_ST.scala 32:46]
  assign _GEN_1132 = 10'ha7 == RADDR ? 10'ha7 : _GEN_1131; // @[RAM_ST.scala 32:46]
  assign _GEN_1133 = 10'ha8 == RADDR ? 10'ha8 : _GEN_1132; // @[RAM_ST.scala 32:46]
  assign _GEN_1134 = 10'ha9 == RADDR ? 10'ha9 : _GEN_1133; // @[RAM_ST.scala 32:46]
  assign _GEN_1135 = 10'haa == RADDR ? 10'haa : _GEN_1134; // @[RAM_ST.scala 32:46]
  assign _GEN_1136 = 10'hab == RADDR ? 10'hab : _GEN_1135; // @[RAM_ST.scala 32:46]
  assign _GEN_1137 = 10'hac == RADDR ? 10'hac : _GEN_1136; // @[RAM_ST.scala 32:46]
  assign _GEN_1138 = 10'had == RADDR ? 10'had : _GEN_1137; // @[RAM_ST.scala 32:46]
  assign _GEN_1139 = 10'hae == RADDR ? 10'hae : _GEN_1138; // @[RAM_ST.scala 32:46]
  assign _GEN_1140 = 10'haf == RADDR ? 10'haf : _GEN_1139; // @[RAM_ST.scala 32:46]
  assign _GEN_1141 = 10'hb0 == RADDR ? 10'hb0 : _GEN_1140; // @[RAM_ST.scala 32:46]
  assign _GEN_1142 = 10'hb1 == RADDR ? 10'hb1 : _GEN_1141; // @[RAM_ST.scala 32:46]
  assign _GEN_1143 = 10'hb2 == RADDR ? 10'hb2 : _GEN_1142; // @[RAM_ST.scala 32:46]
  assign _GEN_1144 = 10'hb3 == RADDR ? 10'hb3 : _GEN_1143; // @[RAM_ST.scala 32:46]
  assign _GEN_1145 = 10'hb4 == RADDR ? 10'hb4 : _GEN_1144; // @[RAM_ST.scala 32:46]
  assign _GEN_1146 = 10'hb5 == RADDR ? 10'hb5 : _GEN_1145; // @[RAM_ST.scala 32:46]
  assign _GEN_1147 = 10'hb6 == RADDR ? 10'hb6 : _GEN_1146; // @[RAM_ST.scala 32:46]
  assign _GEN_1148 = 10'hb7 == RADDR ? 10'hb7 : _GEN_1147; // @[RAM_ST.scala 32:46]
  assign _GEN_1149 = 10'hb8 == RADDR ? 10'hb8 : _GEN_1148; // @[RAM_ST.scala 32:46]
  assign _GEN_1150 = 10'hb9 == RADDR ? 10'hb9 : _GEN_1149; // @[RAM_ST.scala 32:46]
  assign _GEN_1151 = 10'hba == RADDR ? 10'hba : _GEN_1150; // @[RAM_ST.scala 32:46]
  assign _GEN_1152 = 10'hbb == RADDR ? 10'hbb : _GEN_1151; // @[RAM_ST.scala 32:46]
  assign _GEN_1153 = 10'hbc == RADDR ? 10'hbc : _GEN_1152; // @[RAM_ST.scala 32:46]
  assign _GEN_1154 = 10'hbd == RADDR ? 10'hbd : _GEN_1153; // @[RAM_ST.scala 32:46]
  assign _GEN_1155 = 10'hbe == RADDR ? 10'hbe : _GEN_1154; // @[RAM_ST.scala 32:46]
  assign _GEN_1156 = 10'hbf == RADDR ? 10'hbf : _GEN_1155; // @[RAM_ST.scala 32:46]
  assign _GEN_1157 = 10'hc0 == RADDR ? 10'hc0 : _GEN_1156; // @[RAM_ST.scala 32:46]
  assign _GEN_1158 = 10'hc1 == RADDR ? 10'hc1 : _GEN_1157; // @[RAM_ST.scala 32:46]
  assign _GEN_1159 = 10'hc2 == RADDR ? 10'hc2 : _GEN_1158; // @[RAM_ST.scala 32:46]
  assign _GEN_1160 = 10'hc3 == RADDR ? 10'hc3 : _GEN_1159; // @[RAM_ST.scala 32:46]
  assign _GEN_1161 = 10'hc4 == RADDR ? 10'hc4 : _GEN_1160; // @[RAM_ST.scala 32:46]
  assign _GEN_1162 = 10'hc5 == RADDR ? 10'hc5 : _GEN_1161; // @[RAM_ST.scala 32:46]
  assign _GEN_1163 = 10'hc6 == RADDR ? 10'hc6 : _GEN_1162; // @[RAM_ST.scala 32:46]
  assign _GEN_1164 = 10'hc7 == RADDR ? 10'hc7 : _GEN_1163; // @[RAM_ST.scala 32:46]
  assign _GEN_1165 = 10'hc8 == RADDR ? 10'hc8 : _GEN_1164; // @[RAM_ST.scala 32:46]
  assign _GEN_1166 = 10'hc9 == RADDR ? 10'hc9 : _GEN_1165; // @[RAM_ST.scala 32:46]
  assign _GEN_1167 = 10'hca == RADDR ? 10'hca : _GEN_1166; // @[RAM_ST.scala 32:46]
  assign _GEN_1168 = 10'hcb == RADDR ? 10'hcb : _GEN_1167; // @[RAM_ST.scala 32:46]
  assign _GEN_1169 = 10'hcc == RADDR ? 10'hcc : _GEN_1168; // @[RAM_ST.scala 32:46]
  assign _GEN_1170 = 10'hcd == RADDR ? 10'hcd : _GEN_1169; // @[RAM_ST.scala 32:46]
  assign _GEN_1171 = 10'hce == RADDR ? 10'hce : _GEN_1170; // @[RAM_ST.scala 32:46]
  assign _GEN_1172 = 10'hcf == RADDR ? 10'hcf : _GEN_1171; // @[RAM_ST.scala 32:46]
  assign _GEN_1173 = 10'hd0 == RADDR ? 10'hd0 : _GEN_1172; // @[RAM_ST.scala 32:46]
  assign _GEN_1174 = 10'hd1 == RADDR ? 10'hd1 : _GEN_1173; // @[RAM_ST.scala 32:46]
  assign _GEN_1175 = 10'hd2 == RADDR ? 10'hd2 : _GEN_1174; // @[RAM_ST.scala 32:46]
  assign _GEN_1176 = 10'hd3 == RADDR ? 10'hd3 : _GEN_1175; // @[RAM_ST.scala 32:46]
  assign _GEN_1177 = 10'hd4 == RADDR ? 10'hd4 : _GEN_1176; // @[RAM_ST.scala 32:46]
  assign _GEN_1178 = 10'hd5 == RADDR ? 10'hd5 : _GEN_1177; // @[RAM_ST.scala 32:46]
  assign _GEN_1179 = 10'hd6 == RADDR ? 10'hd6 : _GEN_1178; // @[RAM_ST.scala 32:46]
  assign _GEN_1180 = 10'hd7 == RADDR ? 10'hd7 : _GEN_1179; // @[RAM_ST.scala 32:46]
  assign _GEN_1181 = 10'hd8 == RADDR ? 10'hd8 : _GEN_1180; // @[RAM_ST.scala 32:46]
  assign _GEN_1182 = 10'hd9 == RADDR ? 10'hd9 : _GEN_1181; // @[RAM_ST.scala 32:46]
  assign _GEN_1183 = 10'hda == RADDR ? 10'hda : _GEN_1182; // @[RAM_ST.scala 32:46]
  assign _GEN_1184 = 10'hdb == RADDR ? 10'hdb : _GEN_1183; // @[RAM_ST.scala 32:46]
  assign _GEN_1185 = 10'hdc == RADDR ? 10'hdc : _GEN_1184; // @[RAM_ST.scala 32:46]
  assign _GEN_1186 = 10'hdd == RADDR ? 10'hdd : _GEN_1185; // @[RAM_ST.scala 32:46]
  assign _GEN_1187 = 10'hde == RADDR ? 10'hde : _GEN_1186; // @[RAM_ST.scala 32:46]
  assign _GEN_1188 = 10'hdf == RADDR ? 10'hdf : _GEN_1187; // @[RAM_ST.scala 32:46]
  assign _GEN_1189 = 10'he0 == RADDR ? 10'he0 : _GEN_1188; // @[RAM_ST.scala 32:46]
  assign _GEN_1190 = 10'he1 == RADDR ? 10'he1 : _GEN_1189; // @[RAM_ST.scala 32:46]
  assign _GEN_1191 = 10'he2 == RADDR ? 10'he2 : _GEN_1190; // @[RAM_ST.scala 32:46]
  assign _GEN_1192 = 10'he3 == RADDR ? 10'he3 : _GEN_1191; // @[RAM_ST.scala 32:46]
  assign _GEN_1193 = 10'he4 == RADDR ? 10'he4 : _GEN_1192; // @[RAM_ST.scala 32:46]
  assign _GEN_1194 = 10'he5 == RADDR ? 10'he5 : _GEN_1193; // @[RAM_ST.scala 32:46]
  assign _GEN_1195 = 10'he6 == RADDR ? 10'he6 : _GEN_1194; // @[RAM_ST.scala 32:46]
  assign _GEN_1196 = 10'he7 == RADDR ? 10'he7 : _GEN_1195; // @[RAM_ST.scala 32:46]
  assign _GEN_1197 = 10'he8 == RADDR ? 10'he8 : _GEN_1196; // @[RAM_ST.scala 32:46]
  assign _GEN_1198 = 10'he9 == RADDR ? 10'he9 : _GEN_1197; // @[RAM_ST.scala 32:46]
  assign _GEN_1199 = 10'hea == RADDR ? 10'hea : _GEN_1198; // @[RAM_ST.scala 32:46]
  assign _GEN_1200 = 10'heb == RADDR ? 10'heb : _GEN_1199; // @[RAM_ST.scala 32:46]
  assign _GEN_1201 = 10'hec == RADDR ? 10'hec : _GEN_1200; // @[RAM_ST.scala 32:46]
  assign _GEN_1202 = 10'hed == RADDR ? 10'hed : _GEN_1201; // @[RAM_ST.scala 32:46]
  assign _GEN_1203 = 10'hee == RADDR ? 10'hee : _GEN_1202; // @[RAM_ST.scala 32:46]
  assign _GEN_1204 = 10'hef == RADDR ? 10'hef : _GEN_1203; // @[RAM_ST.scala 32:46]
  assign _GEN_1205 = 10'hf0 == RADDR ? 10'hf0 : _GEN_1204; // @[RAM_ST.scala 32:46]
  assign _GEN_1206 = 10'hf1 == RADDR ? 10'hf1 : _GEN_1205; // @[RAM_ST.scala 32:46]
  assign _GEN_1207 = 10'hf2 == RADDR ? 10'hf2 : _GEN_1206; // @[RAM_ST.scala 32:46]
  assign _GEN_1208 = 10'hf3 == RADDR ? 10'hf3 : _GEN_1207; // @[RAM_ST.scala 32:46]
  assign _GEN_1209 = 10'hf4 == RADDR ? 10'hf4 : _GEN_1208; // @[RAM_ST.scala 32:46]
  assign _GEN_1210 = 10'hf5 == RADDR ? 10'hf5 : _GEN_1209; // @[RAM_ST.scala 32:46]
  assign _GEN_1211 = 10'hf6 == RADDR ? 10'hf6 : _GEN_1210; // @[RAM_ST.scala 32:46]
  assign _GEN_1212 = 10'hf7 == RADDR ? 10'hf7 : _GEN_1211; // @[RAM_ST.scala 32:46]
  assign _GEN_1213 = 10'hf8 == RADDR ? 10'hf8 : _GEN_1212; // @[RAM_ST.scala 32:46]
  assign _GEN_1214 = 10'hf9 == RADDR ? 10'hf9 : _GEN_1213; // @[RAM_ST.scala 32:46]
  assign _GEN_1215 = 10'hfa == RADDR ? 10'hfa : _GEN_1214; // @[RAM_ST.scala 32:46]
  assign _GEN_1216 = 10'hfb == RADDR ? 10'hfb : _GEN_1215; // @[RAM_ST.scala 32:46]
  assign _GEN_1217 = 10'hfc == RADDR ? 10'hfc : _GEN_1216; // @[RAM_ST.scala 32:46]
  assign _GEN_1218 = 10'hfd == RADDR ? 10'hfd : _GEN_1217; // @[RAM_ST.scala 32:46]
  assign _GEN_1219 = 10'hfe == RADDR ? 10'hfe : _GEN_1218; // @[RAM_ST.scala 32:46]
  assign _GEN_1220 = 10'hff == RADDR ? 10'hff : _GEN_1219; // @[RAM_ST.scala 32:46]
  assign _GEN_1221 = 10'h100 == RADDR ? 10'h100 : _GEN_1220; // @[RAM_ST.scala 32:46]
  assign _GEN_1222 = 10'h101 == RADDR ? 10'h101 : _GEN_1221; // @[RAM_ST.scala 32:46]
  assign _GEN_1223 = 10'h102 == RADDR ? 10'h102 : _GEN_1222; // @[RAM_ST.scala 32:46]
  assign _GEN_1224 = 10'h103 == RADDR ? 10'h103 : _GEN_1223; // @[RAM_ST.scala 32:46]
  assign _GEN_1225 = 10'h104 == RADDR ? 10'h104 : _GEN_1224; // @[RAM_ST.scala 32:46]
  assign _GEN_1226 = 10'h105 == RADDR ? 10'h105 : _GEN_1225; // @[RAM_ST.scala 32:46]
  assign _GEN_1227 = 10'h106 == RADDR ? 10'h106 : _GEN_1226; // @[RAM_ST.scala 32:46]
  assign _GEN_1228 = 10'h107 == RADDR ? 10'h107 : _GEN_1227; // @[RAM_ST.scala 32:46]
  assign _GEN_1229 = 10'h108 == RADDR ? 10'h108 : _GEN_1228; // @[RAM_ST.scala 32:46]
  assign _GEN_1230 = 10'h109 == RADDR ? 10'h109 : _GEN_1229; // @[RAM_ST.scala 32:46]
  assign _GEN_1231 = 10'h10a == RADDR ? 10'h10a : _GEN_1230; // @[RAM_ST.scala 32:46]
  assign _GEN_1232 = 10'h10b == RADDR ? 10'h10b : _GEN_1231; // @[RAM_ST.scala 32:46]
  assign _GEN_1233 = 10'h10c == RADDR ? 10'h10c : _GEN_1232; // @[RAM_ST.scala 32:46]
  assign _GEN_1234 = 10'h10d == RADDR ? 10'h10d : _GEN_1233; // @[RAM_ST.scala 32:46]
  assign _GEN_1235 = 10'h10e == RADDR ? 10'h10e : _GEN_1234; // @[RAM_ST.scala 32:46]
  assign _GEN_1236 = 10'h10f == RADDR ? 10'h10f : _GEN_1235; // @[RAM_ST.scala 32:46]
  assign _GEN_1237 = 10'h110 == RADDR ? 10'h110 : _GEN_1236; // @[RAM_ST.scala 32:46]
  assign _GEN_1238 = 10'h111 == RADDR ? 10'h111 : _GEN_1237; // @[RAM_ST.scala 32:46]
  assign _GEN_1239 = 10'h112 == RADDR ? 10'h112 : _GEN_1238; // @[RAM_ST.scala 32:46]
  assign _GEN_1240 = 10'h113 == RADDR ? 10'h113 : _GEN_1239; // @[RAM_ST.scala 32:46]
  assign _GEN_1241 = 10'h114 == RADDR ? 10'h114 : _GEN_1240; // @[RAM_ST.scala 32:46]
  assign _GEN_1242 = 10'h115 == RADDR ? 10'h115 : _GEN_1241; // @[RAM_ST.scala 32:46]
  assign _GEN_1243 = 10'h116 == RADDR ? 10'h116 : _GEN_1242; // @[RAM_ST.scala 32:46]
  assign _GEN_1244 = 10'h117 == RADDR ? 10'h117 : _GEN_1243; // @[RAM_ST.scala 32:46]
  assign _GEN_1245 = 10'h118 == RADDR ? 10'h118 : _GEN_1244; // @[RAM_ST.scala 32:46]
  assign _GEN_1246 = 10'h119 == RADDR ? 10'h119 : _GEN_1245; // @[RAM_ST.scala 32:46]
  assign _GEN_1247 = 10'h11a == RADDR ? 10'h11a : _GEN_1246; // @[RAM_ST.scala 32:46]
  assign _GEN_1248 = 10'h11b == RADDR ? 10'h11b : _GEN_1247; // @[RAM_ST.scala 32:46]
  assign _GEN_1249 = 10'h11c == RADDR ? 10'h11c : _GEN_1248; // @[RAM_ST.scala 32:46]
  assign _GEN_1250 = 10'h11d == RADDR ? 10'h11d : _GEN_1249; // @[RAM_ST.scala 32:46]
  assign _GEN_1251 = 10'h11e == RADDR ? 10'h11e : _GEN_1250; // @[RAM_ST.scala 32:46]
  assign _GEN_1252 = 10'h11f == RADDR ? 10'h11f : _GEN_1251; // @[RAM_ST.scala 32:46]
  assign _GEN_1253 = 10'h120 == RADDR ? 10'h120 : _GEN_1252; // @[RAM_ST.scala 32:46]
  assign _GEN_1254 = 10'h121 == RADDR ? 10'h121 : _GEN_1253; // @[RAM_ST.scala 32:46]
  assign _GEN_1255 = 10'h122 == RADDR ? 10'h122 : _GEN_1254; // @[RAM_ST.scala 32:46]
  assign _GEN_1256 = 10'h123 == RADDR ? 10'h123 : _GEN_1255; // @[RAM_ST.scala 32:46]
  assign _GEN_1257 = 10'h124 == RADDR ? 10'h124 : _GEN_1256; // @[RAM_ST.scala 32:46]
  assign _GEN_1258 = 10'h125 == RADDR ? 10'h125 : _GEN_1257; // @[RAM_ST.scala 32:46]
  assign _GEN_1259 = 10'h126 == RADDR ? 10'h126 : _GEN_1258; // @[RAM_ST.scala 32:46]
  assign _GEN_1260 = 10'h127 == RADDR ? 10'h127 : _GEN_1259; // @[RAM_ST.scala 32:46]
  assign _GEN_1261 = 10'h128 == RADDR ? 10'h128 : _GEN_1260; // @[RAM_ST.scala 32:46]
  assign _GEN_1262 = 10'h129 == RADDR ? 10'h129 : _GEN_1261; // @[RAM_ST.scala 32:46]
  assign _GEN_1263 = 10'h12a == RADDR ? 10'h12a : _GEN_1262; // @[RAM_ST.scala 32:46]
  assign _GEN_1264 = 10'h12b == RADDR ? 10'h12b : _GEN_1263; // @[RAM_ST.scala 32:46]
  assign _GEN_1265 = 10'h12c == RADDR ? 10'h12c : _GEN_1264; // @[RAM_ST.scala 32:46]
  assign _GEN_1266 = 10'h12d == RADDR ? 10'h12d : _GEN_1265; // @[RAM_ST.scala 32:46]
  assign _GEN_1267 = 10'h12e == RADDR ? 10'h12e : _GEN_1266; // @[RAM_ST.scala 32:46]
  assign _GEN_1268 = 10'h12f == RADDR ? 10'h12f : _GEN_1267; // @[RAM_ST.scala 32:46]
  assign _GEN_1269 = 10'h130 == RADDR ? 10'h130 : _GEN_1268; // @[RAM_ST.scala 32:46]
  assign _GEN_1270 = 10'h131 == RADDR ? 10'h131 : _GEN_1269; // @[RAM_ST.scala 32:46]
  assign _GEN_1271 = 10'h132 == RADDR ? 10'h132 : _GEN_1270; // @[RAM_ST.scala 32:46]
  assign _GEN_1272 = 10'h133 == RADDR ? 10'h133 : _GEN_1271; // @[RAM_ST.scala 32:46]
  assign _GEN_1273 = 10'h134 == RADDR ? 10'h134 : _GEN_1272; // @[RAM_ST.scala 32:46]
  assign _GEN_1274 = 10'h135 == RADDR ? 10'h135 : _GEN_1273; // @[RAM_ST.scala 32:46]
  assign _GEN_1275 = 10'h136 == RADDR ? 10'h136 : _GEN_1274; // @[RAM_ST.scala 32:46]
  assign _GEN_1276 = 10'h137 == RADDR ? 10'h137 : _GEN_1275; // @[RAM_ST.scala 32:46]
  assign _GEN_1277 = 10'h138 == RADDR ? 10'h138 : _GEN_1276; // @[RAM_ST.scala 32:46]
  assign _GEN_1278 = 10'h139 == RADDR ? 10'h139 : _GEN_1277; // @[RAM_ST.scala 32:46]
  assign _GEN_1279 = 10'h13a == RADDR ? 10'h13a : _GEN_1278; // @[RAM_ST.scala 32:46]
  assign _GEN_1280 = 10'h13b == RADDR ? 10'h13b : _GEN_1279; // @[RAM_ST.scala 32:46]
  assign _GEN_1281 = 10'h13c == RADDR ? 10'h13c : _GEN_1280; // @[RAM_ST.scala 32:46]
  assign _GEN_1282 = 10'h13d == RADDR ? 10'h13d : _GEN_1281; // @[RAM_ST.scala 32:46]
  assign _GEN_1283 = 10'h13e == RADDR ? 10'h13e : _GEN_1282; // @[RAM_ST.scala 32:46]
  assign _GEN_1284 = 10'h13f == RADDR ? 10'h13f : _GEN_1283; // @[RAM_ST.scala 32:46]
  assign _GEN_1285 = 10'h140 == RADDR ? 10'h140 : _GEN_1284; // @[RAM_ST.scala 32:46]
  assign _GEN_1286 = 10'h141 == RADDR ? 10'h141 : _GEN_1285; // @[RAM_ST.scala 32:46]
  assign _GEN_1287 = 10'h142 == RADDR ? 10'h142 : _GEN_1286; // @[RAM_ST.scala 32:46]
  assign _GEN_1288 = 10'h143 == RADDR ? 10'h143 : _GEN_1287; // @[RAM_ST.scala 32:46]
  assign _GEN_1289 = 10'h144 == RADDR ? 10'h144 : _GEN_1288; // @[RAM_ST.scala 32:46]
  assign _GEN_1290 = 10'h145 == RADDR ? 10'h145 : _GEN_1289; // @[RAM_ST.scala 32:46]
  assign _GEN_1291 = 10'h146 == RADDR ? 10'h146 : _GEN_1290; // @[RAM_ST.scala 32:46]
  assign _GEN_1292 = 10'h147 == RADDR ? 10'h147 : _GEN_1291; // @[RAM_ST.scala 32:46]
  assign _GEN_1293 = 10'h148 == RADDR ? 10'h148 : _GEN_1292; // @[RAM_ST.scala 32:46]
  assign _GEN_1294 = 10'h149 == RADDR ? 10'h149 : _GEN_1293; // @[RAM_ST.scala 32:46]
  assign _GEN_1295 = 10'h14a == RADDR ? 10'h14a : _GEN_1294; // @[RAM_ST.scala 32:46]
  assign _GEN_1296 = 10'h14b == RADDR ? 10'h14b : _GEN_1295; // @[RAM_ST.scala 32:46]
  assign _GEN_1297 = 10'h14c == RADDR ? 10'h14c : _GEN_1296; // @[RAM_ST.scala 32:46]
  assign _GEN_1298 = 10'h14d == RADDR ? 10'h14d : _GEN_1297; // @[RAM_ST.scala 32:46]
  assign _GEN_1299 = 10'h14e == RADDR ? 10'h14e : _GEN_1298; // @[RAM_ST.scala 32:46]
  assign _GEN_1300 = 10'h14f == RADDR ? 10'h14f : _GEN_1299; // @[RAM_ST.scala 32:46]
  assign _GEN_1301 = 10'h150 == RADDR ? 10'h150 : _GEN_1300; // @[RAM_ST.scala 32:46]
  assign _GEN_1302 = 10'h151 == RADDR ? 10'h151 : _GEN_1301; // @[RAM_ST.scala 32:46]
  assign _GEN_1303 = 10'h152 == RADDR ? 10'h152 : _GEN_1302; // @[RAM_ST.scala 32:46]
  assign _GEN_1304 = 10'h153 == RADDR ? 10'h153 : _GEN_1303; // @[RAM_ST.scala 32:46]
  assign _GEN_1305 = 10'h154 == RADDR ? 10'h154 : _GEN_1304; // @[RAM_ST.scala 32:46]
  assign _GEN_1306 = 10'h155 == RADDR ? 10'h155 : _GEN_1305; // @[RAM_ST.scala 32:46]
  assign _GEN_1307 = 10'h156 == RADDR ? 10'h156 : _GEN_1306; // @[RAM_ST.scala 32:46]
  assign _GEN_1308 = 10'h157 == RADDR ? 10'h157 : _GEN_1307; // @[RAM_ST.scala 32:46]
  assign _GEN_1309 = 10'h158 == RADDR ? 10'h158 : _GEN_1308; // @[RAM_ST.scala 32:46]
  assign _GEN_1310 = 10'h159 == RADDR ? 10'h159 : _GEN_1309; // @[RAM_ST.scala 32:46]
  assign _GEN_1311 = 10'h15a == RADDR ? 10'h15a : _GEN_1310; // @[RAM_ST.scala 32:46]
  assign _GEN_1312 = 10'h15b == RADDR ? 10'h15b : _GEN_1311; // @[RAM_ST.scala 32:46]
  assign _GEN_1313 = 10'h15c == RADDR ? 10'h15c : _GEN_1312; // @[RAM_ST.scala 32:46]
  assign _GEN_1314 = 10'h15d == RADDR ? 10'h15d : _GEN_1313; // @[RAM_ST.scala 32:46]
  assign _GEN_1315 = 10'h15e == RADDR ? 10'h15e : _GEN_1314; // @[RAM_ST.scala 32:46]
  assign _GEN_1316 = 10'h15f == RADDR ? 10'h15f : _GEN_1315; // @[RAM_ST.scala 32:46]
  assign _GEN_1317 = 10'h160 == RADDR ? 10'h160 : _GEN_1316; // @[RAM_ST.scala 32:46]
  assign _GEN_1318 = 10'h161 == RADDR ? 10'h161 : _GEN_1317; // @[RAM_ST.scala 32:46]
  assign _GEN_1319 = 10'h162 == RADDR ? 10'h162 : _GEN_1318; // @[RAM_ST.scala 32:46]
  assign _GEN_1320 = 10'h163 == RADDR ? 10'h163 : _GEN_1319; // @[RAM_ST.scala 32:46]
  assign _GEN_1321 = 10'h164 == RADDR ? 10'h164 : _GEN_1320; // @[RAM_ST.scala 32:46]
  assign _GEN_1322 = 10'h165 == RADDR ? 10'h165 : _GEN_1321; // @[RAM_ST.scala 32:46]
  assign _GEN_1323 = 10'h166 == RADDR ? 10'h166 : _GEN_1322; // @[RAM_ST.scala 32:46]
  assign _GEN_1324 = 10'h167 == RADDR ? 10'h167 : _GEN_1323; // @[RAM_ST.scala 32:46]
  assign _GEN_1325 = 10'h168 == RADDR ? 10'h168 : _GEN_1324; // @[RAM_ST.scala 32:46]
  assign _GEN_1326 = 10'h169 == RADDR ? 10'h169 : _GEN_1325; // @[RAM_ST.scala 32:46]
  assign _GEN_1327 = 10'h16a == RADDR ? 10'h16a : _GEN_1326; // @[RAM_ST.scala 32:46]
  assign _GEN_1328 = 10'h16b == RADDR ? 10'h16b : _GEN_1327; // @[RAM_ST.scala 32:46]
  assign _GEN_1329 = 10'h16c == RADDR ? 10'h16c : _GEN_1328; // @[RAM_ST.scala 32:46]
  assign _GEN_1330 = 10'h16d == RADDR ? 10'h16d : _GEN_1329; // @[RAM_ST.scala 32:46]
  assign _GEN_1331 = 10'h16e == RADDR ? 10'h16e : _GEN_1330; // @[RAM_ST.scala 32:46]
  assign _GEN_1332 = 10'h16f == RADDR ? 10'h16f : _GEN_1331; // @[RAM_ST.scala 32:46]
  assign _GEN_1333 = 10'h170 == RADDR ? 10'h170 : _GEN_1332; // @[RAM_ST.scala 32:46]
  assign _GEN_1334 = 10'h171 == RADDR ? 10'h171 : _GEN_1333; // @[RAM_ST.scala 32:46]
  assign _GEN_1335 = 10'h172 == RADDR ? 10'h172 : _GEN_1334; // @[RAM_ST.scala 32:46]
  assign _GEN_1336 = 10'h173 == RADDR ? 10'h173 : _GEN_1335; // @[RAM_ST.scala 32:46]
  assign _GEN_1337 = 10'h174 == RADDR ? 10'h174 : _GEN_1336; // @[RAM_ST.scala 32:46]
  assign _GEN_1338 = 10'h175 == RADDR ? 10'h175 : _GEN_1337; // @[RAM_ST.scala 32:46]
  assign _GEN_1339 = 10'h176 == RADDR ? 10'h176 : _GEN_1338; // @[RAM_ST.scala 32:46]
  assign _GEN_1340 = 10'h177 == RADDR ? 10'h177 : _GEN_1339; // @[RAM_ST.scala 32:46]
  assign _GEN_1341 = 10'h178 == RADDR ? 10'h178 : _GEN_1340; // @[RAM_ST.scala 32:46]
  assign _GEN_1342 = 10'h179 == RADDR ? 10'h179 : _GEN_1341; // @[RAM_ST.scala 32:46]
  assign _GEN_1343 = 10'h17a == RADDR ? 10'h17a : _GEN_1342; // @[RAM_ST.scala 32:46]
  assign _GEN_1344 = 10'h17b == RADDR ? 10'h17b : _GEN_1343; // @[RAM_ST.scala 32:46]
  assign _GEN_1345 = 10'h17c == RADDR ? 10'h17c : _GEN_1344; // @[RAM_ST.scala 32:46]
  assign _GEN_1346 = 10'h17d == RADDR ? 10'h17d : _GEN_1345; // @[RAM_ST.scala 32:46]
  assign _GEN_1347 = 10'h17e == RADDR ? 10'h17e : _GEN_1346; // @[RAM_ST.scala 32:46]
  assign _GEN_1348 = 10'h17f == RADDR ? 10'h17f : _GEN_1347; // @[RAM_ST.scala 32:46]
  assign _GEN_1349 = 10'h180 == RADDR ? 10'h180 : _GEN_1348; // @[RAM_ST.scala 32:46]
  assign _GEN_1350 = 10'h181 == RADDR ? 10'h181 : _GEN_1349; // @[RAM_ST.scala 32:46]
  assign _GEN_1351 = 10'h182 == RADDR ? 10'h182 : _GEN_1350; // @[RAM_ST.scala 32:46]
  assign _GEN_1352 = 10'h183 == RADDR ? 10'h183 : _GEN_1351; // @[RAM_ST.scala 32:46]
  assign _GEN_1353 = 10'h184 == RADDR ? 10'h184 : _GEN_1352; // @[RAM_ST.scala 32:46]
  assign _GEN_1354 = 10'h185 == RADDR ? 10'h185 : _GEN_1353; // @[RAM_ST.scala 32:46]
  assign _GEN_1355 = 10'h186 == RADDR ? 10'h186 : _GEN_1354; // @[RAM_ST.scala 32:46]
  assign _GEN_1356 = 10'h187 == RADDR ? 10'h187 : _GEN_1355; // @[RAM_ST.scala 32:46]
  assign _GEN_1357 = 10'h188 == RADDR ? 10'h188 : _GEN_1356; // @[RAM_ST.scala 32:46]
  assign _GEN_1358 = 10'h189 == RADDR ? 10'h189 : _GEN_1357; // @[RAM_ST.scala 32:46]
  assign _GEN_1359 = 10'h18a == RADDR ? 10'h18a : _GEN_1358; // @[RAM_ST.scala 32:46]
  assign _GEN_1360 = 10'h18b == RADDR ? 10'h18b : _GEN_1359; // @[RAM_ST.scala 32:46]
  assign _GEN_1361 = 10'h18c == RADDR ? 10'h18c : _GEN_1360; // @[RAM_ST.scala 32:46]
  assign _GEN_1362 = 10'h18d == RADDR ? 10'h18d : _GEN_1361; // @[RAM_ST.scala 32:46]
  assign _GEN_1363 = 10'h18e == RADDR ? 10'h18e : _GEN_1362; // @[RAM_ST.scala 32:46]
  assign _GEN_1364 = 10'h18f == RADDR ? 10'h18f : _GEN_1363; // @[RAM_ST.scala 32:46]
  assign _GEN_1365 = 10'h190 == RADDR ? 10'h190 : _GEN_1364; // @[RAM_ST.scala 32:46]
  assign _GEN_1366 = 10'h191 == RADDR ? 10'h191 : _GEN_1365; // @[RAM_ST.scala 32:46]
  assign _GEN_1367 = 10'h192 == RADDR ? 10'h192 : _GEN_1366; // @[RAM_ST.scala 32:46]
  assign _GEN_1368 = 10'h193 == RADDR ? 10'h193 : _GEN_1367; // @[RAM_ST.scala 32:46]
  assign _GEN_1369 = 10'h194 == RADDR ? 10'h194 : _GEN_1368; // @[RAM_ST.scala 32:46]
  assign _GEN_1370 = 10'h195 == RADDR ? 10'h195 : _GEN_1369; // @[RAM_ST.scala 32:46]
  assign _GEN_1371 = 10'h196 == RADDR ? 10'h196 : _GEN_1370; // @[RAM_ST.scala 32:46]
  assign _GEN_1372 = 10'h197 == RADDR ? 10'h197 : _GEN_1371; // @[RAM_ST.scala 32:46]
  assign _GEN_1373 = 10'h198 == RADDR ? 10'h198 : _GEN_1372; // @[RAM_ST.scala 32:46]
  assign _GEN_1374 = 10'h199 == RADDR ? 10'h199 : _GEN_1373; // @[RAM_ST.scala 32:46]
  assign _GEN_1375 = 10'h19a == RADDR ? 10'h19a : _GEN_1374; // @[RAM_ST.scala 32:46]
  assign _GEN_1376 = 10'h19b == RADDR ? 10'h19b : _GEN_1375; // @[RAM_ST.scala 32:46]
  assign _GEN_1377 = 10'h19c == RADDR ? 10'h19c : _GEN_1376; // @[RAM_ST.scala 32:46]
  assign _GEN_1378 = 10'h19d == RADDR ? 10'h19d : _GEN_1377; // @[RAM_ST.scala 32:46]
  assign _GEN_1379 = 10'h19e == RADDR ? 10'h19e : _GEN_1378; // @[RAM_ST.scala 32:46]
  assign _GEN_1380 = 10'h19f == RADDR ? 10'h19f : _GEN_1379; // @[RAM_ST.scala 32:46]
  assign _GEN_1381 = 10'h1a0 == RADDR ? 10'h1a0 : _GEN_1380; // @[RAM_ST.scala 32:46]
  assign _GEN_1382 = 10'h1a1 == RADDR ? 10'h1a1 : _GEN_1381; // @[RAM_ST.scala 32:46]
  assign _GEN_1383 = 10'h1a2 == RADDR ? 10'h1a2 : _GEN_1382; // @[RAM_ST.scala 32:46]
  assign _GEN_1384 = 10'h1a3 == RADDR ? 10'h1a3 : _GEN_1383; // @[RAM_ST.scala 32:46]
  assign _GEN_1385 = 10'h1a4 == RADDR ? 10'h1a4 : _GEN_1384; // @[RAM_ST.scala 32:46]
  assign _GEN_1386 = 10'h1a5 == RADDR ? 10'h1a5 : _GEN_1385; // @[RAM_ST.scala 32:46]
  assign _GEN_1387 = 10'h1a6 == RADDR ? 10'h1a6 : _GEN_1386; // @[RAM_ST.scala 32:46]
  assign _GEN_1388 = 10'h1a7 == RADDR ? 10'h1a7 : _GEN_1387; // @[RAM_ST.scala 32:46]
  assign _GEN_1389 = 10'h1a8 == RADDR ? 10'h1a8 : _GEN_1388; // @[RAM_ST.scala 32:46]
  assign _GEN_1390 = 10'h1a9 == RADDR ? 10'h1a9 : _GEN_1389; // @[RAM_ST.scala 32:46]
  assign _GEN_1391 = 10'h1aa == RADDR ? 10'h1aa : _GEN_1390; // @[RAM_ST.scala 32:46]
  assign _GEN_1392 = 10'h1ab == RADDR ? 10'h1ab : _GEN_1391; // @[RAM_ST.scala 32:46]
  assign _GEN_1393 = 10'h1ac == RADDR ? 10'h1ac : _GEN_1392; // @[RAM_ST.scala 32:46]
  assign _GEN_1394 = 10'h1ad == RADDR ? 10'h1ad : _GEN_1393; // @[RAM_ST.scala 32:46]
  assign _GEN_1395 = 10'h1ae == RADDR ? 10'h1ae : _GEN_1394; // @[RAM_ST.scala 32:46]
  assign _GEN_1396 = 10'h1af == RADDR ? 10'h1af : _GEN_1395; // @[RAM_ST.scala 32:46]
  assign _GEN_1397 = 10'h1b0 == RADDR ? 10'h1b0 : _GEN_1396; // @[RAM_ST.scala 32:46]
  assign _GEN_1398 = 10'h1b1 == RADDR ? 10'h1b1 : _GEN_1397; // @[RAM_ST.scala 32:46]
  assign _GEN_1399 = 10'h1b2 == RADDR ? 10'h1b2 : _GEN_1398; // @[RAM_ST.scala 32:46]
  assign _GEN_1400 = 10'h1b3 == RADDR ? 10'h1b3 : _GEN_1399; // @[RAM_ST.scala 32:46]
  assign _GEN_1401 = 10'h1b4 == RADDR ? 10'h1b4 : _GEN_1400; // @[RAM_ST.scala 32:46]
  assign _GEN_1402 = 10'h1b5 == RADDR ? 10'h1b5 : _GEN_1401; // @[RAM_ST.scala 32:46]
  assign _GEN_1403 = 10'h1b6 == RADDR ? 10'h1b6 : _GEN_1402; // @[RAM_ST.scala 32:46]
  assign _GEN_1404 = 10'h1b7 == RADDR ? 10'h1b7 : _GEN_1403; // @[RAM_ST.scala 32:46]
  assign _GEN_1405 = 10'h1b8 == RADDR ? 10'h1b8 : _GEN_1404; // @[RAM_ST.scala 32:46]
  assign _GEN_1406 = 10'h1b9 == RADDR ? 10'h1b9 : _GEN_1405; // @[RAM_ST.scala 32:46]
  assign _GEN_1407 = 10'h1ba == RADDR ? 10'h1ba : _GEN_1406; // @[RAM_ST.scala 32:46]
  assign _GEN_1408 = 10'h1bb == RADDR ? 10'h1bb : _GEN_1407; // @[RAM_ST.scala 32:46]
  assign _GEN_1409 = 10'h1bc == RADDR ? 10'h1bc : _GEN_1408; // @[RAM_ST.scala 32:46]
  assign _GEN_1410 = 10'h1bd == RADDR ? 10'h1bd : _GEN_1409; // @[RAM_ST.scala 32:46]
  assign _GEN_1411 = 10'h1be == RADDR ? 10'h1be : _GEN_1410; // @[RAM_ST.scala 32:46]
  assign _GEN_1412 = 10'h1bf == RADDR ? 10'h1bf : _GEN_1411; // @[RAM_ST.scala 32:46]
  assign _GEN_1413 = 10'h1c0 == RADDR ? 10'h1c0 : _GEN_1412; // @[RAM_ST.scala 32:46]
  assign _GEN_1414 = 10'h1c1 == RADDR ? 10'h1c1 : _GEN_1413; // @[RAM_ST.scala 32:46]
  assign _GEN_1415 = 10'h1c2 == RADDR ? 10'h1c2 : _GEN_1414; // @[RAM_ST.scala 32:46]
  assign _GEN_1416 = 10'h1c3 == RADDR ? 10'h1c3 : _GEN_1415; // @[RAM_ST.scala 32:46]
  assign _GEN_1417 = 10'h1c4 == RADDR ? 10'h1c4 : _GEN_1416; // @[RAM_ST.scala 32:46]
  assign _GEN_1418 = 10'h1c5 == RADDR ? 10'h1c5 : _GEN_1417; // @[RAM_ST.scala 32:46]
  assign _GEN_1419 = 10'h1c6 == RADDR ? 10'h1c6 : _GEN_1418; // @[RAM_ST.scala 32:46]
  assign _GEN_1420 = 10'h1c7 == RADDR ? 10'h1c7 : _GEN_1419; // @[RAM_ST.scala 32:46]
  assign _GEN_1421 = 10'h1c8 == RADDR ? 10'h1c8 : _GEN_1420; // @[RAM_ST.scala 32:46]
  assign _GEN_1422 = 10'h1c9 == RADDR ? 10'h1c9 : _GEN_1421; // @[RAM_ST.scala 32:46]
  assign _GEN_1423 = 10'h1ca == RADDR ? 10'h1ca : _GEN_1422; // @[RAM_ST.scala 32:46]
  assign _GEN_1424 = 10'h1cb == RADDR ? 10'h1cb : _GEN_1423; // @[RAM_ST.scala 32:46]
  assign _GEN_1425 = 10'h1cc == RADDR ? 10'h1cc : _GEN_1424; // @[RAM_ST.scala 32:46]
  assign _GEN_1426 = 10'h1cd == RADDR ? 10'h1cd : _GEN_1425; // @[RAM_ST.scala 32:46]
  assign _GEN_1427 = 10'h1ce == RADDR ? 10'h1ce : _GEN_1426; // @[RAM_ST.scala 32:46]
  assign _GEN_1428 = 10'h1cf == RADDR ? 10'h1cf : _GEN_1427; // @[RAM_ST.scala 32:46]
  assign _GEN_1429 = 10'h1d0 == RADDR ? 10'h1d0 : _GEN_1428; // @[RAM_ST.scala 32:46]
  assign _GEN_1430 = 10'h1d1 == RADDR ? 10'h1d1 : _GEN_1429; // @[RAM_ST.scala 32:46]
  assign _GEN_1431 = 10'h1d2 == RADDR ? 10'h1d2 : _GEN_1430; // @[RAM_ST.scala 32:46]
  assign _GEN_1432 = 10'h1d3 == RADDR ? 10'h1d3 : _GEN_1431; // @[RAM_ST.scala 32:46]
  assign _GEN_1433 = 10'h1d4 == RADDR ? 10'h1d4 : _GEN_1432; // @[RAM_ST.scala 32:46]
  assign _GEN_1434 = 10'h1d5 == RADDR ? 10'h1d5 : _GEN_1433; // @[RAM_ST.scala 32:46]
  assign _GEN_1435 = 10'h1d6 == RADDR ? 10'h1d6 : _GEN_1434; // @[RAM_ST.scala 32:46]
  assign _GEN_1436 = 10'h1d7 == RADDR ? 10'h1d7 : _GEN_1435; // @[RAM_ST.scala 32:46]
  assign _GEN_1437 = 10'h1d8 == RADDR ? 10'h1d8 : _GEN_1436; // @[RAM_ST.scala 32:46]
  assign _GEN_1438 = 10'h1d9 == RADDR ? 10'h1d9 : _GEN_1437; // @[RAM_ST.scala 32:46]
  assign _GEN_1439 = 10'h1da == RADDR ? 10'h1da : _GEN_1438; // @[RAM_ST.scala 32:46]
  assign _GEN_1440 = 10'h1db == RADDR ? 10'h1db : _GEN_1439; // @[RAM_ST.scala 32:46]
  assign _GEN_1441 = 10'h1dc == RADDR ? 10'h1dc : _GEN_1440; // @[RAM_ST.scala 32:46]
  assign _GEN_1442 = 10'h1dd == RADDR ? 10'h1dd : _GEN_1441; // @[RAM_ST.scala 32:46]
  assign _GEN_1443 = 10'h1de == RADDR ? 10'h1de : _GEN_1442; // @[RAM_ST.scala 32:46]
  assign _GEN_1444 = 10'h1df == RADDR ? 10'h1df : _GEN_1443; // @[RAM_ST.scala 32:46]
  assign _GEN_1445 = 10'h1e0 == RADDR ? 10'h1e0 : _GEN_1444; // @[RAM_ST.scala 32:46]
  assign _GEN_1446 = 10'h1e1 == RADDR ? 10'h1e1 : _GEN_1445; // @[RAM_ST.scala 32:46]
  assign _GEN_1447 = 10'h1e2 == RADDR ? 10'h1e2 : _GEN_1446; // @[RAM_ST.scala 32:46]
  assign _GEN_1448 = 10'h1e3 == RADDR ? 10'h1e3 : _GEN_1447; // @[RAM_ST.scala 32:46]
  assign _GEN_1449 = 10'h1e4 == RADDR ? 10'h1e4 : _GEN_1448; // @[RAM_ST.scala 32:46]
  assign _GEN_1450 = 10'h1e5 == RADDR ? 10'h1e5 : _GEN_1449; // @[RAM_ST.scala 32:46]
  assign _GEN_1451 = 10'h1e6 == RADDR ? 10'h1e6 : _GEN_1450; // @[RAM_ST.scala 32:46]
  assign _GEN_1452 = 10'h1e7 == RADDR ? 10'h1e7 : _GEN_1451; // @[RAM_ST.scala 32:46]
  assign _GEN_1453 = 10'h1e8 == RADDR ? 10'h1e8 : _GEN_1452; // @[RAM_ST.scala 32:46]
  assign _GEN_1454 = 10'h1e9 == RADDR ? 10'h1e9 : _GEN_1453; // @[RAM_ST.scala 32:46]
  assign _GEN_1455 = 10'h1ea == RADDR ? 10'h1ea : _GEN_1454; // @[RAM_ST.scala 32:46]
  assign _GEN_1456 = 10'h1eb == RADDR ? 10'h1eb : _GEN_1455; // @[RAM_ST.scala 32:46]
  assign _GEN_1457 = 10'h1ec == RADDR ? 10'h1ec : _GEN_1456; // @[RAM_ST.scala 32:46]
  assign _GEN_1458 = 10'h1ed == RADDR ? 10'h1ed : _GEN_1457; // @[RAM_ST.scala 32:46]
  assign _GEN_1459 = 10'h1ee == RADDR ? 10'h1ee : _GEN_1458; // @[RAM_ST.scala 32:46]
  assign _GEN_1460 = 10'h1ef == RADDR ? 10'h1ef : _GEN_1459; // @[RAM_ST.scala 32:46]
  assign _GEN_1461 = 10'h1f0 == RADDR ? 10'h1f0 : _GEN_1460; // @[RAM_ST.scala 32:46]
  assign _GEN_1462 = 10'h1f1 == RADDR ? 10'h1f1 : _GEN_1461; // @[RAM_ST.scala 32:46]
  assign _GEN_1463 = 10'h1f2 == RADDR ? 10'h1f2 : _GEN_1462; // @[RAM_ST.scala 32:46]
  assign _GEN_1464 = 10'h1f3 == RADDR ? 10'h1f3 : _GEN_1463; // @[RAM_ST.scala 32:46]
  assign _GEN_1465 = 10'h1f4 == RADDR ? 10'h1f4 : _GEN_1464; // @[RAM_ST.scala 32:46]
  assign _GEN_1466 = 10'h1f5 == RADDR ? 10'h1f5 : _GEN_1465; // @[RAM_ST.scala 32:46]
  assign _GEN_1467 = 10'h1f6 == RADDR ? 10'h1f6 : _GEN_1466; // @[RAM_ST.scala 32:46]
  assign _GEN_1468 = 10'h1f7 == RADDR ? 10'h1f7 : _GEN_1467; // @[RAM_ST.scala 32:46]
  assign _GEN_1469 = 10'h1f8 == RADDR ? 10'h1f8 : _GEN_1468; // @[RAM_ST.scala 32:46]
  assign _GEN_1470 = 10'h1f9 == RADDR ? 10'h1f9 : _GEN_1469; // @[RAM_ST.scala 32:46]
  assign _GEN_1471 = 10'h1fa == RADDR ? 10'h1fa : _GEN_1470; // @[RAM_ST.scala 32:46]
  assign _GEN_1472 = 10'h1fb == RADDR ? 10'h1fb : _GEN_1471; // @[RAM_ST.scala 32:46]
  assign _GEN_1473 = 10'h1fc == RADDR ? 10'h1fc : _GEN_1472; // @[RAM_ST.scala 32:46]
  assign _GEN_1474 = 10'h1fd == RADDR ? 10'h1fd : _GEN_1473; // @[RAM_ST.scala 32:46]
  assign _GEN_1475 = 10'h1fe == RADDR ? 10'h1fe : _GEN_1474; // @[RAM_ST.scala 32:46]
  assign _GEN_1476 = 10'h1ff == RADDR ? 10'h1ff : _GEN_1475; // @[RAM_ST.scala 32:46]
  assign _GEN_1477 = 10'h200 == RADDR ? 10'h200 : _GEN_1476; // @[RAM_ST.scala 32:46]
  assign _GEN_1478 = 10'h201 == RADDR ? 10'h201 : _GEN_1477; // @[RAM_ST.scala 32:46]
  assign _GEN_1479 = 10'h202 == RADDR ? 10'h202 : _GEN_1478; // @[RAM_ST.scala 32:46]
  assign _GEN_1480 = 10'h203 == RADDR ? 10'h203 : _GEN_1479; // @[RAM_ST.scala 32:46]
  assign _GEN_1481 = 10'h204 == RADDR ? 10'h204 : _GEN_1480; // @[RAM_ST.scala 32:46]
  assign _GEN_1482 = 10'h205 == RADDR ? 10'h205 : _GEN_1481; // @[RAM_ST.scala 32:46]
  assign _GEN_1483 = 10'h206 == RADDR ? 10'h206 : _GEN_1482; // @[RAM_ST.scala 32:46]
  assign _GEN_1484 = 10'h207 == RADDR ? 10'h207 : _GEN_1483; // @[RAM_ST.scala 32:46]
  assign _GEN_1485 = 10'h208 == RADDR ? 10'h208 : _GEN_1484; // @[RAM_ST.scala 32:46]
  assign _GEN_1486 = 10'h209 == RADDR ? 10'h209 : _GEN_1485; // @[RAM_ST.scala 32:46]
  assign _GEN_1487 = 10'h20a == RADDR ? 10'h20a : _GEN_1486; // @[RAM_ST.scala 32:46]
  assign _GEN_1488 = 10'h20b == RADDR ? 10'h20b : _GEN_1487; // @[RAM_ST.scala 32:46]
  assign _GEN_1489 = 10'h20c == RADDR ? 10'h20c : _GEN_1488; // @[RAM_ST.scala 32:46]
  assign _GEN_1490 = 10'h20d == RADDR ? 10'h20d : _GEN_1489; // @[RAM_ST.scala 32:46]
  assign _GEN_1491 = 10'h20e == RADDR ? 10'h20e : _GEN_1490; // @[RAM_ST.scala 32:46]
  assign _GEN_1492 = 10'h20f == RADDR ? 10'h20f : _GEN_1491; // @[RAM_ST.scala 32:46]
  assign _GEN_1493 = 10'h210 == RADDR ? 10'h210 : _GEN_1492; // @[RAM_ST.scala 32:46]
  assign _GEN_1494 = 10'h211 == RADDR ? 10'h211 : _GEN_1493; // @[RAM_ST.scala 32:46]
  assign _GEN_1495 = 10'h212 == RADDR ? 10'h212 : _GEN_1494; // @[RAM_ST.scala 32:46]
  assign _GEN_1496 = 10'h213 == RADDR ? 10'h213 : _GEN_1495; // @[RAM_ST.scala 32:46]
  assign _GEN_1497 = 10'h214 == RADDR ? 10'h214 : _GEN_1496; // @[RAM_ST.scala 32:46]
  assign _GEN_1498 = 10'h215 == RADDR ? 10'h215 : _GEN_1497; // @[RAM_ST.scala 32:46]
  assign _GEN_1499 = 10'h216 == RADDR ? 10'h216 : _GEN_1498; // @[RAM_ST.scala 32:46]
  assign _GEN_1500 = 10'h217 == RADDR ? 10'h217 : _GEN_1499; // @[RAM_ST.scala 32:46]
  assign _GEN_1501 = 10'h218 == RADDR ? 10'h218 : _GEN_1500; // @[RAM_ST.scala 32:46]
  assign _GEN_1502 = 10'h219 == RADDR ? 10'h219 : _GEN_1501; // @[RAM_ST.scala 32:46]
  assign _GEN_1503 = 10'h21a == RADDR ? 10'h21a : _GEN_1502; // @[RAM_ST.scala 32:46]
  assign _GEN_1504 = 10'h21b == RADDR ? 10'h21b : _GEN_1503; // @[RAM_ST.scala 32:46]
  assign _GEN_1505 = 10'h21c == RADDR ? 10'h21c : _GEN_1504; // @[RAM_ST.scala 32:46]
  assign _GEN_1506 = 10'h21d == RADDR ? 10'h21d : _GEN_1505; // @[RAM_ST.scala 32:46]
  assign _GEN_1507 = 10'h21e == RADDR ? 10'h21e : _GEN_1506; // @[RAM_ST.scala 32:46]
  assign _GEN_1508 = 10'h21f == RADDR ? 10'h21f : _GEN_1507; // @[RAM_ST.scala 32:46]
  assign _GEN_1509 = 10'h220 == RADDR ? 10'h220 : _GEN_1508; // @[RAM_ST.scala 32:46]
  assign _GEN_1510 = 10'h221 == RADDR ? 10'h221 : _GEN_1509; // @[RAM_ST.scala 32:46]
  assign _GEN_1511 = 10'h222 == RADDR ? 10'h222 : _GEN_1510; // @[RAM_ST.scala 32:46]
  assign _GEN_1512 = 10'h223 == RADDR ? 10'h223 : _GEN_1511; // @[RAM_ST.scala 32:46]
  assign _GEN_1513 = 10'h224 == RADDR ? 10'h224 : _GEN_1512; // @[RAM_ST.scala 32:46]
  assign _GEN_1514 = 10'h225 == RADDR ? 10'h225 : _GEN_1513; // @[RAM_ST.scala 32:46]
  assign _GEN_1515 = 10'h226 == RADDR ? 10'h226 : _GEN_1514; // @[RAM_ST.scala 32:46]
  assign _GEN_1516 = 10'h227 == RADDR ? 10'h227 : _GEN_1515; // @[RAM_ST.scala 32:46]
  assign _GEN_1517 = 10'h228 == RADDR ? 10'h228 : _GEN_1516; // @[RAM_ST.scala 32:46]
  assign _GEN_1518 = 10'h229 == RADDR ? 10'h229 : _GEN_1517; // @[RAM_ST.scala 32:46]
  assign _GEN_1519 = 10'h22a == RADDR ? 10'h22a : _GEN_1518; // @[RAM_ST.scala 32:46]
  assign _GEN_1520 = 10'h22b == RADDR ? 10'h22b : _GEN_1519; // @[RAM_ST.scala 32:46]
  assign _GEN_1521 = 10'h22c == RADDR ? 10'h22c : _GEN_1520; // @[RAM_ST.scala 32:46]
  assign _GEN_1522 = 10'h22d == RADDR ? 10'h22d : _GEN_1521; // @[RAM_ST.scala 32:46]
  assign _GEN_1523 = 10'h22e == RADDR ? 10'h22e : _GEN_1522; // @[RAM_ST.scala 32:46]
  assign _GEN_1524 = 10'h22f == RADDR ? 10'h22f : _GEN_1523; // @[RAM_ST.scala 32:46]
  assign _GEN_1525 = 10'h230 == RADDR ? 10'h230 : _GEN_1524; // @[RAM_ST.scala 32:46]
  assign _GEN_1526 = 10'h231 == RADDR ? 10'h231 : _GEN_1525; // @[RAM_ST.scala 32:46]
  assign _GEN_1527 = 10'h232 == RADDR ? 10'h232 : _GEN_1526; // @[RAM_ST.scala 32:46]
  assign _GEN_1528 = 10'h233 == RADDR ? 10'h233 : _GEN_1527; // @[RAM_ST.scala 32:46]
  assign _GEN_1529 = 10'h234 == RADDR ? 10'h234 : _GEN_1528; // @[RAM_ST.scala 32:46]
  assign _GEN_1530 = 10'h235 == RADDR ? 10'h235 : _GEN_1529; // @[RAM_ST.scala 32:46]
  assign _GEN_1531 = 10'h236 == RADDR ? 10'h236 : _GEN_1530; // @[RAM_ST.scala 32:46]
  assign _GEN_1532 = 10'h237 == RADDR ? 10'h237 : _GEN_1531; // @[RAM_ST.scala 32:46]
  assign _GEN_1533 = 10'h238 == RADDR ? 10'h238 : _GEN_1532; // @[RAM_ST.scala 32:46]
  assign _GEN_1534 = 10'h239 == RADDR ? 10'h239 : _GEN_1533; // @[RAM_ST.scala 32:46]
  assign _GEN_1535 = 10'h23a == RADDR ? 10'h23a : _GEN_1534; // @[RAM_ST.scala 32:46]
  assign _GEN_1536 = 10'h23b == RADDR ? 10'h23b : _GEN_1535; // @[RAM_ST.scala 32:46]
  assign _GEN_1537 = 10'h23c == RADDR ? 10'h23c : _GEN_1536; // @[RAM_ST.scala 32:46]
  assign _GEN_1538 = 10'h23d == RADDR ? 10'h23d : _GEN_1537; // @[RAM_ST.scala 32:46]
  assign _GEN_1539 = 10'h23e == RADDR ? 10'h23e : _GEN_1538; // @[RAM_ST.scala 32:46]
  assign _GEN_1540 = 10'h23f == RADDR ? 10'h23f : _GEN_1539; // @[RAM_ST.scala 32:46]
  assign _GEN_1541 = 10'h240 == RADDR ? 10'h240 : _GEN_1540; // @[RAM_ST.scala 32:46]
  assign _GEN_1542 = 10'h241 == RADDR ? 10'h241 : _GEN_1541; // @[RAM_ST.scala 32:46]
  assign _GEN_1543 = 10'h242 == RADDR ? 10'h242 : _GEN_1542; // @[RAM_ST.scala 32:46]
  assign _GEN_1544 = 10'h243 == RADDR ? 10'h243 : _GEN_1543; // @[RAM_ST.scala 32:46]
  assign _GEN_1545 = 10'h244 == RADDR ? 10'h244 : _GEN_1544; // @[RAM_ST.scala 32:46]
  assign _GEN_1546 = 10'h245 == RADDR ? 10'h245 : _GEN_1545; // @[RAM_ST.scala 32:46]
  assign _GEN_1547 = 10'h246 == RADDR ? 10'h246 : _GEN_1546; // @[RAM_ST.scala 32:46]
  assign _GEN_1548 = 10'h247 == RADDR ? 10'h247 : _GEN_1547; // @[RAM_ST.scala 32:46]
  assign _GEN_1549 = 10'h248 == RADDR ? 10'h248 : _GEN_1548; // @[RAM_ST.scala 32:46]
  assign _GEN_1550 = 10'h249 == RADDR ? 10'h249 : _GEN_1549; // @[RAM_ST.scala 32:46]
  assign _GEN_1551 = 10'h24a == RADDR ? 10'h24a : _GEN_1550; // @[RAM_ST.scala 32:46]
  assign _GEN_1552 = 10'h24b == RADDR ? 10'h24b : _GEN_1551; // @[RAM_ST.scala 32:46]
  assign _GEN_1553 = 10'h24c == RADDR ? 10'h24c : _GEN_1552; // @[RAM_ST.scala 32:46]
  assign _GEN_1554 = 10'h24d == RADDR ? 10'h24d : _GEN_1553; // @[RAM_ST.scala 32:46]
  assign _GEN_1555 = 10'h24e == RADDR ? 10'h24e : _GEN_1554; // @[RAM_ST.scala 32:46]
  assign _GEN_1556 = 10'h24f == RADDR ? 10'h24f : _GEN_1555; // @[RAM_ST.scala 32:46]
  assign _GEN_1557 = 10'h250 == RADDR ? 10'h250 : _GEN_1556; // @[RAM_ST.scala 32:46]
  assign _GEN_1558 = 10'h251 == RADDR ? 10'h251 : _GEN_1557; // @[RAM_ST.scala 32:46]
  assign _GEN_1559 = 10'h252 == RADDR ? 10'h252 : _GEN_1558; // @[RAM_ST.scala 32:46]
  assign _GEN_1560 = 10'h253 == RADDR ? 10'h253 : _GEN_1559; // @[RAM_ST.scala 32:46]
  assign _GEN_1561 = 10'h254 == RADDR ? 10'h254 : _GEN_1560; // @[RAM_ST.scala 32:46]
  assign _GEN_1562 = 10'h255 == RADDR ? 10'h255 : _GEN_1561; // @[RAM_ST.scala 32:46]
  assign _GEN_1563 = 10'h256 == RADDR ? 10'h256 : _GEN_1562; // @[RAM_ST.scala 32:46]
  assign _GEN_1564 = 10'h257 == RADDR ? 10'h257 : _GEN_1563; // @[RAM_ST.scala 32:46]
  assign _GEN_1565 = 10'h258 == RADDR ? 10'h258 : _GEN_1564; // @[RAM_ST.scala 32:46]
  assign _GEN_1566 = 10'h259 == RADDR ? 10'h259 : _GEN_1565; // @[RAM_ST.scala 32:46]
  assign _GEN_1567 = 10'h25a == RADDR ? 10'h25a : _GEN_1566; // @[RAM_ST.scala 32:46]
  assign _GEN_1568 = 10'h25b == RADDR ? 10'h25b : _GEN_1567; // @[RAM_ST.scala 32:46]
  assign _GEN_1569 = 10'h25c == RADDR ? 10'h25c : _GEN_1568; // @[RAM_ST.scala 32:46]
  assign _GEN_1570 = 10'h25d == RADDR ? 10'h25d : _GEN_1569; // @[RAM_ST.scala 32:46]
  assign _GEN_1571 = 10'h25e == RADDR ? 10'h25e : _GEN_1570; // @[RAM_ST.scala 32:46]
  assign _GEN_1572 = 10'h25f == RADDR ? 10'h25f : _GEN_1571; // @[RAM_ST.scala 32:46]
  assign _GEN_1573 = 10'h260 == RADDR ? 10'h260 : _GEN_1572; // @[RAM_ST.scala 32:46]
  assign _GEN_1574 = 10'h261 == RADDR ? 10'h261 : _GEN_1573; // @[RAM_ST.scala 32:46]
  assign _GEN_1575 = 10'h262 == RADDR ? 10'h262 : _GEN_1574; // @[RAM_ST.scala 32:46]
  assign _GEN_1576 = 10'h263 == RADDR ? 10'h263 : _GEN_1575; // @[RAM_ST.scala 32:46]
  assign _GEN_1577 = 10'h264 == RADDR ? 10'h264 : _GEN_1576; // @[RAM_ST.scala 32:46]
  assign _GEN_1578 = 10'h265 == RADDR ? 10'h265 : _GEN_1577; // @[RAM_ST.scala 32:46]
  assign _GEN_1579 = 10'h266 == RADDR ? 10'h266 : _GEN_1578; // @[RAM_ST.scala 32:46]
  assign _GEN_1580 = 10'h267 == RADDR ? 10'h267 : _GEN_1579; // @[RAM_ST.scala 32:46]
  assign _GEN_1581 = 10'h268 == RADDR ? 10'h268 : _GEN_1580; // @[RAM_ST.scala 32:46]
  assign _GEN_1582 = 10'h269 == RADDR ? 10'h269 : _GEN_1581; // @[RAM_ST.scala 32:46]
  assign _GEN_1583 = 10'h26a == RADDR ? 10'h26a : _GEN_1582; // @[RAM_ST.scala 32:46]
  assign _GEN_1584 = 10'h26b == RADDR ? 10'h26b : _GEN_1583; // @[RAM_ST.scala 32:46]
  assign _GEN_1585 = 10'h26c == RADDR ? 10'h26c : _GEN_1584; // @[RAM_ST.scala 32:46]
  assign _GEN_1586 = 10'h26d == RADDR ? 10'h26d : _GEN_1585; // @[RAM_ST.scala 32:46]
  assign _GEN_1587 = 10'h26e == RADDR ? 10'h26e : _GEN_1586; // @[RAM_ST.scala 32:46]
  assign _GEN_1588 = 10'h26f == RADDR ? 10'h26f : _GEN_1587; // @[RAM_ST.scala 32:46]
  assign _GEN_1589 = 10'h270 == RADDR ? 10'h270 : _GEN_1588; // @[RAM_ST.scala 32:46]
  assign _GEN_1590 = 10'h271 == RADDR ? 10'h271 : _GEN_1589; // @[RAM_ST.scala 32:46]
  assign _GEN_1591 = 10'h272 == RADDR ? 10'h272 : _GEN_1590; // @[RAM_ST.scala 32:46]
  assign _GEN_1592 = 10'h273 == RADDR ? 10'h273 : _GEN_1591; // @[RAM_ST.scala 32:46]
  assign _GEN_1593 = 10'h274 == RADDR ? 10'h274 : _GEN_1592; // @[RAM_ST.scala 32:46]
  assign _GEN_1594 = 10'h275 == RADDR ? 10'h275 : _GEN_1593; // @[RAM_ST.scala 32:46]
  assign _GEN_1595 = 10'h276 == RADDR ? 10'h276 : _GEN_1594; // @[RAM_ST.scala 32:46]
  assign _GEN_1596 = 10'h277 == RADDR ? 10'h277 : _GEN_1595; // @[RAM_ST.scala 32:46]
  assign _GEN_1597 = 10'h278 == RADDR ? 10'h278 : _GEN_1596; // @[RAM_ST.scala 32:46]
  assign _GEN_1598 = 10'h279 == RADDR ? 10'h279 : _GEN_1597; // @[RAM_ST.scala 32:46]
  assign _GEN_1599 = 10'h27a == RADDR ? 10'h27a : _GEN_1598; // @[RAM_ST.scala 32:46]
  assign _GEN_1600 = 10'h27b == RADDR ? 10'h27b : _GEN_1599; // @[RAM_ST.scala 32:46]
  assign _GEN_1601 = 10'h27c == RADDR ? 10'h27c : _GEN_1600; // @[RAM_ST.scala 32:46]
  assign _GEN_1602 = 10'h27d == RADDR ? 10'h27d : _GEN_1601; // @[RAM_ST.scala 32:46]
  assign _GEN_1603 = 10'h27e == RADDR ? 10'h27e : _GEN_1602; // @[RAM_ST.scala 32:46]
  assign _GEN_1604 = 10'h27f == RADDR ? 10'h27f : _GEN_1603; // @[RAM_ST.scala 32:46]
  assign _GEN_1605 = 10'h280 == RADDR ? 10'h280 : _GEN_1604; // @[RAM_ST.scala 32:46]
  assign _GEN_1606 = 10'h281 == RADDR ? 10'h281 : _GEN_1605; // @[RAM_ST.scala 32:46]
  assign _GEN_1607 = 10'h282 == RADDR ? 10'h282 : _GEN_1606; // @[RAM_ST.scala 32:46]
  assign _GEN_1608 = 10'h283 == RADDR ? 10'h283 : _GEN_1607; // @[RAM_ST.scala 32:46]
  assign _GEN_1609 = 10'h284 == RADDR ? 10'h284 : _GEN_1608; // @[RAM_ST.scala 32:46]
  assign _GEN_1610 = 10'h285 == RADDR ? 10'h285 : _GEN_1609; // @[RAM_ST.scala 32:46]
  assign _GEN_1611 = 10'h286 == RADDR ? 10'h286 : _GEN_1610; // @[RAM_ST.scala 32:46]
  assign _GEN_1612 = 10'h287 == RADDR ? 10'h287 : _GEN_1611; // @[RAM_ST.scala 32:46]
  assign _GEN_1613 = 10'h288 == RADDR ? 10'h288 : _GEN_1612; // @[RAM_ST.scala 32:46]
  assign _GEN_1614 = 10'h289 == RADDR ? 10'h289 : _GEN_1613; // @[RAM_ST.scala 32:46]
  assign _GEN_1615 = 10'h28a == RADDR ? 10'h28a : _GEN_1614; // @[RAM_ST.scala 32:46]
  assign _GEN_1616 = 10'h28b == RADDR ? 10'h28b : _GEN_1615; // @[RAM_ST.scala 32:46]
  assign _GEN_1617 = 10'h28c == RADDR ? 10'h28c : _GEN_1616; // @[RAM_ST.scala 32:46]
  assign _GEN_1618 = 10'h28d == RADDR ? 10'h28d : _GEN_1617; // @[RAM_ST.scala 32:46]
  assign _GEN_1619 = 10'h28e == RADDR ? 10'h28e : _GEN_1618; // @[RAM_ST.scala 32:46]
  assign _GEN_1620 = 10'h28f == RADDR ? 10'h28f : _GEN_1619; // @[RAM_ST.scala 32:46]
  assign _GEN_1621 = 10'h290 == RADDR ? 10'h290 : _GEN_1620; // @[RAM_ST.scala 32:46]
  assign _GEN_1622 = 10'h291 == RADDR ? 10'h291 : _GEN_1621; // @[RAM_ST.scala 32:46]
  assign _GEN_1623 = 10'h292 == RADDR ? 10'h292 : _GEN_1622; // @[RAM_ST.scala 32:46]
  assign _GEN_1624 = 10'h293 == RADDR ? 10'h293 : _GEN_1623; // @[RAM_ST.scala 32:46]
  assign _GEN_1625 = 10'h294 == RADDR ? 10'h294 : _GEN_1624; // @[RAM_ST.scala 32:46]
  assign _GEN_1626 = 10'h295 == RADDR ? 10'h295 : _GEN_1625; // @[RAM_ST.scala 32:46]
  assign _GEN_1627 = 10'h296 == RADDR ? 10'h296 : _GEN_1626; // @[RAM_ST.scala 32:46]
  assign _GEN_1628 = 10'h297 == RADDR ? 10'h297 : _GEN_1627; // @[RAM_ST.scala 32:46]
  assign _GEN_1629 = 10'h298 == RADDR ? 10'h298 : _GEN_1628; // @[RAM_ST.scala 32:46]
  assign _GEN_1630 = 10'h299 == RADDR ? 10'h299 : _GEN_1629; // @[RAM_ST.scala 32:46]
  assign _GEN_1631 = 10'h29a == RADDR ? 10'h29a : _GEN_1630; // @[RAM_ST.scala 32:46]
  assign _GEN_1632 = 10'h29b == RADDR ? 10'h29b : _GEN_1631; // @[RAM_ST.scala 32:46]
  assign _GEN_1633 = 10'h29c == RADDR ? 10'h29c : _GEN_1632; // @[RAM_ST.scala 32:46]
  assign _GEN_1634 = 10'h29d == RADDR ? 10'h29d : _GEN_1633; // @[RAM_ST.scala 32:46]
  assign _GEN_1635 = 10'h29e == RADDR ? 10'h29e : _GEN_1634; // @[RAM_ST.scala 32:46]
  assign _GEN_1636 = 10'h29f == RADDR ? 10'h29f : _GEN_1635; // @[RAM_ST.scala 32:46]
  assign _GEN_1637 = 10'h2a0 == RADDR ? 10'h2a0 : _GEN_1636; // @[RAM_ST.scala 32:46]
  assign _GEN_1638 = 10'h2a1 == RADDR ? 10'h2a1 : _GEN_1637; // @[RAM_ST.scala 32:46]
  assign _GEN_1639 = 10'h2a2 == RADDR ? 10'h2a2 : _GEN_1638; // @[RAM_ST.scala 32:46]
  assign _GEN_1640 = 10'h2a3 == RADDR ? 10'h2a3 : _GEN_1639; // @[RAM_ST.scala 32:46]
  assign _GEN_1641 = 10'h2a4 == RADDR ? 10'h2a4 : _GEN_1640; // @[RAM_ST.scala 32:46]
  assign _GEN_1642 = 10'h2a5 == RADDR ? 10'h2a5 : _GEN_1641; // @[RAM_ST.scala 32:46]
  assign _GEN_1643 = 10'h2a6 == RADDR ? 10'h2a6 : _GEN_1642; // @[RAM_ST.scala 32:46]
  assign _GEN_1644 = 10'h2a7 == RADDR ? 10'h2a7 : _GEN_1643; // @[RAM_ST.scala 32:46]
  assign _GEN_1645 = 10'h2a8 == RADDR ? 10'h2a8 : _GEN_1644; // @[RAM_ST.scala 32:46]
  assign _GEN_1646 = 10'h2a9 == RADDR ? 10'h2a9 : _GEN_1645; // @[RAM_ST.scala 32:46]
  assign _GEN_1647 = 10'h2aa == RADDR ? 10'h2aa : _GEN_1646; // @[RAM_ST.scala 32:46]
  assign _GEN_1648 = 10'h2ab == RADDR ? 10'h2ab : _GEN_1647; // @[RAM_ST.scala 32:46]
  assign _GEN_1649 = 10'h2ac == RADDR ? 10'h2ac : _GEN_1648; // @[RAM_ST.scala 32:46]
  assign _GEN_1650 = 10'h2ad == RADDR ? 10'h2ad : _GEN_1649; // @[RAM_ST.scala 32:46]
  assign _GEN_1651 = 10'h2ae == RADDR ? 10'h2ae : _GEN_1650; // @[RAM_ST.scala 32:46]
  assign _GEN_1652 = 10'h2af == RADDR ? 10'h2af : _GEN_1651; // @[RAM_ST.scala 32:46]
  assign _GEN_1653 = 10'h2b0 == RADDR ? 10'h2b0 : _GEN_1652; // @[RAM_ST.scala 32:46]
  assign _GEN_1654 = 10'h2b1 == RADDR ? 10'h2b1 : _GEN_1653; // @[RAM_ST.scala 32:46]
  assign _GEN_1655 = 10'h2b2 == RADDR ? 10'h2b2 : _GEN_1654; // @[RAM_ST.scala 32:46]
  assign _GEN_1656 = 10'h2b3 == RADDR ? 10'h2b3 : _GEN_1655; // @[RAM_ST.scala 32:46]
  assign _GEN_1657 = 10'h2b4 == RADDR ? 10'h2b4 : _GEN_1656; // @[RAM_ST.scala 32:46]
  assign _GEN_1658 = 10'h2b5 == RADDR ? 10'h2b5 : _GEN_1657; // @[RAM_ST.scala 32:46]
  assign _GEN_1659 = 10'h2b6 == RADDR ? 10'h2b6 : _GEN_1658; // @[RAM_ST.scala 32:46]
  assign _GEN_1660 = 10'h2b7 == RADDR ? 10'h2b7 : _GEN_1659; // @[RAM_ST.scala 32:46]
  assign _GEN_1661 = 10'h2b8 == RADDR ? 10'h2b8 : _GEN_1660; // @[RAM_ST.scala 32:46]
  assign _GEN_1662 = 10'h2b9 == RADDR ? 10'h2b9 : _GEN_1661; // @[RAM_ST.scala 32:46]
  assign _GEN_1663 = 10'h2ba == RADDR ? 10'h2ba : _GEN_1662; // @[RAM_ST.scala 32:46]
  assign _GEN_1664 = 10'h2bb == RADDR ? 10'h2bb : _GEN_1663; // @[RAM_ST.scala 32:46]
  assign _GEN_1665 = 10'h2bc == RADDR ? 10'h2bc : _GEN_1664; // @[RAM_ST.scala 32:46]
  assign _GEN_1666 = 10'h2bd == RADDR ? 10'h2bd : _GEN_1665; // @[RAM_ST.scala 32:46]
  assign _GEN_1667 = 10'h2be == RADDR ? 10'h2be : _GEN_1666; // @[RAM_ST.scala 32:46]
  assign _GEN_1668 = 10'h2bf == RADDR ? 10'h2bf : _GEN_1667; // @[RAM_ST.scala 32:46]
  assign _GEN_1669 = 10'h2c0 == RADDR ? 10'h2c0 : _GEN_1668; // @[RAM_ST.scala 32:46]
  assign _GEN_1670 = 10'h2c1 == RADDR ? 10'h2c1 : _GEN_1669; // @[RAM_ST.scala 32:46]
  assign _GEN_1671 = 10'h2c2 == RADDR ? 10'h2c2 : _GEN_1670; // @[RAM_ST.scala 32:46]
  assign _GEN_1672 = 10'h2c3 == RADDR ? 10'h2c3 : _GEN_1671; // @[RAM_ST.scala 32:46]
  assign _GEN_1673 = 10'h2c4 == RADDR ? 10'h2c4 : _GEN_1672; // @[RAM_ST.scala 32:46]
  assign _GEN_1674 = 10'h2c5 == RADDR ? 10'h2c5 : _GEN_1673; // @[RAM_ST.scala 32:46]
  assign _GEN_1675 = 10'h2c6 == RADDR ? 10'h2c6 : _GEN_1674; // @[RAM_ST.scala 32:46]
  assign _GEN_1676 = 10'h2c7 == RADDR ? 10'h2c7 : _GEN_1675; // @[RAM_ST.scala 32:46]
  assign _GEN_1677 = 10'h2c8 == RADDR ? 10'h2c8 : _GEN_1676; // @[RAM_ST.scala 32:46]
  assign _GEN_1678 = 10'h2c9 == RADDR ? 10'h2c9 : _GEN_1677; // @[RAM_ST.scala 32:46]
  assign _GEN_1679 = 10'h2ca == RADDR ? 10'h2ca : _GEN_1678; // @[RAM_ST.scala 32:46]
  assign _GEN_1680 = 10'h2cb == RADDR ? 10'h2cb : _GEN_1679; // @[RAM_ST.scala 32:46]
  assign _GEN_1681 = 10'h2cc == RADDR ? 10'h2cc : _GEN_1680; // @[RAM_ST.scala 32:46]
  assign _GEN_1682 = 10'h2cd == RADDR ? 10'h2cd : _GEN_1681; // @[RAM_ST.scala 32:46]
  assign _GEN_1683 = 10'h2ce == RADDR ? 10'h2ce : _GEN_1682; // @[RAM_ST.scala 32:46]
  assign _GEN_1684 = 10'h2cf == RADDR ? 10'h2cf : _GEN_1683; // @[RAM_ST.scala 32:46]
  assign _GEN_1685 = 10'h2d0 == RADDR ? 10'h2d0 : _GEN_1684; // @[RAM_ST.scala 32:46]
  assign _GEN_1686 = 10'h2d1 == RADDR ? 10'h2d1 : _GEN_1685; // @[RAM_ST.scala 32:46]
  assign _GEN_1687 = 10'h2d2 == RADDR ? 10'h2d2 : _GEN_1686; // @[RAM_ST.scala 32:46]
  assign _GEN_1688 = 10'h2d3 == RADDR ? 10'h2d3 : _GEN_1687; // @[RAM_ST.scala 32:46]
  assign _GEN_1689 = 10'h2d4 == RADDR ? 10'h2d4 : _GEN_1688; // @[RAM_ST.scala 32:46]
  assign _GEN_1690 = 10'h2d5 == RADDR ? 10'h2d5 : _GEN_1689; // @[RAM_ST.scala 32:46]
  assign _GEN_1691 = 10'h2d6 == RADDR ? 10'h2d6 : _GEN_1690; // @[RAM_ST.scala 32:46]
  assign _GEN_1692 = 10'h2d7 == RADDR ? 10'h2d7 : _GEN_1691; // @[RAM_ST.scala 32:46]
  assign _GEN_1693 = 10'h2d8 == RADDR ? 10'h2d8 : _GEN_1692; // @[RAM_ST.scala 32:46]
  assign _GEN_1694 = 10'h2d9 == RADDR ? 10'h2d9 : _GEN_1693; // @[RAM_ST.scala 32:46]
  assign _GEN_1695 = 10'h2da == RADDR ? 10'h2da : _GEN_1694; // @[RAM_ST.scala 32:46]
  assign _GEN_1696 = 10'h2db == RADDR ? 10'h2db : _GEN_1695; // @[RAM_ST.scala 32:46]
  assign _GEN_1697 = 10'h2dc == RADDR ? 10'h2dc : _GEN_1696; // @[RAM_ST.scala 32:46]
  assign _GEN_1698 = 10'h2dd == RADDR ? 10'h2dd : _GEN_1697; // @[RAM_ST.scala 32:46]
  assign _GEN_1699 = 10'h2de == RADDR ? 10'h2de : _GEN_1698; // @[RAM_ST.scala 32:46]
  assign _GEN_1700 = 10'h2df == RADDR ? 10'h2df : _GEN_1699; // @[RAM_ST.scala 32:46]
  assign _GEN_1701 = 10'h2e0 == RADDR ? 10'h2e0 : _GEN_1700; // @[RAM_ST.scala 32:46]
  assign _GEN_1702 = 10'h2e1 == RADDR ? 10'h2e1 : _GEN_1701; // @[RAM_ST.scala 32:46]
  assign _GEN_1703 = 10'h2e2 == RADDR ? 10'h2e2 : _GEN_1702; // @[RAM_ST.scala 32:46]
  assign _GEN_1704 = 10'h2e3 == RADDR ? 10'h2e3 : _GEN_1703; // @[RAM_ST.scala 32:46]
  assign _GEN_1705 = 10'h2e4 == RADDR ? 10'h2e4 : _GEN_1704; // @[RAM_ST.scala 32:46]
  assign _GEN_1706 = 10'h2e5 == RADDR ? 10'h2e5 : _GEN_1705; // @[RAM_ST.scala 32:46]
  assign _GEN_1707 = 10'h2e6 == RADDR ? 10'h2e6 : _GEN_1706; // @[RAM_ST.scala 32:46]
  assign _GEN_1708 = 10'h2e7 == RADDR ? 10'h2e7 : _GEN_1707; // @[RAM_ST.scala 32:46]
  assign _GEN_1709 = 10'h2e8 == RADDR ? 10'h2e8 : _GEN_1708; // @[RAM_ST.scala 32:46]
  assign _GEN_1710 = 10'h2e9 == RADDR ? 10'h2e9 : _GEN_1709; // @[RAM_ST.scala 32:46]
  assign _GEN_1711 = 10'h2ea == RADDR ? 10'h2ea : _GEN_1710; // @[RAM_ST.scala 32:46]
  assign _GEN_1712 = 10'h2eb == RADDR ? 10'h2eb : _GEN_1711; // @[RAM_ST.scala 32:46]
  assign _GEN_1713 = 10'h2ec == RADDR ? 10'h2ec : _GEN_1712; // @[RAM_ST.scala 32:46]
  assign _GEN_1714 = 10'h2ed == RADDR ? 10'h2ed : _GEN_1713; // @[RAM_ST.scala 32:46]
  assign _GEN_1715 = 10'h2ee == RADDR ? 10'h2ee : _GEN_1714; // @[RAM_ST.scala 32:46]
  assign _GEN_1716 = 10'h2ef == RADDR ? 10'h2ef : _GEN_1715; // @[RAM_ST.scala 32:46]
  assign _GEN_1717 = 10'h2f0 == RADDR ? 10'h2f0 : _GEN_1716; // @[RAM_ST.scala 32:46]
  assign _GEN_1718 = 10'h2f1 == RADDR ? 10'h2f1 : _GEN_1717; // @[RAM_ST.scala 32:46]
  assign _GEN_1719 = 10'h2f2 == RADDR ? 10'h2f2 : _GEN_1718; // @[RAM_ST.scala 32:46]
  assign _GEN_1720 = 10'h2f3 == RADDR ? 10'h2f3 : _GEN_1719; // @[RAM_ST.scala 32:46]
  assign _GEN_1721 = 10'h2f4 == RADDR ? 10'h2f4 : _GEN_1720; // @[RAM_ST.scala 32:46]
  assign _GEN_1722 = 10'h2f5 == RADDR ? 10'h2f5 : _GEN_1721; // @[RAM_ST.scala 32:46]
  assign _GEN_1723 = 10'h2f6 == RADDR ? 10'h2f6 : _GEN_1722; // @[RAM_ST.scala 32:46]
  assign _GEN_1724 = 10'h2f7 == RADDR ? 10'h2f7 : _GEN_1723; // @[RAM_ST.scala 32:46]
  assign _GEN_1725 = 10'h2f8 == RADDR ? 10'h2f8 : _GEN_1724; // @[RAM_ST.scala 32:46]
  assign _GEN_1726 = 10'h2f9 == RADDR ? 10'h2f9 : _GEN_1725; // @[RAM_ST.scala 32:46]
  assign _GEN_1727 = 10'h2fa == RADDR ? 10'h2fa : _GEN_1726; // @[RAM_ST.scala 32:46]
  assign _GEN_1728 = 10'h2fb == RADDR ? 10'h2fb : _GEN_1727; // @[RAM_ST.scala 32:46]
  assign _GEN_1729 = 10'h2fc == RADDR ? 10'h2fc : _GEN_1728; // @[RAM_ST.scala 32:46]
  assign _GEN_1730 = 10'h2fd == RADDR ? 10'h2fd : _GEN_1729; // @[RAM_ST.scala 32:46]
  assign _GEN_1731 = 10'h2fe == RADDR ? 10'h2fe : _GEN_1730; // @[RAM_ST.scala 32:46]
  assign _GEN_1732 = 10'h2ff == RADDR ? 10'h2ff : _GEN_1731; // @[RAM_ST.scala 32:46]
  assign _GEN_1733 = 10'h300 == RADDR ? 10'h300 : _GEN_1732; // @[RAM_ST.scala 32:46]
  assign _GEN_1734 = 10'h301 == RADDR ? 10'h301 : _GEN_1733; // @[RAM_ST.scala 32:46]
  assign _GEN_1735 = 10'h302 == RADDR ? 10'h302 : _GEN_1734; // @[RAM_ST.scala 32:46]
  assign _GEN_1736 = 10'h303 == RADDR ? 10'h303 : _GEN_1735; // @[RAM_ST.scala 32:46]
  assign _GEN_1737 = 10'h304 == RADDR ? 10'h304 : _GEN_1736; // @[RAM_ST.scala 32:46]
  assign _GEN_1738 = 10'h305 == RADDR ? 10'h305 : _GEN_1737; // @[RAM_ST.scala 32:46]
  assign _GEN_1739 = 10'h306 == RADDR ? 10'h306 : _GEN_1738; // @[RAM_ST.scala 32:46]
  assign _GEN_1740 = 10'h307 == RADDR ? 10'h307 : _GEN_1739; // @[RAM_ST.scala 32:46]
  assign _GEN_1741 = 10'h308 == RADDR ? 10'h308 : _GEN_1740; // @[RAM_ST.scala 32:46]
  assign _GEN_1742 = 10'h309 == RADDR ? 10'h309 : _GEN_1741; // @[RAM_ST.scala 32:46]
  assign _GEN_1743 = 10'h30a == RADDR ? 10'h30a : _GEN_1742; // @[RAM_ST.scala 32:46]
  assign _GEN_1744 = 10'h30b == RADDR ? 10'h30b : _GEN_1743; // @[RAM_ST.scala 32:46]
  assign _GEN_1745 = 10'h30c == RADDR ? 10'h30c : _GEN_1744; // @[RAM_ST.scala 32:46]
  assign _GEN_1746 = 10'h30d == RADDR ? 10'h30d : _GEN_1745; // @[RAM_ST.scala 32:46]
  assign _GEN_1747 = 10'h30e == RADDR ? 10'h30e : _GEN_1746; // @[RAM_ST.scala 32:46]
  assign _GEN_1748 = 10'h30f == RADDR ? 10'h30f : _GEN_1747; // @[RAM_ST.scala 32:46]
  assign _GEN_1749 = 10'h310 == RADDR ? 10'h310 : _GEN_1748; // @[RAM_ST.scala 32:46]
  assign _GEN_1750 = 10'h311 == RADDR ? 10'h311 : _GEN_1749; // @[RAM_ST.scala 32:46]
  assign _GEN_1751 = 10'h312 == RADDR ? 10'h312 : _GEN_1750; // @[RAM_ST.scala 32:46]
  assign _GEN_1752 = 10'h313 == RADDR ? 10'h313 : _GEN_1751; // @[RAM_ST.scala 32:46]
  assign _GEN_1753 = 10'h314 == RADDR ? 10'h314 : _GEN_1752; // @[RAM_ST.scala 32:46]
  assign _GEN_1754 = 10'h315 == RADDR ? 10'h315 : _GEN_1753; // @[RAM_ST.scala 32:46]
  assign _GEN_1755 = 10'h316 == RADDR ? 10'h316 : _GEN_1754; // @[RAM_ST.scala 32:46]
  assign _GEN_1756 = 10'h317 == RADDR ? 10'h317 : _GEN_1755; // @[RAM_ST.scala 32:46]
  assign _GEN_1757 = 10'h318 == RADDR ? 10'h318 : _GEN_1756; // @[RAM_ST.scala 32:46]
  assign _GEN_1758 = 10'h319 == RADDR ? 10'h319 : _GEN_1757; // @[RAM_ST.scala 32:46]
  assign _GEN_1759 = 10'h31a == RADDR ? 10'h31a : _GEN_1758; // @[RAM_ST.scala 32:46]
  assign _GEN_1760 = 10'h31b == RADDR ? 10'h31b : _GEN_1759; // @[RAM_ST.scala 32:46]
  assign _GEN_1761 = 10'h31c == RADDR ? 10'h31c : _GEN_1760; // @[RAM_ST.scala 32:46]
  assign _GEN_1762 = 10'h31d == RADDR ? 10'h31d : _GEN_1761; // @[RAM_ST.scala 32:46]
  assign _GEN_1763 = 10'h31e == RADDR ? 10'h31e : _GEN_1762; // @[RAM_ST.scala 32:46]
  assign _GEN_1764 = 10'h31f == RADDR ? 10'h31f : _GEN_1763; // @[RAM_ST.scala 32:46]
  assign _GEN_1765 = 10'h320 == RADDR ? 10'h320 : _GEN_1764; // @[RAM_ST.scala 32:46]
  assign _GEN_1766 = 10'h321 == RADDR ? 10'h321 : _GEN_1765; // @[RAM_ST.scala 32:46]
  assign _GEN_1767 = 10'h322 == RADDR ? 10'h322 : _GEN_1766; // @[RAM_ST.scala 32:46]
  assign _GEN_1768 = 10'h323 == RADDR ? 10'h323 : _GEN_1767; // @[RAM_ST.scala 32:46]
  assign _GEN_1769 = 10'h324 == RADDR ? 10'h324 : _GEN_1768; // @[RAM_ST.scala 32:46]
  assign _GEN_1770 = 10'h325 == RADDR ? 10'h325 : _GEN_1769; // @[RAM_ST.scala 32:46]
  assign _GEN_1771 = 10'h326 == RADDR ? 10'h326 : _GEN_1770; // @[RAM_ST.scala 32:46]
  assign _GEN_1772 = 10'h327 == RADDR ? 10'h327 : _GEN_1771; // @[RAM_ST.scala 32:46]
  assign _GEN_1773 = 10'h328 == RADDR ? 10'h328 : _GEN_1772; // @[RAM_ST.scala 32:46]
  assign _GEN_1774 = 10'h329 == RADDR ? 10'h329 : _GEN_1773; // @[RAM_ST.scala 32:46]
  assign _GEN_1775 = 10'h32a == RADDR ? 10'h32a : _GEN_1774; // @[RAM_ST.scala 32:46]
  assign _GEN_1776 = 10'h32b == RADDR ? 10'h32b : _GEN_1775; // @[RAM_ST.scala 32:46]
  assign _GEN_1777 = 10'h32c == RADDR ? 10'h32c : _GEN_1776; // @[RAM_ST.scala 32:46]
  assign _GEN_1778 = 10'h32d == RADDR ? 10'h32d : _GEN_1777; // @[RAM_ST.scala 32:46]
  assign _GEN_1779 = 10'h32e == RADDR ? 10'h32e : _GEN_1778; // @[RAM_ST.scala 32:46]
  assign _GEN_1780 = 10'h32f == RADDR ? 10'h32f : _GEN_1779; // @[RAM_ST.scala 32:46]
  assign _GEN_1781 = 10'h330 == RADDR ? 10'h330 : _GEN_1780; // @[RAM_ST.scala 32:46]
  assign _GEN_1782 = 10'h331 == RADDR ? 10'h331 : _GEN_1781; // @[RAM_ST.scala 32:46]
  assign _GEN_1783 = 10'h332 == RADDR ? 10'h332 : _GEN_1782; // @[RAM_ST.scala 32:46]
  assign _GEN_1784 = 10'h333 == RADDR ? 10'h333 : _GEN_1783; // @[RAM_ST.scala 32:46]
  assign _GEN_1785 = 10'h334 == RADDR ? 10'h334 : _GEN_1784; // @[RAM_ST.scala 32:46]
  assign _GEN_1786 = 10'h335 == RADDR ? 10'h335 : _GEN_1785; // @[RAM_ST.scala 32:46]
  assign _GEN_1787 = 10'h336 == RADDR ? 10'h336 : _GEN_1786; // @[RAM_ST.scala 32:46]
  assign _GEN_1788 = 10'h337 == RADDR ? 10'h337 : _GEN_1787; // @[RAM_ST.scala 32:46]
  assign _GEN_1789 = 10'h338 == RADDR ? 10'h338 : _GEN_1788; // @[RAM_ST.scala 32:46]
  assign _GEN_1790 = 10'h339 == RADDR ? 10'h339 : _GEN_1789; // @[RAM_ST.scala 32:46]
  assign _GEN_1791 = 10'h33a == RADDR ? 10'h33a : _GEN_1790; // @[RAM_ST.scala 32:46]
  assign _GEN_1792 = 10'h33b == RADDR ? 10'h33b : _GEN_1791; // @[RAM_ST.scala 32:46]
  assign _GEN_1793 = 10'h33c == RADDR ? 10'h33c : _GEN_1792; // @[RAM_ST.scala 32:46]
  assign _GEN_1794 = 10'h33d == RADDR ? 10'h33d : _GEN_1793; // @[RAM_ST.scala 32:46]
  assign _GEN_1795 = 10'h33e == RADDR ? 10'h33e : _GEN_1794; // @[RAM_ST.scala 32:46]
  assign _GEN_1796 = 10'h33f == RADDR ? 10'h33f : _GEN_1795; // @[RAM_ST.scala 32:46]
  assign _GEN_1797 = 10'h340 == RADDR ? 10'h340 : _GEN_1796; // @[RAM_ST.scala 32:46]
  assign _GEN_1798 = 10'h341 == RADDR ? 10'h341 : _GEN_1797; // @[RAM_ST.scala 32:46]
  assign _GEN_1799 = 10'h342 == RADDR ? 10'h342 : _GEN_1798; // @[RAM_ST.scala 32:46]
  assign _GEN_1800 = 10'h343 == RADDR ? 10'h343 : _GEN_1799; // @[RAM_ST.scala 32:46]
  assign _GEN_1801 = 10'h344 == RADDR ? 10'h344 : _GEN_1800; // @[RAM_ST.scala 32:46]
  assign _GEN_1802 = 10'h345 == RADDR ? 10'h345 : _GEN_1801; // @[RAM_ST.scala 32:46]
  assign _GEN_1803 = 10'h346 == RADDR ? 10'h346 : _GEN_1802; // @[RAM_ST.scala 32:46]
  assign _GEN_1804 = 10'h347 == RADDR ? 10'h347 : _GEN_1803; // @[RAM_ST.scala 32:46]
  assign _GEN_1805 = 10'h348 == RADDR ? 10'h348 : _GEN_1804; // @[RAM_ST.scala 32:46]
  assign _GEN_1806 = 10'h349 == RADDR ? 10'h349 : _GEN_1805; // @[RAM_ST.scala 32:46]
  assign _GEN_1807 = 10'h34a == RADDR ? 10'h34a : _GEN_1806; // @[RAM_ST.scala 32:46]
  assign _GEN_1808 = 10'h34b == RADDR ? 10'h34b : _GEN_1807; // @[RAM_ST.scala 32:46]
  assign _GEN_1809 = 10'h34c == RADDR ? 10'h34c : _GEN_1808; // @[RAM_ST.scala 32:46]
  assign _GEN_1810 = 10'h34d == RADDR ? 10'h34d : _GEN_1809; // @[RAM_ST.scala 32:46]
  assign _GEN_1811 = 10'h34e == RADDR ? 10'h34e : _GEN_1810; // @[RAM_ST.scala 32:46]
  assign _GEN_1812 = 10'h34f == RADDR ? 10'h34f : _GEN_1811; // @[RAM_ST.scala 32:46]
  assign _GEN_1813 = 10'h350 == RADDR ? 10'h350 : _GEN_1812; // @[RAM_ST.scala 32:46]
  assign _GEN_1814 = 10'h351 == RADDR ? 10'h351 : _GEN_1813; // @[RAM_ST.scala 32:46]
  assign _GEN_1815 = 10'h352 == RADDR ? 10'h352 : _GEN_1814; // @[RAM_ST.scala 32:46]
  assign _GEN_1816 = 10'h353 == RADDR ? 10'h353 : _GEN_1815; // @[RAM_ST.scala 32:46]
  assign _GEN_1817 = 10'h354 == RADDR ? 10'h354 : _GEN_1816; // @[RAM_ST.scala 32:46]
  assign _GEN_1818 = 10'h355 == RADDR ? 10'h355 : _GEN_1817; // @[RAM_ST.scala 32:46]
  assign _GEN_1819 = 10'h356 == RADDR ? 10'h356 : _GEN_1818; // @[RAM_ST.scala 32:46]
  assign _GEN_1820 = 10'h357 == RADDR ? 10'h357 : _GEN_1819; // @[RAM_ST.scala 32:46]
  assign _GEN_1821 = 10'h358 == RADDR ? 10'h358 : _GEN_1820; // @[RAM_ST.scala 32:46]
  assign _GEN_1822 = 10'h359 == RADDR ? 10'h359 : _GEN_1821; // @[RAM_ST.scala 32:46]
  assign _GEN_1823 = 10'h35a == RADDR ? 10'h35a : _GEN_1822; // @[RAM_ST.scala 32:46]
  assign _GEN_1824 = 10'h35b == RADDR ? 10'h35b : _GEN_1823; // @[RAM_ST.scala 32:46]
  assign _GEN_1825 = 10'h35c == RADDR ? 10'h35c : _GEN_1824; // @[RAM_ST.scala 32:46]
  assign _GEN_1826 = 10'h35d == RADDR ? 10'h35d : _GEN_1825; // @[RAM_ST.scala 32:46]
  assign _GEN_1827 = 10'h35e == RADDR ? 10'h35e : _GEN_1826; // @[RAM_ST.scala 32:46]
  assign _GEN_1828 = 10'h35f == RADDR ? 10'h35f : _GEN_1827; // @[RAM_ST.scala 32:46]
  assign _GEN_1829 = 10'h360 == RADDR ? 10'h360 : _GEN_1828; // @[RAM_ST.scala 32:46]
  assign _GEN_1830 = 10'h361 == RADDR ? 10'h361 : _GEN_1829; // @[RAM_ST.scala 32:46]
  assign _GEN_1831 = 10'h362 == RADDR ? 10'h362 : _GEN_1830; // @[RAM_ST.scala 32:46]
  assign _GEN_1832 = 10'h363 == RADDR ? 10'h363 : _GEN_1831; // @[RAM_ST.scala 32:46]
  assign _GEN_1833 = 10'h364 == RADDR ? 10'h364 : _GEN_1832; // @[RAM_ST.scala 32:46]
  assign _GEN_1834 = 10'h365 == RADDR ? 10'h365 : _GEN_1833; // @[RAM_ST.scala 32:46]
  assign _GEN_1835 = 10'h366 == RADDR ? 10'h366 : _GEN_1834; // @[RAM_ST.scala 32:46]
  assign _GEN_1836 = 10'h367 == RADDR ? 10'h367 : _GEN_1835; // @[RAM_ST.scala 32:46]
  assign _GEN_1837 = 10'h368 == RADDR ? 10'h368 : _GEN_1836; // @[RAM_ST.scala 32:46]
  assign _GEN_1838 = 10'h369 == RADDR ? 10'h369 : _GEN_1837; // @[RAM_ST.scala 32:46]
  assign _GEN_1839 = 10'h36a == RADDR ? 10'h36a : _GEN_1838; // @[RAM_ST.scala 32:46]
  assign _GEN_1840 = 10'h36b == RADDR ? 10'h36b : _GEN_1839; // @[RAM_ST.scala 32:46]
  assign _GEN_1841 = 10'h36c == RADDR ? 10'h36c : _GEN_1840; // @[RAM_ST.scala 32:46]
  assign _GEN_1842 = 10'h36d == RADDR ? 10'h36d : _GEN_1841; // @[RAM_ST.scala 32:46]
  assign _GEN_1843 = 10'h36e == RADDR ? 10'h36e : _GEN_1842; // @[RAM_ST.scala 32:46]
  assign _GEN_1844 = 10'h36f == RADDR ? 10'h36f : _GEN_1843; // @[RAM_ST.scala 32:46]
  assign _GEN_1845 = 10'h370 == RADDR ? 10'h370 : _GEN_1844; // @[RAM_ST.scala 32:46]
  assign _GEN_1846 = 10'h371 == RADDR ? 10'h371 : _GEN_1845; // @[RAM_ST.scala 32:46]
  assign _GEN_1847 = 10'h372 == RADDR ? 10'h372 : _GEN_1846; // @[RAM_ST.scala 32:46]
  assign _GEN_1848 = 10'h373 == RADDR ? 10'h373 : _GEN_1847; // @[RAM_ST.scala 32:46]
  assign _GEN_1849 = 10'h374 == RADDR ? 10'h374 : _GEN_1848; // @[RAM_ST.scala 32:46]
  assign _GEN_1850 = 10'h375 == RADDR ? 10'h375 : _GEN_1849; // @[RAM_ST.scala 32:46]
  assign _GEN_1851 = 10'h376 == RADDR ? 10'h376 : _GEN_1850; // @[RAM_ST.scala 32:46]
  assign _GEN_1852 = 10'h377 == RADDR ? 10'h377 : _GEN_1851; // @[RAM_ST.scala 32:46]
  assign _GEN_1853 = 10'h378 == RADDR ? 10'h378 : _GEN_1852; // @[RAM_ST.scala 32:46]
  assign _GEN_1854 = 10'h379 == RADDR ? 10'h379 : _GEN_1853; // @[RAM_ST.scala 32:46]
  assign _GEN_1855 = 10'h37a == RADDR ? 10'h37a : _GEN_1854; // @[RAM_ST.scala 32:46]
  assign _GEN_1856 = 10'h37b == RADDR ? 10'h37b : _GEN_1855; // @[RAM_ST.scala 32:46]
  assign _GEN_1857 = 10'h37c == RADDR ? 10'h37c : _GEN_1856; // @[RAM_ST.scala 32:46]
  assign _GEN_1858 = 10'h37d == RADDR ? 10'h37d : _GEN_1857; // @[RAM_ST.scala 32:46]
  assign _GEN_1859 = 10'h37e == RADDR ? 10'h37e : _GEN_1858; // @[RAM_ST.scala 32:46]
  assign _GEN_1860 = 10'h37f == RADDR ? 10'h37f : _GEN_1859; // @[RAM_ST.scala 32:46]
  assign _GEN_1861 = 10'h380 == RADDR ? 10'h380 : _GEN_1860; // @[RAM_ST.scala 32:46]
  assign _GEN_1862 = 10'h381 == RADDR ? 10'h381 : _GEN_1861; // @[RAM_ST.scala 32:46]
  assign _GEN_1863 = 10'h382 == RADDR ? 10'h382 : _GEN_1862; // @[RAM_ST.scala 32:46]
  assign _GEN_1864 = 10'h383 == RADDR ? 10'h383 : _GEN_1863; // @[RAM_ST.scala 32:46]
  assign _GEN_1865 = 10'h384 == RADDR ? 10'h384 : _GEN_1864; // @[RAM_ST.scala 32:46]
  assign _GEN_1866 = 10'h385 == RADDR ? 10'h385 : _GEN_1865; // @[RAM_ST.scala 32:46]
  assign _GEN_1867 = 10'h386 == RADDR ? 10'h386 : _GEN_1866; // @[RAM_ST.scala 32:46]
  assign _GEN_1868 = 10'h387 == RADDR ? 10'h387 : _GEN_1867; // @[RAM_ST.scala 32:46]
  assign _GEN_1869 = 10'h388 == RADDR ? 10'h388 : _GEN_1868; // @[RAM_ST.scala 32:46]
  assign _GEN_1870 = 10'h389 == RADDR ? 10'h389 : _GEN_1869; // @[RAM_ST.scala 32:46]
  assign _GEN_1871 = 10'h38a == RADDR ? 10'h38a : _GEN_1870; // @[RAM_ST.scala 32:46]
  assign _GEN_1872 = 10'h38b == RADDR ? 10'h38b : _GEN_1871; // @[RAM_ST.scala 32:46]
  assign _GEN_1873 = 10'h38c == RADDR ? 10'h38c : _GEN_1872; // @[RAM_ST.scala 32:46]
  assign _GEN_1874 = 10'h38d == RADDR ? 10'h38d : _GEN_1873; // @[RAM_ST.scala 32:46]
  assign _GEN_1875 = 10'h38e == RADDR ? 10'h38e : _GEN_1874; // @[RAM_ST.scala 32:46]
  assign _GEN_1876 = 10'h38f == RADDR ? 10'h38f : _GEN_1875; // @[RAM_ST.scala 32:46]
  assign _GEN_1877 = 10'h390 == RADDR ? 10'h390 : _GEN_1876; // @[RAM_ST.scala 32:46]
  assign _GEN_1878 = 10'h391 == RADDR ? 10'h391 : _GEN_1877; // @[RAM_ST.scala 32:46]
  assign _GEN_1879 = 10'h392 == RADDR ? 10'h392 : _GEN_1878; // @[RAM_ST.scala 32:46]
  assign _GEN_1880 = 10'h393 == RADDR ? 10'h393 : _GEN_1879; // @[RAM_ST.scala 32:46]
  assign _GEN_1881 = 10'h394 == RADDR ? 10'h394 : _GEN_1880; // @[RAM_ST.scala 32:46]
  assign _GEN_1882 = 10'h395 == RADDR ? 10'h395 : _GEN_1881; // @[RAM_ST.scala 32:46]
  assign _GEN_1883 = 10'h396 == RADDR ? 10'h396 : _GEN_1882; // @[RAM_ST.scala 32:46]
  assign _GEN_1884 = 10'h397 == RADDR ? 10'h397 : _GEN_1883; // @[RAM_ST.scala 32:46]
  assign _GEN_1885 = 10'h398 == RADDR ? 10'h398 : _GEN_1884; // @[RAM_ST.scala 32:46]
  assign _GEN_1886 = 10'h399 == RADDR ? 10'h399 : _GEN_1885; // @[RAM_ST.scala 32:46]
  assign _GEN_1887 = 10'h39a == RADDR ? 10'h39a : _GEN_1886; // @[RAM_ST.scala 32:46]
  assign _GEN_1888 = 10'h39b == RADDR ? 10'h39b : _GEN_1887; // @[RAM_ST.scala 32:46]
  assign _GEN_1889 = 10'h39c == RADDR ? 10'h39c : _GEN_1888; // @[RAM_ST.scala 32:46]
  assign _GEN_1890 = 10'h39d == RADDR ? 10'h39d : _GEN_1889; // @[RAM_ST.scala 32:46]
  assign _GEN_1891 = 10'h39e == RADDR ? 10'h39e : _GEN_1890; // @[RAM_ST.scala 32:46]
  assign _GEN_1892 = 10'h39f == RADDR ? 10'h39f : _GEN_1891; // @[RAM_ST.scala 32:46]
  assign _GEN_1893 = 10'h3a0 == RADDR ? 10'h3a0 : _GEN_1892; // @[RAM_ST.scala 32:46]
  assign _GEN_1894 = 10'h3a1 == RADDR ? 10'h3a1 : _GEN_1893; // @[RAM_ST.scala 32:46]
  assign _GEN_1895 = 10'h3a2 == RADDR ? 10'h3a2 : _GEN_1894; // @[RAM_ST.scala 32:46]
  assign _GEN_1896 = 10'h3a3 == RADDR ? 10'h3a3 : _GEN_1895; // @[RAM_ST.scala 32:46]
  assign _GEN_1897 = 10'h3a4 == RADDR ? 10'h3a4 : _GEN_1896; // @[RAM_ST.scala 32:46]
  assign _GEN_1898 = 10'h3a5 == RADDR ? 10'h3a5 : _GEN_1897; // @[RAM_ST.scala 32:46]
  assign _GEN_1899 = 10'h3a6 == RADDR ? 10'h3a6 : _GEN_1898; // @[RAM_ST.scala 32:46]
  assign _GEN_1900 = 10'h3a7 == RADDR ? 10'h3a7 : _GEN_1899; // @[RAM_ST.scala 32:46]
  assign _GEN_1901 = 10'h3a8 == RADDR ? 10'h3a8 : _GEN_1900; // @[RAM_ST.scala 32:46]
  assign _GEN_1902 = 10'h3a9 == RADDR ? 10'h3a9 : _GEN_1901; // @[RAM_ST.scala 32:46]
  assign _GEN_1903 = 10'h3aa == RADDR ? 10'h3aa : _GEN_1902; // @[RAM_ST.scala 32:46]
  assign _GEN_1904 = 10'h3ab == RADDR ? 10'h3ab : _GEN_1903; // @[RAM_ST.scala 32:46]
  assign _GEN_1905 = 10'h3ac == RADDR ? 10'h3ac : _GEN_1904; // @[RAM_ST.scala 32:46]
  assign _GEN_1906 = 10'h3ad == RADDR ? 10'h3ad : _GEN_1905; // @[RAM_ST.scala 32:46]
  assign _GEN_1907 = 10'h3ae == RADDR ? 10'h3ae : _GEN_1906; // @[RAM_ST.scala 32:46]
  assign _GEN_1908 = 10'h3af == RADDR ? 10'h3af : _GEN_1907; // @[RAM_ST.scala 32:46]
  assign _GEN_1909 = 10'h3b0 == RADDR ? 10'h3b0 : _GEN_1908; // @[RAM_ST.scala 32:46]
  assign _GEN_1910 = 10'h3b1 == RADDR ? 10'h3b1 : _GEN_1909; // @[RAM_ST.scala 32:46]
  assign _GEN_1911 = 10'h3b2 == RADDR ? 10'h3b2 : _GEN_1910; // @[RAM_ST.scala 32:46]
  assign _GEN_1912 = 10'h3b3 == RADDR ? 10'h3b3 : _GEN_1911; // @[RAM_ST.scala 32:46]
  assign _GEN_1913 = 10'h3b4 == RADDR ? 10'h3b4 : _GEN_1912; // @[RAM_ST.scala 32:46]
  assign _GEN_1914 = 10'h3b5 == RADDR ? 10'h3b5 : _GEN_1913; // @[RAM_ST.scala 32:46]
  assign _GEN_1915 = 10'h3b6 == RADDR ? 10'h3b6 : _GEN_1914; // @[RAM_ST.scala 32:46]
  assign _GEN_1916 = 10'h3b7 == RADDR ? 10'h3b7 : _GEN_1915; // @[RAM_ST.scala 32:46]
  assign _GEN_1917 = 10'h3b8 == RADDR ? 10'h3b8 : _GEN_1916; // @[RAM_ST.scala 32:46]
  assign _GEN_1918 = 10'h3b9 == RADDR ? 10'h3b9 : _GEN_1917; // @[RAM_ST.scala 32:46]
  assign _GEN_1919 = 10'h3ba == RADDR ? 10'h3ba : _GEN_1918; // @[RAM_ST.scala 32:46]
  assign _GEN_1920 = 10'h3bb == RADDR ? 10'h3bb : _GEN_1919; // @[RAM_ST.scala 32:46]
  assign _GEN_1921 = 10'h3bc == RADDR ? 10'h3bc : _GEN_1920; // @[RAM_ST.scala 32:46]
  assign _GEN_1922 = 10'h3bd == RADDR ? 10'h3bd : _GEN_1921; // @[RAM_ST.scala 32:46]
  assign _GEN_1923 = 10'h3be == RADDR ? 10'h3be : _GEN_1922; // @[RAM_ST.scala 32:46]
  assign _GEN_1924 = 10'h3bf == RADDR ? 10'h3bf : _GEN_1923; // @[RAM_ST.scala 32:46]
  assign _T_4 = {{1'd0}, _GEN_1924}; // @[RAM_ST.scala 32:46]
  assign _T_11 = ram__T_9_data;
  assign RDATA_0 = _T_11[7:0]; // @[RAM_ST.scala 32:9]
  assign RDATA_1 = _T_11[15:8]; // @[RAM_ST.scala 32:9]
  assign write_elem_counter_CE = WE; // @[RAM_ST.scala 23:25]
  assign read_elem_counter_CE = RE; // @[RAM_ST.scala 24:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 960; initvar = initvar+1)
    ram[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram__T_9_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ram__T_9_addr_pipe_0 = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram__T_3_en & ram__T_3_mask) begin
      ram[ram__T_3_addr] <= ram__T_3_data; // @[RAM_ST.scala 29:24]
    end
    ram__T_9_en_pipe_0 <= read_elem_counter_valid;
    if (read_elem_counter_valid) begin
      ram__T_9_addr_pipe_0 <= _T_4[9:0];
    end
  end
endmodule
module ShiftT(
  input        clock,
  input        reset,
  input        valid_up,
  input  [7:0] I_0,
  input  [7:0] I_1,
  output [7:0] O_0,
  output [7:0] O_1
);
  wire  RAM_ST_clock; // @[ShiftT.scala 39:29]
  wire  RAM_ST_RE; // @[ShiftT.scala 39:29]
  wire [9:0] RAM_ST_RADDR; // @[ShiftT.scala 39:29]
  wire [7:0] RAM_ST_RDATA_0; // @[ShiftT.scala 39:29]
  wire [7:0] RAM_ST_RDATA_1; // @[ShiftT.scala 39:29]
  wire  RAM_ST_WE; // @[ShiftT.scala 39:29]
  wire [9:0] RAM_ST_WADDR; // @[ShiftT.scala 39:29]
  wire [7:0] RAM_ST_WDATA_0; // @[ShiftT.scala 39:29]
  wire [7:0] RAM_ST_WDATA_1; // @[ShiftT.scala 39:29]
  wire  NestedCounters_CE; // @[ShiftT.scala 41:31]
  wire  NestedCounters_valid; // @[ShiftT.scala 41:31]
  reg [9:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[Counter.scala 37:24]
  wire [9:0] _T_3; // @[Counter.scala 38:22]
  RAM_ST RAM_ST ( // @[ShiftT.scala 39:29]
    .clock(RAM_ST_clock),
    .RE(RAM_ST_RE),
    .RADDR(RAM_ST_RADDR),
    .RDATA_0(RAM_ST_RDATA_0),
    .RDATA_1(RAM_ST_RDATA_1),
    .WE(RAM_ST_WE),
    .WADDR(RAM_ST_WADDR),
    .WDATA_0(RAM_ST_WDATA_0),
    .WDATA_1(RAM_ST_WDATA_1)
  );
  NestedCounters_1 NestedCounters ( // @[ShiftT.scala 41:31]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign _T_1 = value == 10'h3bf; // @[Counter.scala 37:24]
  assign _T_3 = value + 10'h1; // @[Counter.scala 38:22]
  assign O_0 = RAM_ST_RDATA_0; // @[ShiftT.scala 51:7]
  assign O_1 = RAM_ST_RDATA_1; // @[ShiftT.scala 51:7]
  assign RAM_ST_clock = clock;
  assign RAM_ST_RE = valid_up; // @[ShiftT.scala 49:20]
  assign RAM_ST_RADDR = _T_1 ? 10'h0 : _T_3; // @[ShiftT.scala 46:76 ShiftT.scala 47:38]
  assign RAM_ST_WE = valid_up; // @[ShiftT.scala 48:20]
  assign RAM_ST_WADDR = value; // @[ShiftT.scala 45:23]
  assign RAM_ST_WDATA_0 = I_0; // @[ShiftT.scala 50:23]
  assign RAM_ST_WDATA_1 = I_1; // @[ShiftT.scala 50:23]
  assign NestedCounters_CE = valid_up; // @[ShiftT.scala 42:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[9:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 10'h0;
    end else if (valid_up) begin
      if (_T_1) begin
        value <= 10'h0;
      end else begin
        value <= _T_3;
      end
    end
  end
endmodule
module ShiftTS(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  output [7:0] O_0,
  output [7:0] O_1
);
  wire  ShiftT_clock; // @[ShiftTS.scala 32:26]
  wire  ShiftT_reset; // @[ShiftTS.scala 32:26]
  wire  ShiftT_valid_up; // @[ShiftTS.scala 32:26]
  wire [7:0] ShiftT_I_0; // @[ShiftTS.scala 32:26]
  wire [7:0] ShiftT_I_1; // @[ShiftTS.scala 32:26]
  wire [7:0] ShiftT_O_0; // @[ShiftTS.scala 32:26]
  wire [7:0] ShiftT_O_1; // @[ShiftTS.scala 32:26]
  ShiftT ShiftT ( // @[ShiftTS.scala 32:26]
    .clock(ShiftT_clock),
    .reset(ShiftT_reset),
    .valid_up(ShiftT_valid_up),
    .I_0(ShiftT_I_0),
    .I_1(ShiftT_I_1),
    .O_0(ShiftT_O_0),
    .O_1(ShiftT_O_1)
  );
  assign valid_down = valid_up; // @[ShiftTS.scala 58:14]
  assign O_0 = ShiftT_O_0; // @[ShiftTS.scala 51:36]
  assign O_1 = ShiftT_O_1; // @[ShiftTS.scala 51:36]
  assign ShiftT_clock = clock;
  assign ShiftT_reset = reset;
  assign ShiftT_valid_up = valid_up; // @[ShiftTS.scala 53:29]
  assign ShiftT_I_0 = I_0; // @[ShiftTS.scala 50:25]
  assign ShiftT_I_1 = I_1; // @[ShiftTS.scala 50:25]
endmodule
module ShiftT_2(
  input        clock,
  input  [7:0] I_0,
  output [7:0] O_0
);
  reg [7:0] _T_0; // @[ShiftT.scala 24:82]
  reg [31:0] _RAND_0;
  assign O_0 = _T_0; // @[ShiftT.scala 24:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0 <= I_0;
  end
endmodule
module ShiftTS_2(
  input        clock,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  output [7:0] O_0,
  output [7:0] O_1
);
  wire  ShiftT_clock; // @[ShiftTS.scala 32:26]
  wire [7:0] ShiftT_I_0; // @[ShiftTS.scala 32:26]
  wire [7:0] ShiftT_O_0; // @[ShiftTS.scala 32:26]
  ShiftT_2 ShiftT ( // @[ShiftTS.scala 32:26]
    .clock(ShiftT_clock),
    .I_0(ShiftT_I_0),
    .O_0(ShiftT_O_0)
  );
  assign valid_down = valid_up; // @[ShiftTS.scala 58:14]
  assign O_0 = ShiftT_O_0; // @[ShiftTS.scala 51:36]
  assign O_1 = I_0; // @[ShiftTS.scala 40:36]
  assign ShiftT_clock = clock;
  assign ShiftT_I_0 = I_1; // @[ShiftTS.scala 50:25]
endmodule
module SSeqTupleCreator(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  input  [7:0] I1,
  output [7:0] O_0,
  output [7:0] O_1
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0 = I0; // @[Tuple.scala 12:32]
  assign O_1 = I1; // @[Tuple.scala 13:32]
endmodule
module Map2S(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_1_0,
  output [7:0] O_1_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1; // @[Map2S.scala 10:86]
  SSeqTupleCreator fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1)
  );
  SSeqTupleCreator other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_1_0 = other_ops_0_O_0; // @[Map2S.scala 24:12]
  assign O_1_1 = other_ops_0_O_1; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
endmodule
module Map2T(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_1_0,
  output [7:0] O_1_1
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_1; // @[Map2T.scala 8:20]
  Map2S op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0(op_I0_0),
    .I0_1(op_I0_1),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0 = op_O_0_0; // @[Map2T.scala 17:7]
  assign O_0_1 = op_O_0_1; // @[Map2T.scala 17:7]
  assign O_1_0 = op_O_1_0; // @[Map2T.scala 17:7]
  assign O_1_1 = op_O_1_1; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0 = I0_0; // @[Map2T.scala 15:11]
  assign op_I0_1 = I0_1; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleAppender(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I1,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0 = I0_0; // @[Tuple.scala 24:34]
  assign O_1 = I0_1; // @[Tuple.scala 24:34]
  assign O_2 = I1; // @[Tuple.scala 26:32]
endmodule
module Map2S_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2; // @[Map2S.scala 10:86]
  SSeqTupleAppender fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  SSeqTupleAppender other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I1(other_ops_0_I1),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_0_2 = fst_op_O_2; // @[Map2S.scala 19:8]
  assign O_1_0 = other_ops_0_O_0; // @[Map2S.scala 24:12]
  assign O_1_1 = other_ops_0_O_1; // @[Map2S.scala 24:12]
  assign O_1_2 = other_ops_0_O_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
endmodule
module Map2T_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_2; // @[Map2T.scala 8:20]
  Map2S_1 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0(op_I0_0_0),
    .I0_0_1(op_I0_0_1),
    .I0_1_0(op_I0_1_0),
    .I0_1_1(op_I0_1_1),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_0_2(op_O_0_2),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_1_2(op_O_1_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0 = op_O_0_0; // @[Map2T.scala 17:7]
  assign O_0_1 = op_O_0_1; // @[Map2T.scala 17:7]
  assign O_0_2 = op_O_0_2; // @[Map2T.scala 17:7]
  assign O_1_0 = op_O_1_0; // @[Map2T.scala 17:7]
  assign O_1_1 = op_O_1_1; // @[Map2T.scala 17:7]
  assign O_1_2 = op_O_1_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0 = I0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1 = I0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0 = I0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1 = I0_1_1; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
endmodule
module PartitionS(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0 = I_0_0; // @[Partition.scala 15:39]
  assign O_0_0_1 = I_0_1; // @[Partition.scala 15:39]
  assign O_0_0_2 = I_0_2; // @[Partition.scala 15:39]
  assign O_1_0_0 = I_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1 = I_1_1; // @[Partition.scala 15:39]
  assign O_1_0_2 = I_1_2; // @[Partition.scala 15:39]
endmodule
module MapT(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_2; // @[MapT.scala 8:20]
  PartitionS op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0(op_I_0_0),
    .I_0_1(op_I_0_1),
    .I_0_2(op_I_0_2),
    .I_1_0(op_I_1_0),
    .I_1_1(op_I_1_1),
    .I_1_2(op_I_1_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_2 = op_O_0_0_2; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_0_2 = op_O_1_0_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0 = I_0_0; // @[MapT.scala 14:10]
  assign op_I_0_1 = I_0_1; // @[MapT.scala 14:10]
  assign op_I_0_2 = I_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0 = I_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1 = I_1_1; // @[MapT.scala 14:10]
  assign op_I_1_2 = I_1_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleToSSeq(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0 = I_0; // @[Tuple.scala 41:5]
  assign O_1 = I_1; // @[Tuple.scala 41:5]
  assign O_2 = I_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0(op_inst_I_0),
    .I_1(op_inst_I_1),
    .I_2(op_inst_I_2),
    .O_0(op_inst_O_0),
    .O_1(op_inst_O_1),
    .O_2(op_inst_O_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0 = op_inst_O_0; // @[Remove1S.scala 14:5]
  assign O_1 = op_inst_O_1; // @[Remove1S.scala 14:5]
  assign O_2 = op_inst_O_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0 = I_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1 = I_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2 = I_0_2; // @[Remove1S.scala 13:13]
endmodule
module MapS(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2; // @[MapS.scala 10:86]
  Remove1S fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  Remove1S other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_1_2 = other_ops_0_O_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
endmodule
module MapT_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_2; // @[MapT.scala 8:20]
  MapS op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_0_2(op_O_0_2),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_1_2(op_O_1_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0 = op_O_0_0; // @[MapT.scala 15:7]
  assign O_0_1 = op_O_0_1; // @[MapT.scala 15:7]
  assign O_0_2 = op_O_0_2; // @[MapT.scala 15:7]
  assign O_1_0 = op_O_1_0; // @[MapT.scala 15:7]
  assign O_1_1 = op_O_1_1; // @[MapT.scala 15:7]
  assign O_1_2 = op_O_1_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleCreator_2(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I0_2,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0_0 = I0_0; // @[Tuple.scala 12:32]
  assign O_0_1 = I0_1; // @[Tuple.scala 12:32]
  assign O_0_2 = I0_2; // @[Tuple.scala 12:32]
  assign O_1_0 = I1_0; // @[Tuple.scala 13:32]
  assign O_1_1 = I1_1; // @[Tuple.scala 13:32]
  assign O_1_2 = I1_2; // @[Tuple.scala 13:32]
endmodule
module Map2S_4(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_0_2,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_1_2,
  input  [7:0] I1_0_0,
  input  [7:0] I1_0_1,
  input  [7:0] I1_0_2,
  input  [7:0] I1_1_0,
  input  [7:0] I1_1_1,
  input  [7:0] I1_1_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_2; // @[Map2S.scala 10:86]
  SSeqTupleCreator_2 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I0_2(other_ops_0_I0_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[Map2S.scala 24:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[Map2S.scala 24:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[Map2S.scala 24:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2 = I0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = I1_1_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = I1_1_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = I1_1_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_4(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_0_2,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_1_2,
  input  [7:0] I1_0_0,
  input  [7:0] I1_0_1,
  input  [7:0] I1_0_2,
  input  [7:0] I1_1_0,
  input  [7:0] I1_1_1,
  input  [7:0] I1_1_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_1_2; // @[Map2T.scala 8:20]
  Map2S_4 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0(op_I0_0_0),
    .I0_0_1(op_I0_0_1),
    .I0_0_2(op_I0_0_2),
    .I0_1_0(op_I0_1_0),
    .I0_1_1(op_I0_1_1),
    .I0_1_2(op_I0_1_2),
    .I1_0_0(op_I1_0_0),
    .I1_0_1(op_I1_0_1),
    .I1_0_2(op_I1_0_2),
    .I1_1_0(op_I1_1_0),
    .I1_1_1(op_I1_1_1),
    .I1_1_2(op_I1_1_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0 = op_O_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_1 = op_O_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_2 = op_O_0_0_2; // @[Map2T.scala 17:7]
  assign O_0_1_0 = op_O_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_1_1 = op_O_0_1_1; // @[Map2T.scala 17:7]
  assign O_0_1_2 = op_O_0_1_2; // @[Map2T.scala 17:7]
  assign O_1_0_0 = op_O_1_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_1 = op_O_1_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_2 = op_O_1_0_2; // @[Map2T.scala 17:7]
  assign O_1_1_0 = op_O_1_1_0; // @[Map2T.scala 17:7]
  assign O_1_1_1 = op_O_1_1_1; // @[Map2T.scala 17:7]
  assign O_1_1_2 = op_O_1_1_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0 = I0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1 = I0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_2 = I0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0 = I0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1 = I0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_1_2 = I0_1_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0 = I1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_1 = I1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_0_2 = I1_0_2; // @[Map2T.scala 16:11]
  assign op_I1_1_0 = I1_1_0; // @[Map2T.scala 16:11]
  assign op_I1_1_1 = I1_1_1; // @[Map2T.scala 16:11]
  assign op_I1_1_2 = I1_1_2; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleAppender_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_0_2,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_1_2,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0_0 = I0_0_0; // @[Tuple.scala 24:34]
  assign O_0_1 = I0_0_1; // @[Tuple.scala 24:34]
  assign O_0_2 = I0_0_2; // @[Tuple.scala 24:34]
  assign O_1_0 = I0_1_0; // @[Tuple.scala 24:34]
  assign O_1_1 = I0_1_1; // @[Tuple.scala 24:34]
  assign O_1_2 = I0_1_2; // @[Tuple.scala 24:34]
  assign O_2_0 = I1_0; // @[Tuple.scala 26:32]
  assign O_2_1 = I1_1; // @[Tuple.scala 26:32]
  assign O_2_2 = I1_2; // @[Tuple.scala 26:32]
endmodule
module Map2S_7(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_0_0_1,
  input  [7:0] I0_0_0_2,
  input  [7:0] I0_0_1_0,
  input  [7:0] I0_0_1_1,
  input  [7:0] I0_0_1_2,
  input  [7:0] I0_1_0_0,
  input  [7:0] I0_1_0_1,
  input  [7:0] I0_1_0_2,
  input  [7:0] I0_1_1_0,
  input  [7:0] I0_1_1_1,
  input  [7:0] I0_1_1_2,
  input  [7:0] I1_0_0,
  input  [7:0] I1_0_1,
  input  [7:0] I1_0_2,
  input  [7:0] I1_1_0,
  input  [7:0] I1_1_1,
  input  [7:0] I1_1_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_0_2_0,
  output [7:0] O_0_2_1,
  output [7:0] O_0_2_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2,
  output [7:0] O_1_2_0,
  output [7:0] O_1_2_1,
  output [7:0] O_1_2_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_2; // @[Map2S.scala 10:86]
  SSeqTupleAppender_3 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I0_0_2(fst_op_I0_0_2),
    .I0_1_0(fst_op_I0_1_0),
    .I0_1_1(fst_op_I0_1_1),
    .I0_1_2(fst_op_I0_1_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0(other_ops_0_I0_0_0),
    .I0_0_1(other_ops_0_I0_0_1),
    .I0_0_2(other_ops_0_I0_0_2),
    .I0_1_0(other_ops_0_I0_1_0),
    .I0_1_1(other_ops_0_I0_1_1),
    .I0_1_2(other_ops_0_I0_1_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2),
    .O_2_0(other_ops_0_O_2_0),
    .O_2_1(other_ops_0_O_2_1),
    .O_2_2(other_ops_0_O_2_2)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[Map2S.scala 19:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[Map2S.scala 19:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[Map2S.scala 24:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[Map2S.scala 24:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[Map2S.scala 24:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[Map2S.scala 24:12]
  assign O_1_2_0 = other_ops_0_O_2_0; // @[Map2S.scala 24:12]
  assign O_1_2_1 = other_ops_0_O_2_1; // @[Map2S.scala 24:12]
  assign O_1_2_2 = other_ops_0_O_2_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_2 = I0_0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_0 = I0_0_1_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_1 = I0_0_1_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_2 = I0_0_1_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0 = I0_1_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_1 = I0_1_0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_2 = I0_1_0_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_0 = I0_1_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_1 = I0_1_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_2 = I0_1_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = I1_1_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = I1_1_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = I1_1_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_7(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_0_0_1,
  input  [7:0] I0_0_0_2,
  input  [7:0] I0_0_1_0,
  input  [7:0] I0_0_1_1,
  input  [7:0] I0_0_1_2,
  input  [7:0] I0_1_0_0,
  input  [7:0] I0_1_0_1,
  input  [7:0] I0_1_0_2,
  input  [7:0] I0_1_1_0,
  input  [7:0] I0_1_1_1,
  input  [7:0] I0_1_1_2,
  input  [7:0] I1_0_0,
  input  [7:0] I1_0_1,
  input  [7:0] I1_0_2,
  input  [7:0] I1_1_0,
  input  [7:0] I1_1_1,
  input  [7:0] I1_1_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_0_2_0,
  output [7:0] O_0_2_1,
  output [7:0] O_0_2_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2,
  output [7:0] O_1_2_0,
  output [7:0] O_1_2_1,
  output [7:0] O_1_2_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_2_2; // @[Map2T.scala 8:20]
  Map2S_7 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0_0(op_I0_0_0_0),
    .I0_0_0_1(op_I0_0_0_1),
    .I0_0_0_2(op_I0_0_0_2),
    .I0_0_1_0(op_I0_0_1_0),
    .I0_0_1_1(op_I0_0_1_1),
    .I0_0_1_2(op_I0_0_1_2),
    .I0_1_0_0(op_I0_1_0_0),
    .I0_1_0_1(op_I0_1_0_1),
    .I0_1_0_2(op_I0_1_0_2),
    .I0_1_1_0(op_I0_1_1_0),
    .I0_1_1_1(op_I0_1_1_1),
    .I0_1_1_2(op_I0_1_1_2),
    .I1_0_0(op_I1_0_0),
    .I1_0_1(op_I1_0_1),
    .I1_0_2(op_I1_0_2),
    .I1_1_0(op_I1_1_0),
    .I1_1_1(op_I1_1_1),
    .I1_1_2(op_I1_1_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_0_2_0(op_O_0_2_0),
    .O_0_2_1(op_O_0_2_1),
    .O_0_2_2(op_O_0_2_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_1_2_0(op_O_1_2_0),
    .O_1_2_1(op_O_1_2_1),
    .O_1_2_2(op_O_1_2_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0 = op_O_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_1 = op_O_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_2 = op_O_0_0_2; // @[Map2T.scala 17:7]
  assign O_0_1_0 = op_O_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_1_1 = op_O_0_1_1; // @[Map2T.scala 17:7]
  assign O_0_1_2 = op_O_0_1_2; // @[Map2T.scala 17:7]
  assign O_0_2_0 = op_O_0_2_0; // @[Map2T.scala 17:7]
  assign O_0_2_1 = op_O_0_2_1; // @[Map2T.scala 17:7]
  assign O_0_2_2 = op_O_0_2_2; // @[Map2T.scala 17:7]
  assign O_1_0_0 = op_O_1_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_1 = op_O_1_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_2 = op_O_1_0_2; // @[Map2T.scala 17:7]
  assign O_1_1_0 = op_O_1_1_0; // @[Map2T.scala 17:7]
  assign O_1_1_1 = op_O_1_1_1; // @[Map2T.scala 17:7]
  assign O_1_1_2 = op_O_1_1_2; // @[Map2T.scala 17:7]
  assign O_1_2_0 = op_O_1_2_0; // @[Map2T.scala 17:7]
  assign O_1_2_1 = op_O_1_2_1; // @[Map2T.scala 17:7]
  assign O_1_2_2 = op_O_1_2_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0_0 = I0_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_0_1 = I0_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_0_2 = I0_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_0_1_0 = I0_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1_1 = I0_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_0_1_2 = I0_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0 = I0_1_0_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_1 = I0_1_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0_2 = I0_1_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_1_0 = I0_1_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1_1 = I0_1_1_1; // @[Map2T.scala 15:11]
  assign op_I0_1_1_2 = I0_1_1_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0 = I1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_1 = I1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_0_2 = I1_0_2; // @[Map2T.scala 16:11]
  assign op_I1_1_0 = I1_1_0; // @[Map2T.scala 16:11]
  assign op_I1_1_1 = I1_1_1; // @[Map2T.scala 16:11]
  assign op_I1_1_2 = I1_1_2; // @[Map2T.scala 16:11]
endmodule
module PartitionS_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  input  [7:0] I_1_1_0,
  input  [7:0] I_1_1_1,
  input  [7:0] I_1_1_2,
  input  [7:0] I_1_2_0,
  input  [7:0] I_1_2_1,
  input  [7:0] I_1_2_2,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_0_2,
  output [7:0] O_0_0_1_0,
  output [7:0] O_0_0_1_1,
  output [7:0] O_0_0_1_2,
  output [7:0] O_0_0_2_0,
  output [7:0] O_0_0_2_1,
  output [7:0] O_0_0_2_2,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_0_2,
  output [7:0] O_1_0_1_0,
  output [7:0] O_1_0_1_1,
  output [7:0] O_1_0_1_2,
  output [7:0] O_1_0_2_0,
  output [7:0] O_1_0_2_1,
  output [7:0] O_1_0_2_2
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0_0 = I_0_0_0; // @[Partition.scala 15:39]
  assign O_0_0_0_1 = I_0_0_1; // @[Partition.scala 15:39]
  assign O_0_0_0_2 = I_0_0_2; // @[Partition.scala 15:39]
  assign O_0_0_1_0 = I_0_1_0; // @[Partition.scala 15:39]
  assign O_0_0_1_1 = I_0_1_1; // @[Partition.scala 15:39]
  assign O_0_0_1_2 = I_0_1_2; // @[Partition.scala 15:39]
  assign O_0_0_2_0 = I_0_2_0; // @[Partition.scala 15:39]
  assign O_0_0_2_1 = I_0_2_1; // @[Partition.scala 15:39]
  assign O_0_0_2_2 = I_0_2_2; // @[Partition.scala 15:39]
  assign O_1_0_0_0 = I_1_0_0; // @[Partition.scala 15:39]
  assign O_1_0_0_1 = I_1_0_1; // @[Partition.scala 15:39]
  assign O_1_0_0_2 = I_1_0_2; // @[Partition.scala 15:39]
  assign O_1_0_1_0 = I_1_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1_1 = I_1_1_1; // @[Partition.scala 15:39]
  assign O_1_0_1_2 = I_1_1_2; // @[Partition.scala 15:39]
  assign O_1_0_2_0 = I_1_2_0; // @[Partition.scala 15:39]
  assign O_1_0_2_1 = I_1_2_1; // @[Partition.scala 15:39]
  assign O_1_0_2_2 = I_1_2_2; // @[Partition.scala 15:39]
endmodule
module MapT_6(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  input  [7:0] I_1_1_0,
  input  [7:0] I_1_1_1,
  input  [7:0] I_1_1_2,
  input  [7:0] I_1_2_0,
  input  [7:0] I_1_2_1,
  input  [7:0] I_1_2_2,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_0_2,
  output [7:0] O_0_0_1_0,
  output [7:0] O_0_0_1_1,
  output [7:0] O_0_0_1_2,
  output [7:0] O_0_0_2_0,
  output [7:0] O_0_0_2_1,
  output [7:0] O_0_0_2_2,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_0_2,
  output [7:0] O_1_0_1_0,
  output [7:0] O_1_0_1_1,
  output [7:0] O_1_0_1_2,
  output [7:0] O_1_0_2_0,
  output [7:0] O_1_0_2_1,
  output [7:0] O_1_0_2_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_2_2; // @[MapT.scala 8:20]
  PartitionS_3 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .O_0_0_0_0(op_O_0_0_0_0),
    .O_0_0_0_1(op_O_0_0_0_1),
    .O_0_0_0_2(op_O_0_0_0_2),
    .O_0_0_1_0(op_O_0_0_1_0),
    .O_0_0_1_1(op_O_0_0_1_1),
    .O_0_0_1_2(op_O_0_0_1_2),
    .O_0_0_2_0(op_O_0_0_2_0),
    .O_0_0_2_1(op_O_0_0_2_1),
    .O_0_0_2_2(op_O_0_0_2_2),
    .O_1_0_0_0(op_O_1_0_0_0),
    .O_1_0_0_1(op_O_1_0_0_1),
    .O_1_0_0_2(op_O_1_0_0_2),
    .O_1_0_1_0(op_O_1_0_1_0),
    .O_1_0_1_1(op_O_1_0_1_1),
    .O_1_0_1_2(op_O_1_0_1_2),
    .O_1_0_2_0(op_O_1_0_2_0),
    .O_1_0_2_1(op_O_1_0_2_1),
    .O_1_0_2_2(op_O_1_0_2_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0_0 = op_O_0_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_0_1 = op_O_0_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_0_2 = op_O_0_0_0_2; // @[MapT.scala 15:7]
  assign O_0_0_1_0 = op_O_0_0_1_0; // @[MapT.scala 15:7]
  assign O_0_0_1_1 = op_O_0_0_1_1; // @[MapT.scala 15:7]
  assign O_0_0_1_2 = op_O_0_0_1_2; // @[MapT.scala 15:7]
  assign O_0_0_2_0 = op_O_0_0_2_0; // @[MapT.scala 15:7]
  assign O_0_0_2_1 = op_O_0_0_2_1; // @[MapT.scala 15:7]
  assign O_0_0_2_2 = op_O_0_0_2_2; // @[MapT.scala 15:7]
  assign O_1_0_0_0 = op_O_1_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0_1 = op_O_1_0_0_1; // @[MapT.scala 15:7]
  assign O_1_0_0_2 = op_O_1_0_0_2; // @[MapT.scala 15:7]
  assign O_1_0_1_0 = op_O_1_0_1_0; // @[MapT.scala 15:7]
  assign O_1_0_1_1 = op_O_1_0_1_1; // @[MapT.scala 15:7]
  assign O_1_0_1_2 = op_O_1_0_1_2; // @[MapT.scala 15:7]
  assign O_1_0_2_0 = op_O_1_0_2_0; // @[MapT.scala 15:7]
  assign O_1_0_2_1 = op_O_1_0_2_1; // @[MapT.scala 15:7]
  assign O_1_0_2_2 = op_O_1_0_2_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleToSSeq_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_2_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0_0 = I_0_0; // @[Tuple.scala 41:5]
  assign O_0_1 = I_0_1; // @[Tuple.scala 41:5]
  assign O_0_2 = I_0_2; // @[Tuple.scala 41:5]
  assign O_1_0 = I_1_0; // @[Tuple.scala 41:5]
  assign O_1_1 = I_1_1; // @[Tuple.scala 41:5]
  assign O_1_2 = I_1_2; // @[Tuple.scala 41:5]
  assign O_2_0 = I_2_0; // @[Tuple.scala 41:5]
  assign O_2_1 = I_2_1; // @[Tuple.scala 41:5]
  assign O_2_2 = I_2_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq_3 op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0_0(op_inst_I_0_0),
    .I_0_1(op_inst_I_0_1),
    .I_0_2(op_inst_I_0_2),
    .I_1_0(op_inst_I_1_0),
    .I_1_1(op_inst_I_1_1),
    .I_1_2(op_inst_I_1_2),
    .I_2_0(op_inst_I_2_0),
    .I_2_1(op_inst_I_2_1),
    .I_2_2(op_inst_I_2_2),
    .O_0_0(op_inst_O_0_0),
    .O_0_1(op_inst_O_0_1),
    .O_0_2(op_inst_O_0_2),
    .O_1_0(op_inst_O_1_0),
    .O_1_1(op_inst_O_1_1),
    .O_1_2(op_inst_O_1_2),
    .O_2_0(op_inst_O_2_0),
    .O_2_1(op_inst_O_2_1),
    .O_2_2(op_inst_O_2_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0_0 = op_inst_O_0_0; // @[Remove1S.scala 14:5]
  assign O_0_1 = op_inst_O_0_1; // @[Remove1S.scala 14:5]
  assign O_0_2 = op_inst_O_0_2; // @[Remove1S.scala 14:5]
  assign O_1_0 = op_inst_O_1_0; // @[Remove1S.scala 14:5]
  assign O_1_1 = op_inst_O_1_1; // @[Remove1S.scala 14:5]
  assign O_1_2 = op_inst_O_1_2; // @[Remove1S.scala 14:5]
  assign O_2_0 = op_inst_O_2_0; // @[Remove1S.scala 14:5]
  assign O_2_1 = op_inst_O_2_1; // @[Remove1S.scala 14:5]
  assign O_2_2 = op_inst_O_2_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0_0 = I_0_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_1 = I_0_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_2 = I_0_0_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_0 = I_0_1_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_1 = I_0_1_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_2 = I_0_1_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_0 = I_0_2_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_1 = I_0_2_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_2 = I_0_2_2; // @[Remove1S.scala 13:13]
endmodule
module MapS_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0_0,
  input  [7:0] I_0_0_0_1,
  input  [7:0] I_0_0_0_2,
  input  [7:0] I_0_0_1_0,
  input  [7:0] I_0_0_1_1,
  input  [7:0] I_0_0_1_2,
  input  [7:0] I_0_0_2_0,
  input  [7:0] I_0_0_2_1,
  input  [7:0] I_0_0_2_2,
  input  [7:0] I_1_0_0_0,
  input  [7:0] I_1_0_0_1,
  input  [7:0] I_1_0_0_2,
  input  [7:0] I_1_0_1_0,
  input  [7:0] I_1_0_1_1,
  input  [7:0] I_1_0_1_2,
  input  [7:0] I_1_0_2_0,
  input  [7:0] I_1_0_2_1,
  input  [7:0] I_1_0_2_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_0_2_0,
  output [7:0] O_0_2_1,
  output [7:0] O_0_2_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2,
  output [7:0] O_1_2_0,
  output [7:0] O_1_2_1,
  output [7:0] O_1_2_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2_2; // @[MapS.scala 10:86]
  Remove1S_3 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0_0(fst_op_I_0_0_0),
    .I_0_0_1(fst_op_I_0_0_1),
    .I_0_0_2(fst_op_I_0_0_2),
    .I_0_1_0(fst_op_I_0_1_0),
    .I_0_1_1(fst_op_I_0_1_1),
    .I_0_1_2(fst_op_I_0_1_2),
    .I_0_2_0(fst_op_I_0_2_0),
    .I_0_2_1(fst_op_I_0_2_1),
    .I_0_2_2(fst_op_I_0_2_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  Remove1S_3 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0_0(other_ops_0_I_0_0_0),
    .I_0_0_1(other_ops_0_I_0_0_1),
    .I_0_0_2(other_ops_0_I_0_0_2),
    .I_0_1_0(other_ops_0_I_0_1_0),
    .I_0_1_1(other_ops_0_I_0_1_1),
    .I_0_1_2(other_ops_0_I_0_1_2),
    .I_0_2_0(other_ops_0_I_0_2_0),
    .I_0_2_1(other_ops_0_I_0_2_1),
    .I_0_2_2(other_ops_0_I_0_2_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2),
    .O_2_0(other_ops_0_O_2_0),
    .O_2_1(other_ops_0_O_2_1),
    .O_2_2(other_ops_0_O_2_2)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[MapS.scala 17:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[MapS.scala 17:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[MapS.scala 17:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[MapS.scala 17:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[MapS.scala 17:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[MapS.scala 17:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[MapS.scala 17:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[MapS.scala 21:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[MapS.scala 21:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[MapS.scala 21:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[MapS.scala 21:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[MapS.scala 21:12]
  assign O_1_2_0 = other_ops_0_O_2_0; // @[MapS.scala 21:12]
  assign O_1_2_1 = other_ops_0_O_2_1; // @[MapS.scala 21:12]
  assign O_1_2_2 = other_ops_0_O_2_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0_0 = I_0_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_1 = I_0_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_2 = I_0_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_0 = I_0_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_1 = I_0_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_2 = I_0_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_0 = I_0_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_1 = I_0_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_2 = I_0_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0_0 = I_1_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_1 = I_1_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_2 = I_1_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_0 = I_1_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_1 = I_1_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_2 = I_1_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_0 = I_1_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_1 = I_1_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_2 = I_1_0_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_7(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0_0,
  input  [7:0] I_0_0_0_1,
  input  [7:0] I_0_0_0_2,
  input  [7:0] I_0_0_1_0,
  input  [7:0] I_0_0_1_1,
  input  [7:0] I_0_0_1_2,
  input  [7:0] I_0_0_2_0,
  input  [7:0] I_0_0_2_1,
  input  [7:0] I_0_0_2_2,
  input  [7:0] I_1_0_0_0,
  input  [7:0] I_1_0_0_1,
  input  [7:0] I_1_0_0_2,
  input  [7:0] I_1_0_1_0,
  input  [7:0] I_1_0_1_1,
  input  [7:0] I_1_0_1_2,
  input  [7:0] I_1_0_2_0,
  input  [7:0] I_1_0_2_1,
  input  [7:0] I_1_0_2_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_0_2_0,
  output [7:0] O_0_2_1,
  output [7:0] O_0_2_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2,
  output [7:0] O_1_2_0,
  output [7:0] O_1_2_1,
  output [7:0] O_1_2_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_2_2; // @[MapT.scala 8:20]
  MapS_3 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0_0(op_I_0_0_0_0),
    .I_0_0_0_1(op_I_0_0_0_1),
    .I_0_0_0_2(op_I_0_0_0_2),
    .I_0_0_1_0(op_I_0_0_1_0),
    .I_0_0_1_1(op_I_0_0_1_1),
    .I_0_0_1_2(op_I_0_0_1_2),
    .I_0_0_2_0(op_I_0_0_2_0),
    .I_0_0_2_1(op_I_0_0_2_1),
    .I_0_0_2_2(op_I_0_0_2_2),
    .I_1_0_0_0(op_I_1_0_0_0),
    .I_1_0_0_1(op_I_1_0_0_1),
    .I_1_0_0_2(op_I_1_0_0_2),
    .I_1_0_1_0(op_I_1_0_1_0),
    .I_1_0_1_1(op_I_1_0_1_1),
    .I_1_0_1_2(op_I_1_0_1_2),
    .I_1_0_2_0(op_I_1_0_2_0),
    .I_1_0_2_1(op_I_1_0_2_1),
    .I_1_0_2_2(op_I_1_0_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_0_2_0(op_O_0_2_0),
    .O_0_2_1(op_O_0_2_1),
    .O_0_2_2(op_O_0_2_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_1_2_0(op_O_1_2_0),
    .O_1_2_1(op_O_1_2_1),
    .O_1_2_2(op_O_1_2_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_2 = op_O_0_0_2; // @[MapT.scala 15:7]
  assign O_0_1_0 = op_O_0_1_0; // @[MapT.scala 15:7]
  assign O_0_1_1 = op_O_0_1_1; // @[MapT.scala 15:7]
  assign O_0_1_2 = op_O_0_1_2; // @[MapT.scala 15:7]
  assign O_0_2_0 = op_O_0_2_0; // @[MapT.scala 15:7]
  assign O_0_2_1 = op_O_0_2_1; // @[MapT.scala 15:7]
  assign O_0_2_2 = op_O_0_2_2; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_0_2 = op_O_1_0_2; // @[MapT.scala 15:7]
  assign O_1_1_0 = op_O_1_1_0; // @[MapT.scala 15:7]
  assign O_1_1_1 = op_O_1_1_1; // @[MapT.scala 15:7]
  assign O_1_1_2 = op_O_1_1_2; // @[MapT.scala 15:7]
  assign O_1_2_0 = op_O_1_2_0; // @[MapT.scala 15:7]
  assign O_1_2_1 = op_O_1_2_1; // @[MapT.scala 15:7]
  assign O_1_2_2 = op_O_1_2_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0_0 = I_0_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_0_1 = I_0_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_0_2 = I_0_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_0_1_0 = I_0_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1_1 = I_0_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_0_1_2 = I_0_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_0_2_0 = I_0_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_0_2_1 = I_0_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2_2 = I_0_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0_0 = I_1_0_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_0_1 = I_1_0_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0_2 = I_1_0_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0_1_0 = I_1_0_1_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1_1 = I_1_0_1_1; // @[MapT.scala 14:10]
  assign op_I_1_0_1_2 = I_1_0_1_2; // @[MapT.scala 14:10]
  assign op_I_1_0_2_0 = I_1_0_2_0; // @[MapT.scala 14:10]
  assign op_I_1_0_2_1 = I_1_0_2_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2_2 = I_1_0_2_2; // @[MapT.scala 14:10]
endmodule
module InitialDelayCounter(
  input   clock,
  input   reset,
  output  valid_down
);
  reg  value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire  _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 1'h1; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 1'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 1'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module AtomTuple(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  input  [7:0] I1,
  output [7:0] O_t0b,
  output [7:0] O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b = I1; // @[Tuple.scala 50:9]
endmodule
module Map2S_8(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I0_2,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  output [7:0] O_0_t0b,
  output [7:0] O_0_t1b,
  output [7:0] O_1_t0b,
  output [7:0] O_1_t1b,
  output [7:0] O_2_t0b,
  output [7:0] O_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  AtomTuple other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_t0b(other_ops_0_O_t0b),
    .O_t1b(other_ops_0_O_t1b)
  );
  AtomTuple other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_t0b(other_ops_1_O_t0b),
    .O_t1b(other_ops_1_O_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign O_1_t0b = other_ops_0_O_t0b; // @[Map2S.scala 24:12]
  assign O_1_t1b = other_ops_0_O_t1b; // @[Map2S.scala 24:12]
  assign O_2_t0b = other_ops_1_O_t0b; // @[Map2S.scala 24:12]
  assign O_2_t1b = other_ops_1_O_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
endmodule
module Map2S_9(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_0_2,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_1_2,
  input  [7:0] I0_2_0,
  input  [7:0] I0_2_1,
  input  [7:0] I0_2_2,
  output [7:0] O_0_0_t0b,
  output [7:0] O_0_0_t1b,
  output [7:0] O_0_1_t0b,
  output [7:0] O_0_1_t1b,
  output [7:0] O_0_2_t0b,
  output [7:0] O_0_2_t1b,
  output [7:0] O_1_0_t0b,
  output [7:0] O_1_0_t1b,
  output [7:0] O_1_1_t0b,
  output [7:0] O_1_1_t1b,
  output [7:0] O_1_2_t0b,
  output [7:0] O_1_2_t1b,
  output [7:0] O_2_0_t0b,
  output [7:0] O_2_0_t1b,
  output [7:0] O_2_1_t0b,
  output [7:0] O_2_1_t1b,
  output [7:0] O_2_2_t0b,
  output [7:0] O_2_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_t1b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  Map2S_8 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b),
    .O_1_t0b(fst_op_O_1_t0b),
    .O_1_t1b(fst_op_O_1_t1b),
    .O_2_t0b(fst_op_O_2_t0b),
    .O_2_t1b(fst_op_O_2_t1b)
  );
  Map2S_8 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I0_2(other_ops_0_I0_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_t0b(other_ops_0_O_0_t0b),
    .O_0_t1b(other_ops_0_O_0_t1b),
    .O_1_t0b(other_ops_0_O_1_t0b),
    .O_1_t1b(other_ops_0_O_1_t1b),
    .O_2_t0b(other_ops_0_O_2_t0b),
    .O_2_t1b(other_ops_0_O_2_t1b)
  );
  Map2S_8 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I0_2(other_ops_1_I0_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_t0b(other_ops_1_O_0_t0b),
    .O_0_t1b(other_ops_1_O_0_t1b),
    .O_1_t0b(other_ops_1_O_1_t0b),
    .O_1_t1b(other_ops_1_O_1_t1b),
    .O_2_t0b(other_ops_1_O_2_t0b),
    .O_2_t1b(other_ops_1_O_2_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign O_0_1_t0b = fst_op_O_1_t0b; // @[Map2S.scala 19:8]
  assign O_0_1_t1b = fst_op_O_1_t1b; // @[Map2S.scala 19:8]
  assign O_0_2_t0b = fst_op_O_2_t0b; // @[Map2S.scala 19:8]
  assign O_0_2_t1b = fst_op_O_2_t1b; // @[Map2S.scala 19:8]
  assign O_1_0_t0b = other_ops_0_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_1_0_t1b = other_ops_0_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_1_1_t0b = other_ops_0_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_1_1_t1b = other_ops_0_O_1_t1b; // @[Map2S.scala 24:12]
  assign O_1_2_t0b = other_ops_0_O_2_t0b; // @[Map2S.scala 24:12]
  assign O_1_2_t1b = other_ops_0_O_2_t1b; // @[Map2S.scala 24:12]
  assign O_2_0_t0b = other_ops_1_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_2_0_t1b = other_ops_1_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_2_1_t0b = other_ops_1_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_2_1_t1b = other_ops_1_O_1_t1b; // @[Map2S.scala 24:12]
  assign O_2_2_t0b = other_ops_1_O_2_t0b; // @[Map2S.scala 24:12]
  assign O_2_2_t1b = other_ops_1_O_2_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = 8'h1; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = 8'h2; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = 8'h1; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2 = I0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = 8'h2; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = 8'h4; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = 8'h2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2 = I0_2_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = 8'h1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = 8'h2; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = 8'h1; // @[Map2S.scala 23:43]
endmodule
module Mul(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  wire [7:0] BlackBoxMulUInt8_I0; // @[Arithmetic.scala 165:27]
  wire [7:0] BlackBoxMulUInt8_I1; // @[Arithmetic.scala 165:27]
  wire [15:0] BlackBoxMulUInt8_O; // @[Arithmetic.scala 165:27]
  wire  BlackBoxMulUInt8_clock; // @[Arithmetic.scala 165:27]
  reg  _T_1; // @[Arithmetic.scala 217:42]
  reg [31:0] _RAND_0;
  reg  _T_2; // @[Arithmetic.scala 217:34]
  reg [31:0] _RAND_1;
  reg  _T_3; // @[Arithmetic.scala 217:26]
  reg [31:0] _RAND_2;
  BlackBoxMulUInt8 BlackBoxMulUInt8 ( // @[Arithmetic.scala 165:27]
    .I0(BlackBoxMulUInt8_I0),
    .I1(BlackBoxMulUInt8_I1),
    .O(BlackBoxMulUInt8_O),
    .clock(BlackBoxMulUInt8_clock)
  );
  assign valid_down = _T_3; // @[Arithmetic.scala 217:16]
  assign O = BlackBoxMulUInt8_O[7:0]; // @[Arithmetic.scala 168:7]
  assign BlackBoxMulUInt8_I0 = I_t0b; // @[Arithmetic.scala 166:21]
  assign BlackBoxMulUInt8_I1 = I_t1b; // @[Arithmetic.scala 167:21]
  assign BlackBoxMulUInt8_clock = clock; // @[Arithmetic.scala 169:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_2 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_3 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
    if (reset) begin
      _T_2 <= 1'h0;
    end else begin
      _T_2 <= _T_1;
    end
    if (reset) begin
      _T_3 <= 1'h0;
    end else begin
      _T_3 <= _T_2;
    end
  end
endmodule
module MapS_4(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  input  [7:0] I_1_t0b,
  input  [7:0] I_1_t1b,
  input  [7:0] I_2_t0b,
  input  [7:0] I_2_t1b,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  Mul fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  Mul other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_t0b(other_ops_0_I_t0b),
    .I_t1b(other_ops_0_I_t1b),
    .O(other_ops_0_O)
  );
  Mul other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_t0b(other_ops_1_I_t0b),
    .I_t1b(other_ops_1_I_t1b),
    .O(other_ops_1_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_t0b = I_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_t1b = I_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_t0b = I_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_t1b = I_2_t1b; // @[MapS.scala 20:41]
endmodule
module MapS_5(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_t0b,
  input  [7:0] I_0_0_t1b,
  input  [7:0] I_0_1_t0b,
  input  [7:0] I_0_1_t1b,
  input  [7:0] I_0_2_t0b,
  input  [7:0] I_0_2_t1b,
  input  [7:0] I_1_0_t0b,
  input  [7:0] I_1_0_t1b,
  input  [7:0] I_1_1_t0b,
  input  [7:0] I_1_1_t1b,
  input  [7:0] I_1_2_t0b,
  input  [7:0] I_1_2_t1b,
  input  [7:0] I_2_0_t0b,
  input  [7:0] I_2_0_t1b,
  input  [7:0] I_2_1_t0b,
  input  [7:0] I_2_1_t1b,
  input  [7:0] I_2_2_t0b,
  input  [7:0] I_2_2_t1b,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  MapS_4 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .I_1_t0b(fst_op_I_1_t0b),
    .I_1_t1b(fst_op_I_1_t1b),
    .I_2_t0b(fst_op_I_2_t0b),
    .I_2_t1b(fst_op_I_2_t1b),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  MapS_4 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_t0b(other_ops_0_I_0_t0b),
    .I_0_t1b(other_ops_0_I_0_t1b),
    .I_1_t0b(other_ops_0_I_1_t0b),
    .I_1_t1b(other_ops_0_I_1_t1b),
    .I_2_t0b(other_ops_0_I_2_t0b),
    .I_2_t1b(other_ops_0_I_2_t1b),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  MapS_4 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_t0b(other_ops_1_I_0_t0b),
    .I_0_t1b(other_ops_1_I_0_t1b),
    .I_1_t0b(other_ops_1_I_1_t0b),
    .I_1_t1b(other_ops_1_I_1_t1b),
    .I_2_t0b(other_ops_1_I_2_t0b),
    .I_2_t1b(other_ops_1_I_2_t1b),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_1_2 = other_ops_0_O_2; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign O_2_1 = other_ops_1_O_1; // @[MapS.scala 21:12]
  assign O_2_2 = other_ops_1_O_2; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t0b = I_0_1_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t1b = I_0_1_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_2_t0b = I_0_2_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_2_t1b = I_0_2_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_t0b = I_1_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_t1b = I_1_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t0b = I_1_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t1b = I_1_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_t0b = I_1_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_t1b = I_1_2_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_t0b = I_2_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_t1b = I_2_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_t0b = I_2_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_t1b = I_2_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_t0b = I_2_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_t1b = I_2_2_t1b; // @[MapS.scala 20:41]
endmodule
module AddNoValid(
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  assign O = I_t0b + I_t1b; // @[Arithmetic.scala 122:7]
endmodule
module ReduceS(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  output [7:0] O_0
);
  wire [7:0] AddNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_O; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_1_I_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_1_I_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_1_O; // @[ReduceS.scala 20:43]
  reg [7:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg [7:0] _T_1; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_1;
  reg [7:0] _T_2; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_2;
  reg [7:0] _T_3; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_3;
  reg  _T_4; // @[ReduceS.scala 47:32]
  reg [31:0] _RAND_4;
  reg  _T_5; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_5;
  AddNoValid AddNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  AddNoValid AddNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_1_I_t0b),
    .I_t1b(AddNoValid_1_I_t1b),
    .O(AddNoValid_1_O)
  );
  assign valid_down = _T_5; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign AddNoValid_I_t0b = _T_1; // @[ReduceS.scala 43:18]
  assign AddNoValid_I_t1b = AddNoValid_1_O; // @[ReduceS.scala 36:18]
  assign AddNoValid_1_I_t0b = _T_3; // @[ReduceS.scala 43:18]
  assign AddNoValid_1_I_t1b = _T_2; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= AddNoValid_O;
    _T_1 <= I_0;
    _T_2 <= I_1;
    _T_3 <= I_2;
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= valid_up;
    end
    _T_5 <= _T_4;
  end
endmodule
module MapS_6(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_2_2,
  output [7:0] O_0_0,
  output [7:0] O_1_0,
  output [7:0] O_2_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  ReduceS fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .I_2(fst_op_I_2),
    .O_0(fst_op_O_0)
  );
  ReduceS other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0(other_ops_0_I_0),
    .I_1(other_ops_0_I_1),
    .I_2(other_ops_0_I_2),
    .O_0(other_ops_0_O_0)
  );
  ReduceS other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0(other_ops_1_I_0),
    .I_1(other_ops_1_I_1),
    .I_2(other_ops_1_I_2),
    .O_0(other_ops_1_O_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_2 = I_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0 = I_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1 = I_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2 = I_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0 = I_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1 = I_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2 = I_2_2; // @[MapS.scala 20:41]
endmodule
module MapSNoValid(
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  output [7:0] O_0
);
  wire [7:0] fst_op_I_t0b; // @[MapS.scala 28:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 28:22]
  wire [7:0] fst_op_O; // @[MapS.scala 28:22]
  AddNoValid fst_op ( // @[MapS.scala 28:22]
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign O_0 = fst_op_O; // @[MapS.scala 35:8]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 34:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 34:12]
endmodule
module ReduceS_1(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_1_0,
  input  [7:0] I_2_0,
  output [7:0] O_0_0
);
  wire [7:0] MapSNoValid_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_O_0; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_1_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_1_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_1_O_0; // @[ReduceS.scala 20:43]
  reg [7:0] _T_0; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg [7:0] _T_1_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_1;
  reg [7:0] _T_2_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_2;
  reg [7:0] _T_3_0; // @[ReduceS.scala 43:46]
  reg [31:0] _RAND_3;
  reg  _T_4; // @[ReduceS.scala 47:32]
  reg [31:0] _RAND_4;
  reg  _T_5; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_5;
  MapSNoValid MapSNoValid ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_I_0_t0b),
    .I_0_t1b(MapSNoValid_I_0_t1b),
    .O_0(MapSNoValid_O_0)
  );
  MapSNoValid MapSNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_1_I_0_t0b),
    .I_0_t1b(MapSNoValid_1_I_0_t1b),
    .O_0(MapSNoValid_1_O_0)
  );
  assign valid_down = _T_5; // @[ReduceS.scala 47:14]
  assign O_0_0 = _T_0; // @[ReduceS.scala 27:14]
  assign MapSNoValid_I_0_t0b = _T_1_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_I_0_t1b = MapSNoValid_1_O_0; // @[ReduceS.scala 36:18]
  assign MapSNoValid_1_I_0_t0b = _T_3_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_1_I_0_t1b = _T_2_0; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1_0 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2_0 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3_0 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0 <= MapSNoValid_O_0;
    _T_1_0 <= I_0_0;
    _T_2_0 <= I_1_0;
    _T_3_0 <= I_2_0;
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= valid_up;
    end
    _T_5 <= _T_4;
  end
endmodule
module InitialDelayCounter_1(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [3:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [3:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 4'h8; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 4'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 4'h8; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 4'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module AtomTuple_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  output [7:0] O_t0b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
endmodule
module Map2S_10(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  output [7:0] O_0_t0b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  AtomTuple_1 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .O_t0b(fst_op_O_t0b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
endmodule
module Map2S_11(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  output [7:0] O_0_0_t0b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  Map2S_10 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .O_0_t0b(fst_op_O_0_t0b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
endmodule
module Div(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  output [7:0] O
);
  wire [7:0] BlackBoxMulUInt8_I0; // @[Arithmetic.scala 342:27]
  wire [7:0] BlackBoxMulUInt8_I1; // @[Arithmetic.scala 342:27]
  wire [15:0] BlackBoxMulUInt8_O; // @[Arithmetic.scala 342:27]
  wire  BlackBoxMulUInt8_clock; // @[Arithmetic.scala 342:27]
  reg  _T_3; // @[Arithmetic.scala 370:42]
  reg [31:0] _RAND_0;
  reg  _T_4; // @[Arithmetic.scala 370:34]
  reg [31:0] _RAND_1;
  reg  _T_5; // @[Arithmetic.scala 370:26]
  reg [31:0] _RAND_2;
  BlackBoxMulUInt8 BlackBoxMulUInt8 ( // @[Arithmetic.scala 342:27]
    .I0(BlackBoxMulUInt8_I0),
    .I1(BlackBoxMulUInt8_I1),
    .O(BlackBoxMulUInt8_O),
    .clock(BlackBoxMulUInt8_clock)
  );
  assign valid_down = _T_5; // @[Arithmetic.scala 370:16]
  assign O = BlackBoxMulUInt8_O[14:7]; // @[Arithmetic.scala 345:7]
  assign BlackBoxMulUInt8_I0 = I_t0b; // @[Arithmetic.scala 343:21]
  assign BlackBoxMulUInt8_I1 = 8'h8; // @[Arithmetic.scala 344:21]
  assign BlackBoxMulUInt8_clock = clock; // @[Arithmetic.scala 346:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_3 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_4 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_5 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_3 <= 1'h0;
    end else begin
      _T_3 <= valid_up;
    end
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= _T_3;
    end
    if (reset) begin
      _T_5 <= 1'h0;
    end else begin
      _T_5 <= _T_4;
    end
  end
endmodule
module MapS_7(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_t0b,
  output [7:0] O_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  Div fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
endmodule
module MapS_8(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_t0b,
  output [7:0] O_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  MapS_7 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
endmodule
module Module_0(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_2_2,
  output [7:0] O_0_0
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n110_valid_up; // @[Top.scala 18:22]
  wire  n110_valid_down; // @[Top.scala 18:22]
  wire [7:0] n110_I0_0_0; // @[Top.scala 18:22]
  wire [7:0] n110_I0_0_1; // @[Top.scala 18:22]
  wire [7:0] n110_I0_0_2; // @[Top.scala 18:22]
  wire [7:0] n110_I0_1_0; // @[Top.scala 18:22]
  wire [7:0] n110_I0_1_1; // @[Top.scala 18:22]
  wire [7:0] n110_I0_1_2; // @[Top.scala 18:22]
  wire [7:0] n110_I0_2_0; // @[Top.scala 18:22]
  wire [7:0] n110_I0_2_1; // @[Top.scala 18:22]
  wire [7:0] n110_I0_2_2; // @[Top.scala 18:22]
  wire [7:0] n110_O_0_0_t0b; // @[Top.scala 18:22]
  wire [7:0] n110_O_0_0_t1b; // @[Top.scala 18:22]
  wire [7:0] n110_O_0_1_t0b; // @[Top.scala 18:22]
  wire [7:0] n110_O_0_1_t1b; // @[Top.scala 18:22]
  wire [7:0] n110_O_0_2_t0b; // @[Top.scala 18:22]
  wire [7:0] n110_O_0_2_t1b; // @[Top.scala 18:22]
  wire [7:0] n110_O_1_0_t0b; // @[Top.scala 18:22]
  wire [7:0] n110_O_1_0_t1b; // @[Top.scala 18:22]
  wire [7:0] n110_O_1_1_t0b; // @[Top.scala 18:22]
  wire [7:0] n110_O_1_1_t1b; // @[Top.scala 18:22]
  wire [7:0] n110_O_1_2_t0b; // @[Top.scala 18:22]
  wire [7:0] n110_O_1_2_t1b; // @[Top.scala 18:22]
  wire [7:0] n110_O_2_0_t0b; // @[Top.scala 18:22]
  wire [7:0] n110_O_2_0_t1b; // @[Top.scala 18:22]
  wire [7:0] n110_O_2_1_t0b; // @[Top.scala 18:22]
  wire [7:0] n110_O_2_1_t1b; // @[Top.scala 18:22]
  wire [7:0] n110_O_2_2_t0b; // @[Top.scala 18:22]
  wire [7:0] n110_O_2_2_t1b; // @[Top.scala 18:22]
  wire  n121_clock; // @[Top.scala 22:22]
  wire  n121_reset; // @[Top.scala 22:22]
  wire  n121_valid_up; // @[Top.scala 22:22]
  wire  n121_valid_down; // @[Top.scala 22:22]
  wire [7:0] n121_I_0_0_t0b; // @[Top.scala 22:22]
  wire [7:0] n121_I_0_0_t1b; // @[Top.scala 22:22]
  wire [7:0] n121_I_0_1_t0b; // @[Top.scala 22:22]
  wire [7:0] n121_I_0_1_t1b; // @[Top.scala 22:22]
  wire [7:0] n121_I_0_2_t0b; // @[Top.scala 22:22]
  wire [7:0] n121_I_0_2_t1b; // @[Top.scala 22:22]
  wire [7:0] n121_I_1_0_t0b; // @[Top.scala 22:22]
  wire [7:0] n121_I_1_0_t1b; // @[Top.scala 22:22]
  wire [7:0] n121_I_1_1_t0b; // @[Top.scala 22:22]
  wire [7:0] n121_I_1_1_t1b; // @[Top.scala 22:22]
  wire [7:0] n121_I_1_2_t0b; // @[Top.scala 22:22]
  wire [7:0] n121_I_1_2_t1b; // @[Top.scala 22:22]
  wire [7:0] n121_I_2_0_t0b; // @[Top.scala 22:22]
  wire [7:0] n121_I_2_0_t1b; // @[Top.scala 22:22]
  wire [7:0] n121_I_2_1_t0b; // @[Top.scala 22:22]
  wire [7:0] n121_I_2_1_t1b; // @[Top.scala 22:22]
  wire [7:0] n121_I_2_2_t0b; // @[Top.scala 22:22]
  wire [7:0] n121_I_2_2_t1b; // @[Top.scala 22:22]
  wire [7:0] n121_O_0_0; // @[Top.scala 22:22]
  wire [7:0] n121_O_0_1; // @[Top.scala 22:22]
  wire [7:0] n121_O_0_2; // @[Top.scala 22:22]
  wire [7:0] n121_O_1_0; // @[Top.scala 22:22]
  wire [7:0] n121_O_1_1; // @[Top.scala 22:22]
  wire [7:0] n121_O_1_2; // @[Top.scala 22:22]
  wire [7:0] n121_O_2_0; // @[Top.scala 22:22]
  wire [7:0] n121_O_2_1; // @[Top.scala 22:22]
  wire [7:0] n121_O_2_2; // @[Top.scala 22:22]
  wire  n126_clock; // @[Top.scala 25:22]
  wire  n126_reset; // @[Top.scala 25:22]
  wire  n126_valid_up; // @[Top.scala 25:22]
  wire  n126_valid_down; // @[Top.scala 25:22]
  wire [7:0] n126_I_0_0; // @[Top.scala 25:22]
  wire [7:0] n126_I_0_1; // @[Top.scala 25:22]
  wire [7:0] n126_I_0_2; // @[Top.scala 25:22]
  wire [7:0] n126_I_1_0; // @[Top.scala 25:22]
  wire [7:0] n126_I_1_1; // @[Top.scala 25:22]
  wire [7:0] n126_I_1_2; // @[Top.scala 25:22]
  wire [7:0] n126_I_2_0; // @[Top.scala 25:22]
  wire [7:0] n126_I_2_1; // @[Top.scala 25:22]
  wire [7:0] n126_I_2_2; // @[Top.scala 25:22]
  wire [7:0] n126_O_0_0; // @[Top.scala 25:22]
  wire [7:0] n126_O_1_0; // @[Top.scala 25:22]
  wire [7:0] n126_O_2_0; // @[Top.scala 25:22]
  wire  n131_clock; // @[Top.scala 28:22]
  wire  n131_reset; // @[Top.scala 28:22]
  wire  n131_valid_up; // @[Top.scala 28:22]
  wire  n131_valid_down; // @[Top.scala 28:22]
  wire [7:0] n131_I_0_0; // @[Top.scala 28:22]
  wire [7:0] n131_I_1_0; // @[Top.scala 28:22]
  wire [7:0] n131_I_2_0; // @[Top.scala 28:22]
  wire [7:0] n131_O_0_0; // @[Top.scala 28:22]
  wire  InitialDelayCounter_1_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_valid_down; // @[Const.scala 11:33]
  wire  n134_valid_up; // @[Top.scala 32:22]
  wire  n134_valid_down; // @[Top.scala 32:22]
  wire [7:0] n134_I0_0_0; // @[Top.scala 32:22]
  wire [7:0] n134_O_0_0_t0b; // @[Top.scala 32:22]
  wire  n145_clock; // @[Top.scala 36:22]
  wire  n145_reset; // @[Top.scala 36:22]
  wire  n145_valid_up; // @[Top.scala 36:22]
  wire  n145_valid_down; // @[Top.scala 36:22]
  wire [7:0] n145_I_0_0_t0b; // @[Top.scala 36:22]
  wire [7:0] n145_O_0_0; // @[Top.scala 36:22]
  InitialDelayCounter InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  Map2S_9 n110 ( // @[Top.scala 18:22]
    .valid_up(n110_valid_up),
    .valid_down(n110_valid_down),
    .I0_0_0(n110_I0_0_0),
    .I0_0_1(n110_I0_0_1),
    .I0_0_2(n110_I0_0_2),
    .I0_1_0(n110_I0_1_0),
    .I0_1_1(n110_I0_1_1),
    .I0_1_2(n110_I0_1_2),
    .I0_2_0(n110_I0_2_0),
    .I0_2_1(n110_I0_2_1),
    .I0_2_2(n110_I0_2_2),
    .O_0_0_t0b(n110_O_0_0_t0b),
    .O_0_0_t1b(n110_O_0_0_t1b),
    .O_0_1_t0b(n110_O_0_1_t0b),
    .O_0_1_t1b(n110_O_0_1_t1b),
    .O_0_2_t0b(n110_O_0_2_t0b),
    .O_0_2_t1b(n110_O_0_2_t1b),
    .O_1_0_t0b(n110_O_1_0_t0b),
    .O_1_0_t1b(n110_O_1_0_t1b),
    .O_1_1_t0b(n110_O_1_1_t0b),
    .O_1_1_t1b(n110_O_1_1_t1b),
    .O_1_2_t0b(n110_O_1_2_t0b),
    .O_1_2_t1b(n110_O_1_2_t1b),
    .O_2_0_t0b(n110_O_2_0_t0b),
    .O_2_0_t1b(n110_O_2_0_t1b),
    .O_2_1_t0b(n110_O_2_1_t0b),
    .O_2_1_t1b(n110_O_2_1_t1b),
    .O_2_2_t0b(n110_O_2_2_t0b),
    .O_2_2_t1b(n110_O_2_2_t1b)
  );
  MapS_5 n121 ( // @[Top.scala 22:22]
    .clock(n121_clock),
    .reset(n121_reset),
    .valid_up(n121_valid_up),
    .valid_down(n121_valid_down),
    .I_0_0_t0b(n121_I_0_0_t0b),
    .I_0_0_t1b(n121_I_0_0_t1b),
    .I_0_1_t0b(n121_I_0_1_t0b),
    .I_0_1_t1b(n121_I_0_1_t1b),
    .I_0_2_t0b(n121_I_0_2_t0b),
    .I_0_2_t1b(n121_I_0_2_t1b),
    .I_1_0_t0b(n121_I_1_0_t0b),
    .I_1_0_t1b(n121_I_1_0_t1b),
    .I_1_1_t0b(n121_I_1_1_t0b),
    .I_1_1_t1b(n121_I_1_1_t1b),
    .I_1_2_t0b(n121_I_1_2_t0b),
    .I_1_2_t1b(n121_I_1_2_t1b),
    .I_2_0_t0b(n121_I_2_0_t0b),
    .I_2_0_t1b(n121_I_2_0_t1b),
    .I_2_1_t0b(n121_I_2_1_t0b),
    .I_2_1_t1b(n121_I_2_1_t1b),
    .I_2_2_t0b(n121_I_2_2_t0b),
    .I_2_2_t1b(n121_I_2_2_t1b),
    .O_0_0(n121_O_0_0),
    .O_0_1(n121_O_0_1),
    .O_0_2(n121_O_0_2),
    .O_1_0(n121_O_1_0),
    .O_1_1(n121_O_1_1),
    .O_1_2(n121_O_1_2),
    .O_2_0(n121_O_2_0),
    .O_2_1(n121_O_2_1),
    .O_2_2(n121_O_2_2)
  );
  MapS_6 n126 ( // @[Top.scala 25:22]
    .clock(n126_clock),
    .reset(n126_reset),
    .valid_up(n126_valid_up),
    .valid_down(n126_valid_down),
    .I_0_0(n126_I_0_0),
    .I_0_1(n126_I_0_1),
    .I_0_2(n126_I_0_2),
    .I_1_0(n126_I_1_0),
    .I_1_1(n126_I_1_1),
    .I_1_2(n126_I_1_2),
    .I_2_0(n126_I_2_0),
    .I_2_1(n126_I_2_1),
    .I_2_2(n126_I_2_2),
    .O_0_0(n126_O_0_0),
    .O_1_0(n126_O_1_0),
    .O_2_0(n126_O_2_0)
  );
  ReduceS_1 n131 ( // @[Top.scala 28:22]
    .clock(n131_clock),
    .reset(n131_reset),
    .valid_up(n131_valid_up),
    .valid_down(n131_valid_down),
    .I_0_0(n131_I_0_0),
    .I_1_0(n131_I_1_0),
    .I_2_0(n131_I_2_0),
    .O_0_0(n131_O_0_0)
  );
  InitialDelayCounter_1 InitialDelayCounter_1 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_1_clock),
    .reset(InitialDelayCounter_1_reset),
    .valid_down(InitialDelayCounter_1_valid_down)
  );
  Map2S_11 n134 ( // @[Top.scala 32:22]
    .valid_up(n134_valid_up),
    .valid_down(n134_valid_down),
    .I0_0_0(n134_I0_0_0),
    .O_0_0_t0b(n134_O_0_0_t0b)
  );
  MapS_8 n145 ( // @[Top.scala 36:22]
    .clock(n145_clock),
    .reset(n145_reset),
    .valid_up(n145_valid_up),
    .valid_down(n145_valid_down),
    .I_0_0_t0b(n145_I_0_0_t0b),
    .O_0_0(n145_O_0_0)
  );
  assign valid_down = n145_valid_down; // @[Top.scala 40:16]
  assign O_0_0 = n145_O_0_0; // @[Top.scala 39:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n110_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 21:19]
  assign n110_I0_0_0 = I_0_0; // @[Top.scala 19:13]
  assign n110_I0_0_1 = I_0_1; // @[Top.scala 19:13]
  assign n110_I0_0_2 = I_0_2; // @[Top.scala 19:13]
  assign n110_I0_1_0 = I_1_0; // @[Top.scala 19:13]
  assign n110_I0_1_1 = I_1_1; // @[Top.scala 19:13]
  assign n110_I0_1_2 = I_1_2; // @[Top.scala 19:13]
  assign n110_I0_2_0 = I_2_0; // @[Top.scala 19:13]
  assign n110_I0_2_1 = I_2_1; // @[Top.scala 19:13]
  assign n110_I0_2_2 = I_2_2; // @[Top.scala 19:13]
  assign n121_clock = clock;
  assign n121_reset = reset;
  assign n121_valid_up = n110_valid_down; // @[Top.scala 24:19]
  assign n121_I_0_0_t0b = n110_O_0_0_t0b; // @[Top.scala 23:12]
  assign n121_I_0_0_t1b = n110_O_0_0_t1b; // @[Top.scala 23:12]
  assign n121_I_0_1_t0b = n110_O_0_1_t0b; // @[Top.scala 23:12]
  assign n121_I_0_1_t1b = n110_O_0_1_t1b; // @[Top.scala 23:12]
  assign n121_I_0_2_t0b = n110_O_0_2_t0b; // @[Top.scala 23:12]
  assign n121_I_0_2_t1b = n110_O_0_2_t1b; // @[Top.scala 23:12]
  assign n121_I_1_0_t0b = n110_O_1_0_t0b; // @[Top.scala 23:12]
  assign n121_I_1_0_t1b = n110_O_1_0_t1b; // @[Top.scala 23:12]
  assign n121_I_1_1_t0b = n110_O_1_1_t0b; // @[Top.scala 23:12]
  assign n121_I_1_1_t1b = n110_O_1_1_t1b; // @[Top.scala 23:12]
  assign n121_I_1_2_t0b = n110_O_1_2_t0b; // @[Top.scala 23:12]
  assign n121_I_1_2_t1b = n110_O_1_2_t1b; // @[Top.scala 23:12]
  assign n121_I_2_0_t0b = n110_O_2_0_t0b; // @[Top.scala 23:12]
  assign n121_I_2_0_t1b = n110_O_2_0_t1b; // @[Top.scala 23:12]
  assign n121_I_2_1_t0b = n110_O_2_1_t0b; // @[Top.scala 23:12]
  assign n121_I_2_1_t1b = n110_O_2_1_t1b; // @[Top.scala 23:12]
  assign n121_I_2_2_t0b = n110_O_2_2_t0b; // @[Top.scala 23:12]
  assign n121_I_2_2_t1b = n110_O_2_2_t1b; // @[Top.scala 23:12]
  assign n126_clock = clock;
  assign n126_reset = reset;
  assign n126_valid_up = n121_valid_down; // @[Top.scala 27:19]
  assign n126_I_0_0 = n121_O_0_0; // @[Top.scala 26:12]
  assign n126_I_0_1 = n121_O_0_1; // @[Top.scala 26:12]
  assign n126_I_0_2 = n121_O_0_2; // @[Top.scala 26:12]
  assign n126_I_1_0 = n121_O_1_0; // @[Top.scala 26:12]
  assign n126_I_1_1 = n121_O_1_1; // @[Top.scala 26:12]
  assign n126_I_1_2 = n121_O_1_2; // @[Top.scala 26:12]
  assign n126_I_2_0 = n121_O_2_0; // @[Top.scala 26:12]
  assign n126_I_2_1 = n121_O_2_1; // @[Top.scala 26:12]
  assign n126_I_2_2 = n121_O_2_2; // @[Top.scala 26:12]
  assign n131_clock = clock;
  assign n131_reset = reset;
  assign n131_valid_up = n126_valid_down; // @[Top.scala 30:19]
  assign n131_I_0_0 = n126_O_0_0; // @[Top.scala 29:12]
  assign n131_I_1_0 = n126_O_1_0; // @[Top.scala 29:12]
  assign n131_I_2_0 = n126_O_2_0; // @[Top.scala 29:12]
  assign InitialDelayCounter_1_clock = clock;
  assign InitialDelayCounter_1_reset = reset;
  assign n134_valid_up = n131_valid_down & InitialDelayCounter_1_valid_down; // @[Top.scala 35:19]
  assign n134_I0_0_0 = n131_O_0_0; // @[Top.scala 33:13]
  assign n145_clock = clock;
  assign n145_reset = reset;
  assign n145_valid_up = n134_valid_down; // @[Top.scala 38:19]
  assign n145_I_0_0_t0b = n134_O_0_0_t0b; // @[Top.scala 37:12]
endmodule
module MapS_9(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  input  [7:0] I_1_1_0,
  input  [7:0] I_1_1_1,
  input  [7:0] I_1_1_2,
  input  [7:0] I_1_2_0,
  input  [7:0] I_1_2_1,
  input  [7:0] I_1_2_2,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  Module_0 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .I_1_0(fst_op_I_1_0),
    .I_1_1(fst_op_I_1_1),
    .I_1_2(fst_op_I_1_2),
    .I_2_0(fst_op_I_2_0),
    .I_2_1(fst_op_I_2_1),
    .I_2_2(fst_op_I_2_2),
    .O_0_0(fst_op_O_0_0)
  );
  Module_0 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .I_1_0(other_ops_0_I_1_0),
    .I_1_1(other_ops_0_I_1_1),
    .I_1_2(other_ops_0_I_1_2),
    .I_2_0(other_ops_0_I_2_0),
    .I_2_1(other_ops_0_I_2_1),
    .I_2_2(other_ops_0_I_2_2),
    .O_0_0(other_ops_0_O_0_0)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_1_0 = I_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_1_1 = I_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_1_2 = I_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_2_0 = I_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_2_1 = I_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_2_2 = I_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_0 = I_1_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_1 = I_1_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_2 = I_1_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_0 = I_1_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_1 = I_1_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_2 = I_1_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_8(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  input  [7:0] I_1_1_0,
  input  [7:0] I_1_1_1,
  input  [7:0] I_1_1_2,
  input  [7:0] I_1_2_0,
  input  [7:0] I_1_2_1,
  input  [7:0] I_1_2_2,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[MapT.scala 8:20]
  MapS_9 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_1_0_0(op_O_1_0_0)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
endmodule
module Passthrough(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_1_0_0,
  output [7:0] O_0_0,
  output [7:0] O_1_0
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0_0 = I_0_0_0; // @[Passthrough.scala 17:68]
  assign O_1_0 = I_1_0_0; // @[Passthrough.scala 17:68]
endmodule
module Passthrough_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_1_0,
  output [7:0] O_0,
  output [7:0] O_1
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0 = I_0_0; // @[Passthrough.scala 17:68]
  assign O_1 = I_1_0; // @[Passthrough.scala 17:68]
endmodule
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  output [7:0] O_0,
  output [7:0] O_1
);
  wire  n1_clock; // @[Top.scala 46:20]
  wire  n1_reset; // @[Top.scala 46:20]
  wire  n1_valid_up; // @[Top.scala 46:20]
  wire  n1_valid_down; // @[Top.scala 46:20]
  wire [7:0] n1_I_0; // @[Top.scala 46:20]
  wire [7:0] n1_I_1; // @[Top.scala 46:20]
  wire [7:0] n1_O_0; // @[Top.scala 46:20]
  wire [7:0] n1_O_1; // @[Top.scala 46:20]
  wire  n2_clock; // @[Top.scala 49:20]
  wire  n2_reset; // @[Top.scala 49:20]
  wire  n2_valid_up; // @[Top.scala 49:20]
  wire  n2_valid_down; // @[Top.scala 49:20]
  wire [7:0] n2_I_0; // @[Top.scala 49:20]
  wire [7:0] n2_I_1; // @[Top.scala 49:20]
  wire [7:0] n2_O_0; // @[Top.scala 49:20]
  wire [7:0] n2_O_1; // @[Top.scala 49:20]
  wire  n3_clock; // @[Top.scala 52:20]
  wire  n3_reset; // @[Top.scala 52:20]
  wire  n3_valid_up; // @[Top.scala 52:20]
  wire  n3_valid_down; // @[Top.scala 52:20]
  wire [7:0] n3_I_0; // @[Top.scala 52:20]
  wire [7:0] n3_I_1; // @[Top.scala 52:20]
  wire [7:0] n3_O_0; // @[Top.scala 52:20]
  wire [7:0] n3_O_1; // @[Top.scala 52:20]
  wire  n4_clock; // @[Top.scala 55:20]
  wire  n4_valid_up; // @[Top.scala 55:20]
  wire  n4_valid_down; // @[Top.scala 55:20]
  wire [7:0] n4_I_0; // @[Top.scala 55:20]
  wire [7:0] n4_I_1; // @[Top.scala 55:20]
  wire [7:0] n4_O_0; // @[Top.scala 55:20]
  wire [7:0] n4_O_1; // @[Top.scala 55:20]
  wire  n5_clock; // @[Top.scala 58:20]
  wire  n5_valid_up; // @[Top.scala 58:20]
  wire  n5_valid_down; // @[Top.scala 58:20]
  wire [7:0] n5_I_0; // @[Top.scala 58:20]
  wire [7:0] n5_I_1; // @[Top.scala 58:20]
  wire [7:0] n5_O_0; // @[Top.scala 58:20]
  wire [7:0] n5_O_1; // @[Top.scala 58:20]
  wire  n6_valid_up; // @[Top.scala 61:20]
  wire  n6_valid_down; // @[Top.scala 61:20]
  wire [7:0] n6_I0_0; // @[Top.scala 61:20]
  wire [7:0] n6_I0_1; // @[Top.scala 61:20]
  wire [7:0] n6_I1_0; // @[Top.scala 61:20]
  wire [7:0] n6_I1_1; // @[Top.scala 61:20]
  wire [7:0] n6_O_0_0; // @[Top.scala 61:20]
  wire [7:0] n6_O_0_1; // @[Top.scala 61:20]
  wire [7:0] n6_O_1_0; // @[Top.scala 61:20]
  wire [7:0] n6_O_1_1; // @[Top.scala 61:20]
  wire  n13_valid_up; // @[Top.scala 65:21]
  wire  n13_valid_down; // @[Top.scala 65:21]
  wire [7:0] n13_I0_0_0; // @[Top.scala 65:21]
  wire [7:0] n13_I0_0_1; // @[Top.scala 65:21]
  wire [7:0] n13_I0_1_0; // @[Top.scala 65:21]
  wire [7:0] n13_I0_1_1; // @[Top.scala 65:21]
  wire [7:0] n13_I1_0; // @[Top.scala 65:21]
  wire [7:0] n13_I1_1; // @[Top.scala 65:21]
  wire [7:0] n13_O_0_0; // @[Top.scala 65:21]
  wire [7:0] n13_O_0_1; // @[Top.scala 65:21]
  wire [7:0] n13_O_0_2; // @[Top.scala 65:21]
  wire [7:0] n13_O_1_0; // @[Top.scala 65:21]
  wire [7:0] n13_O_1_1; // @[Top.scala 65:21]
  wire [7:0] n13_O_1_2; // @[Top.scala 65:21]
  wire  n22_valid_up; // @[Top.scala 69:21]
  wire  n22_valid_down; // @[Top.scala 69:21]
  wire [7:0] n22_I_0_0; // @[Top.scala 69:21]
  wire [7:0] n22_I_0_1; // @[Top.scala 69:21]
  wire [7:0] n22_I_0_2; // @[Top.scala 69:21]
  wire [7:0] n22_I_1_0; // @[Top.scala 69:21]
  wire [7:0] n22_I_1_1; // @[Top.scala 69:21]
  wire [7:0] n22_I_1_2; // @[Top.scala 69:21]
  wire [7:0] n22_O_0_0_0; // @[Top.scala 69:21]
  wire [7:0] n22_O_0_0_1; // @[Top.scala 69:21]
  wire [7:0] n22_O_0_0_2; // @[Top.scala 69:21]
  wire [7:0] n22_O_1_0_0; // @[Top.scala 69:21]
  wire [7:0] n22_O_1_0_1; // @[Top.scala 69:21]
  wire [7:0] n22_O_1_0_2; // @[Top.scala 69:21]
  wire  n29_valid_up; // @[Top.scala 72:21]
  wire  n29_valid_down; // @[Top.scala 72:21]
  wire [7:0] n29_I_0_0_0; // @[Top.scala 72:21]
  wire [7:0] n29_I_0_0_1; // @[Top.scala 72:21]
  wire [7:0] n29_I_0_0_2; // @[Top.scala 72:21]
  wire [7:0] n29_I_1_0_0; // @[Top.scala 72:21]
  wire [7:0] n29_I_1_0_1; // @[Top.scala 72:21]
  wire [7:0] n29_I_1_0_2; // @[Top.scala 72:21]
  wire [7:0] n29_O_0_0; // @[Top.scala 72:21]
  wire [7:0] n29_O_0_1; // @[Top.scala 72:21]
  wire [7:0] n29_O_0_2; // @[Top.scala 72:21]
  wire [7:0] n29_O_1_0; // @[Top.scala 72:21]
  wire [7:0] n29_O_1_1; // @[Top.scala 72:21]
  wire [7:0] n29_O_1_2; // @[Top.scala 72:21]
  wire  n30_clock; // @[Top.scala 75:21]
  wire  n30_valid_up; // @[Top.scala 75:21]
  wire  n30_valid_down; // @[Top.scala 75:21]
  wire [7:0] n30_I_0; // @[Top.scala 75:21]
  wire [7:0] n30_I_1; // @[Top.scala 75:21]
  wire [7:0] n30_O_0; // @[Top.scala 75:21]
  wire [7:0] n30_O_1; // @[Top.scala 75:21]
  wire  n31_clock; // @[Top.scala 78:21]
  wire  n31_valid_up; // @[Top.scala 78:21]
  wire  n31_valid_down; // @[Top.scala 78:21]
  wire [7:0] n31_I_0; // @[Top.scala 78:21]
  wire [7:0] n31_I_1; // @[Top.scala 78:21]
  wire [7:0] n31_O_0; // @[Top.scala 78:21]
  wire [7:0] n31_O_1; // @[Top.scala 78:21]
  wire  n32_valid_up; // @[Top.scala 81:21]
  wire  n32_valid_down; // @[Top.scala 81:21]
  wire [7:0] n32_I0_0; // @[Top.scala 81:21]
  wire [7:0] n32_I0_1; // @[Top.scala 81:21]
  wire [7:0] n32_I1_0; // @[Top.scala 81:21]
  wire [7:0] n32_I1_1; // @[Top.scala 81:21]
  wire [7:0] n32_O_0_0; // @[Top.scala 81:21]
  wire [7:0] n32_O_0_1; // @[Top.scala 81:21]
  wire [7:0] n32_O_1_0; // @[Top.scala 81:21]
  wire [7:0] n32_O_1_1; // @[Top.scala 81:21]
  wire  n39_valid_up; // @[Top.scala 85:21]
  wire  n39_valid_down; // @[Top.scala 85:21]
  wire [7:0] n39_I0_0_0; // @[Top.scala 85:21]
  wire [7:0] n39_I0_0_1; // @[Top.scala 85:21]
  wire [7:0] n39_I0_1_0; // @[Top.scala 85:21]
  wire [7:0] n39_I0_1_1; // @[Top.scala 85:21]
  wire [7:0] n39_I1_0; // @[Top.scala 85:21]
  wire [7:0] n39_I1_1; // @[Top.scala 85:21]
  wire [7:0] n39_O_0_0; // @[Top.scala 85:21]
  wire [7:0] n39_O_0_1; // @[Top.scala 85:21]
  wire [7:0] n39_O_0_2; // @[Top.scala 85:21]
  wire [7:0] n39_O_1_0; // @[Top.scala 85:21]
  wire [7:0] n39_O_1_1; // @[Top.scala 85:21]
  wire [7:0] n39_O_1_2; // @[Top.scala 85:21]
  wire  n48_valid_up; // @[Top.scala 89:21]
  wire  n48_valid_down; // @[Top.scala 89:21]
  wire [7:0] n48_I_0_0; // @[Top.scala 89:21]
  wire [7:0] n48_I_0_1; // @[Top.scala 89:21]
  wire [7:0] n48_I_0_2; // @[Top.scala 89:21]
  wire [7:0] n48_I_1_0; // @[Top.scala 89:21]
  wire [7:0] n48_I_1_1; // @[Top.scala 89:21]
  wire [7:0] n48_I_1_2; // @[Top.scala 89:21]
  wire [7:0] n48_O_0_0_0; // @[Top.scala 89:21]
  wire [7:0] n48_O_0_0_1; // @[Top.scala 89:21]
  wire [7:0] n48_O_0_0_2; // @[Top.scala 89:21]
  wire [7:0] n48_O_1_0_0; // @[Top.scala 89:21]
  wire [7:0] n48_O_1_0_1; // @[Top.scala 89:21]
  wire [7:0] n48_O_1_0_2; // @[Top.scala 89:21]
  wire  n55_valid_up; // @[Top.scala 92:21]
  wire  n55_valid_down; // @[Top.scala 92:21]
  wire [7:0] n55_I_0_0_0; // @[Top.scala 92:21]
  wire [7:0] n55_I_0_0_1; // @[Top.scala 92:21]
  wire [7:0] n55_I_0_0_2; // @[Top.scala 92:21]
  wire [7:0] n55_I_1_0_0; // @[Top.scala 92:21]
  wire [7:0] n55_I_1_0_1; // @[Top.scala 92:21]
  wire [7:0] n55_I_1_0_2; // @[Top.scala 92:21]
  wire [7:0] n55_O_0_0; // @[Top.scala 92:21]
  wire [7:0] n55_O_0_1; // @[Top.scala 92:21]
  wire [7:0] n55_O_0_2; // @[Top.scala 92:21]
  wire [7:0] n55_O_1_0; // @[Top.scala 92:21]
  wire [7:0] n55_O_1_1; // @[Top.scala 92:21]
  wire [7:0] n55_O_1_2; // @[Top.scala 92:21]
  wire  n56_valid_up; // @[Top.scala 95:21]
  wire  n56_valid_down; // @[Top.scala 95:21]
  wire [7:0] n56_I0_0_0; // @[Top.scala 95:21]
  wire [7:0] n56_I0_0_1; // @[Top.scala 95:21]
  wire [7:0] n56_I0_0_2; // @[Top.scala 95:21]
  wire [7:0] n56_I0_1_0; // @[Top.scala 95:21]
  wire [7:0] n56_I0_1_1; // @[Top.scala 95:21]
  wire [7:0] n56_I0_1_2; // @[Top.scala 95:21]
  wire [7:0] n56_I1_0_0; // @[Top.scala 95:21]
  wire [7:0] n56_I1_0_1; // @[Top.scala 95:21]
  wire [7:0] n56_I1_0_2; // @[Top.scala 95:21]
  wire [7:0] n56_I1_1_0; // @[Top.scala 95:21]
  wire [7:0] n56_I1_1_1; // @[Top.scala 95:21]
  wire [7:0] n56_I1_1_2; // @[Top.scala 95:21]
  wire [7:0] n56_O_0_0_0; // @[Top.scala 95:21]
  wire [7:0] n56_O_0_0_1; // @[Top.scala 95:21]
  wire [7:0] n56_O_0_0_2; // @[Top.scala 95:21]
  wire [7:0] n56_O_0_1_0; // @[Top.scala 95:21]
  wire [7:0] n56_O_0_1_1; // @[Top.scala 95:21]
  wire [7:0] n56_O_0_1_2; // @[Top.scala 95:21]
  wire [7:0] n56_O_1_0_0; // @[Top.scala 95:21]
  wire [7:0] n56_O_1_0_1; // @[Top.scala 95:21]
  wire [7:0] n56_O_1_0_2; // @[Top.scala 95:21]
  wire [7:0] n56_O_1_1_0; // @[Top.scala 95:21]
  wire [7:0] n56_O_1_1_1; // @[Top.scala 95:21]
  wire [7:0] n56_O_1_1_2; // @[Top.scala 95:21]
  wire  n63_clock; // @[Top.scala 99:21]
  wire  n63_valid_up; // @[Top.scala 99:21]
  wire  n63_valid_down; // @[Top.scala 99:21]
  wire [7:0] n63_I_0; // @[Top.scala 99:21]
  wire [7:0] n63_I_1; // @[Top.scala 99:21]
  wire [7:0] n63_O_0; // @[Top.scala 99:21]
  wire [7:0] n63_O_1; // @[Top.scala 99:21]
  wire  n64_clock; // @[Top.scala 102:21]
  wire  n64_valid_up; // @[Top.scala 102:21]
  wire  n64_valid_down; // @[Top.scala 102:21]
  wire [7:0] n64_I_0; // @[Top.scala 102:21]
  wire [7:0] n64_I_1; // @[Top.scala 102:21]
  wire [7:0] n64_O_0; // @[Top.scala 102:21]
  wire [7:0] n64_O_1; // @[Top.scala 102:21]
  wire  n65_valid_up; // @[Top.scala 105:21]
  wire  n65_valid_down; // @[Top.scala 105:21]
  wire [7:0] n65_I0_0; // @[Top.scala 105:21]
  wire [7:0] n65_I0_1; // @[Top.scala 105:21]
  wire [7:0] n65_I1_0; // @[Top.scala 105:21]
  wire [7:0] n65_I1_1; // @[Top.scala 105:21]
  wire [7:0] n65_O_0_0; // @[Top.scala 105:21]
  wire [7:0] n65_O_0_1; // @[Top.scala 105:21]
  wire [7:0] n65_O_1_0; // @[Top.scala 105:21]
  wire [7:0] n65_O_1_1; // @[Top.scala 105:21]
  wire  n72_valid_up; // @[Top.scala 109:21]
  wire  n72_valid_down; // @[Top.scala 109:21]
  wire [7:0] n72_I0_0_0; // @[Top.scala 109:21]
  wire [7:0] n72_I0_0_1; // @[Top.scala 109:21]
  wire [7:0] n72_I0_1_0; // @[Top.scala 109:21]
  wire [7:0] n72_I0_1_1; // @[Top.scala 109:21]
  wire [7:0] n72_I1_0; // @[Top.scala 109:21]
  wire [7:0] n72_I1_1; // @[Top.scala 109:21]
  wire [7:0] n72_O_0_0; // @[Top.scala 109:21]
  wire [7:0] n72_O_0_1; // @[Top.scala 109:21]
  wire [7:0] n72_O_0_2; // @[Top.scala 109:21]
  wire [7:0] n72_O_1_0; // @[Top.scala 109:21]
  wire [7:0] n72_O_1_1; // @[Top.scala 109:21]
  wire [7:0] n72_O_1_2; // @[Top.scala 109:21]
  wire  n81_valid_up; // @[Top.scala 113:21]
  wire  n81_valid_down; // @[Top.scala 113:21]
  wire [7:0] n81_I_0_0; // @[Top.scala 113:21]
  wire [7:0] n81_I_0_1; // @[Top.scala 113:21]
  wire [7:0] n81_I_0_2; // @[Top.scala 113:21]
  wire [7:0] n81_I_1_0; // @[Top.scala 113:21]
  wire [7:0] n81_I_1_1; // @[Top.scala 113:21]
  wire [7:0] n81_I_1_2; // @[Top.scala 113:21]
  wire [7:0] n81_O_0_0_0; // @[Top.scala 113:21]
  wire [7:0] n81_O_0_0_1; // @[Top.scala 113:21]
  wire [7:0] n81_O_0_0_2; // @[Top.scala 113:21]
  wire [7:0] n81_O_1_0_0; // @[Top.scala 113:21]
  wire [7:0] n81_O_1_0_1; // @[Top.scala 113:21]
  wire [7:0] n81_O_1_0_2; // @[Top.scala 113:21]
  wire  n88_valid_up; // @[Top.scala 116:21]
  wire  n88_valid_down; // @[Top.scala 116:21]
  wire [7:0] n88_I_0_0_0; // @[Top.scala 116:21]
  wire [7:0] n88_I_0_0_1; // @[Top.scala 116:21]
  wire [7:0] n88_I_0_0_2; // @[Top.scala 116:21]
  wire [7:0] n88_I_1_0_0; // @[Top.scala 116:21]
  wire [7:0] n88_I_1_0_1; // @[Top.scala 116:21]
  wire [7:0] n88_I_1_0_2; // @[Top.scala 116:21]
  wire [7:0] n88_O_0_0; // @[Top.scala 116:21]
  wire [7:0] n88_O_0_1; // @[Top.scala 116:21]
  wire [7:0] n88_O_0_2; // @[Top.scala 116:21]
  wire [7:0] n88_O_1_0; // @[Top.scala 116:21]
  wire [7:0] n88_O_1_1; // @[Top.scala 116:21]
  wire [7:0] n88_O_1_2; // @[Top.scala 116:21]
  wire  n89_valid_up; // @[Top.scala 119:21]
  wire  n89_valid_down; // @[Top.scala 119:21]
  wire [7:0] n89_I0_0_0_0; // @[Top.scala 119:21]
  wire [7:0] n89_I0_0_0_1; // @[Top.scala 119:21]
  wire [7:0] n89_I0_0_0_2; // @[Top.scala 119:21]
  wire [7:0] n89_I0_0_1_0; // @[Top.scala 119:21]
  wire [7:0] n89_I0_0_1_1; // @[Top.scala 119:21]
  wire [7:0] n89_I0_0_1_2; // @[Top.scala 119:21]
  wire [7:0] n89_I0_1_0_0; // @[Top.scala 119:21]
  wire [7:0] n89_I0_1_0_1; // @[Top.scala 119:21]
  wire [7:0] n89_I0_1_0_2; // @[Top.scala 119:21]
  wire [7:0] n89_I0_1_1_0; // @[Top.scala 119:21]
  wire [7:0] n89_I0_1_1_1; // @[Top.scala 119:21]
  wire [7:0] n89_I0_1_1_2; // @[Top.scala 119:21]
  wire [7:0] n89_I1_0_0; // @[Top.scala 119:21]
  wire [7:0] n89_I1_0_1; // @[Top.scala 119:21]
  wire [7:0] n89_I1_0_2; // @[Top.scala 119:21]
  wire [7:0] n89_I1_1_0; // @[Top.scala 119:21]
  wire [7:0] n89_I1_1_1; // @[Top.scala 119:21]
  wire [7:0] n89_I1_1_2; // @[Top.scala 119:21]
  wire [7:0] n89_O_0_0_0; // @[Top.scala 119:21]
  wire [7:0] n89_O_0_0_1; // @[Top.scala 119:21]
  wire [7:0] n89_O_0_0_2; // @[Top.scala 119:21]
  wire [7:0] n89_O_0_1_0; // @[Top.scala 119:21]
  wire [7:0] n89_O_0_1_1; // @[Top.scala 119:21]
  wire [7:0] n89_O_0_1_2; // @[Top.scala 119:21]
  wire [7:0] n89_O_0_2_0; // @[Top.scala 119:21]
  wire [7:0] n89_O_0_2_1; // @[Top.scala 119:21]
  wire [7:0] n89_O_0_2_2; // @[Top.scala 119:21]
  wire [7:0] n89_O_1_0_0; // @[Top.scala 119:21]
  wire [7:0] n89_O_1_0_1; // @[Top.scala 119:21]
  wire [7:0] n89_O_1_0_2; // @[Top.scala 119:21]
  wire [7:0] n89_O_1_1_0; // @[Top.scala 119:21]
  wire [7:0] n89_O_1_1_1; // @[Top.scala 119:21]
  wire [7:0] n89_O_1_1_2; // @[Top.scala 119:21]
  wire [7:0] n89_O_1_2_0; // @[Top.scala 119:21]
  wire [7:0] n89_O_1_2_1; // @[Top.scala 119:21]
  wire [7:0] n89_O_1_2_2; // @[Top.scala 119:21]
  wire  n98_valid_up; // @[Top.scala 123:21]
  wire  n98_valid_down; // @[Top.scala 123:21]
  wire [7:0] n98_I_0_0_0; // @[Top.scala 123:21]
  wire [7:0] n98_I_0_0_1; // @[Top.scala 123:21]
  wire [7:0] n98_I_0_0_2; // @[Top.scala 123:21]
  wire [7:0] n98_I_0_1_0; // @[Top.scala 123:21]
  wire [7:0] n98_I_0_1_1; // @[Top.scala 123:21]
  wire [7:0] n98_I_0_1_2; // @[Top.scala 123:21]
  wire [7:0] n98_I_0_2_0; // @[Top.scala 123:21]
  wire [7:0] n98_I_0_2_1; // @[Top.scala 123:21]
  wire [7:0] n98_I_0_2_2; // @[Top.scala 123:21]
  wire [7:0] n98_I_1_0_0; // @[Top.scala 123:21]
  wire [7:0] n98_I_1_0_1; // @[Top.scala 123:21]
  wire [7:0] n98_I_1_0_2; // @[Top.scala 123:21]
  wire [7:0] n98_I_1_1_0; // @[Top.scala 123:21]
  wire [7:0] n98_I_1_1_1; // @[Top.scala 123:21]
  wire [7:0] n98_I_1_1_2; // @[Top.scala 123:21]
  wire [7:0] n98_I_1_2_0; // @[Top.scala 123:21]
  wire [7:0] n98_I_1_2_1; // @[Top.scala 123:21]
  wire [7:0] n98_I_1_2_2; // @[Top.scala 123:21]
  wire [7:0] n98_O_0_0_0_0; // @[Top.scala 123:21]
  wire [7:0] n98_O_0_0_0_1; // @[Top.scala 123:21]
  wire [7:0] n98_O_0_0_0_2; // @[Top.scala 123:21]
  wire [7:0] n98_O_0_0_1_0; // @[Top.scala 123:21]
  wire [7:0] n98_O_0_0_1_1; // @[Top.scala 123:21]
  wire [7:0] n98_O_0_0_1_2; // @[Top.scala 123:21]
  wire [7:0] n98_O_0_0_2_0; // @[Top.scala 123:21]
  wire [7:0] n98_O_0_0_2_1; // @[Top.scala 123:21]
  wire [7:0] n98_O_0_0_2_2; // @[Top.scala 123:21]
  wire [7:0] n98_O_1_0_0_0; // @[Top.scala 123:21]
  wire [7:0] n98_O_1_0_0_1; // @[Top.scala 123:21]
  wire [7:0] n98_O_1_0_0_2; // @[Top.scala 123:21]
  wire [7:0] n98_O_1_0_1_0; // @[Top.scala 123:21]
  wire [7:0] n98_O_1_0_1_1; // @[Top.scala 123:21]
  wire [7:0] n98_O_1_0_1_2; // @[Top.scala 123:21]
  wire [7:0] n98_O_1_0_2_0; // @[Top.scala 123:21]
  wire [7:0] n98_O_1_0_2_1; // @[Top.scala 123:21]
  wire [7:0] n98_O_1_0_2_2; // @[Top.scala 123:21]
  wire  n105_valid_up; // @[Top.scala 126:22]
  wire  n105_valid_down; // @[Top.scala 126:22]
  wire [7:0] n105_I_0_0_0_0; // @[Top.scala 126:22]
  wire [7:0] n105_I_0_0_0_1; // @[Top.scala 126:22]
  wire [7:0] n105_I_0_0_0_2; // @[Top.scala 126:22]
  wire [7:0] n105_I_0_0_1_0; // @[Top.scala 126:22]
  wire [7:0] n105_I_0_0_1_1; // @[Top.scala 126:22]
  wire [7:0] n105_I_0_0_1_2; // @[Top.scala 126:22]
  wire [7:0] n105_I_0_0_2_0; // @[Top.scala 126:22]
  wire [7:0] n105_I_0_0_2_1; // @[Top.scala 126:22]
  wire [7:0] n105_I_0_0_2_2; // @[Top.scala 126:22]
  wire [7:0] n105_I_1_0_0_0; // @[Top.scala 126:22]
  wire [7:0] n105_I_1_0_0_1; // @[Top.scala 126:22]
  wire [7:0] n105_I_1_0_0_2; // @[Top.scala 126:22]
  wire [7:0] n105_I_1_0_1_0; // @[Top.scala 126:22]
  wire [7:0] n105_I_1_0_1_1; // @[Top.scala 126:22]
  wire [7:0] n105_I_1_0_1_2; // @[Top.scala 126:22]
  wire [7:0] n105_I_1_0_2_0; // @[Top.scala 126:22]
  wire [7:0] n105_I_1_0_2_1; // @[Top.scala 126:22]
  wire [7:0] n105_I_1_0_2_2; // @[Top.scala 126:22]
  wire [7:0] n105_O_0_0_0; // @[Top.scala 126:22]
  wire [7:0] n105_O_0_0_1; // @[Top.scala 126:22]
  wire [7:0] n105_O_0_0_2; // @[Top.scala 126:22]
  wire [7:0] n105_O_0_1_0; // @[Top.scala 126:22]
  wire [7:0] n105_O_0_1_1; // @[Top.scala 126:22]
  wire [7:0] n105_O_0_1_2; // @[Top.scala 126:22]
  wire [7:0] n105_O_0_2_0; // @[Top.scala 126:22]
  wire [7:0] n105_O_0_2_1; // @[Top.scala 126:22]
  wire [7:0] n105_O_0_2_2; // @[Top.scala 126:22]
  wire [7:0] n105_O_1_0_0; // @[Top.scala 126:22]
  wire [7:0] n105_O_1_0_1; // @[Top.scala 126:22]
  wire [7:0] n105_O_1_0_2; // @[Top.scala 126:22]
  wire [7:0] n105_O_1_1_0; // @[Top.scala 126:22]
  wire [7:0] n105_O_1_1_1; // @[Top.scala 126:22]
  wire [7:0] n105_O_1_1_2; // @[Top.scala 126:22]
  wire [7:0] n105_O_1_2_0; // @[Top.scala 126:22]
  wire [7:0] n105_O_1_2_1; // @[Top.scala 126:22]
  wire [7:0] n105_O_1_2_2; // @[Top.scala 126:22]
  wire  n147_clock; // @[Top.scala 129:22]
  wire  n147_reset; // @[Top.scala 129:22]
  wire  n147_valid_up; // @[Top.scala 129:22]
  wire  n147_valid_down; // @[Top.scala 129:22]
  wire [7:0] n147_I_0_0_0; // @[Top.scala 129:22]
  wire [7:0] n147_I_0_0_1; // @[Top.scala 129:22]
  wire [7:0] n147_I_0_0_2; // @[Top.scala 129:22]
  wire [7:0] n147_I_0_1_0; // @[Top.scala 129:22]
  wire [7:0] n147_I_0_1_1; // @[Top.scala 129:22]
  wire [7:0] n147_I_0_1_2; // @[Top.scala 129:22]
  wire [7:0] n147_I_0_2_0; // @[Top.scala 129:22]
  wire [7:0] n147_I_0_2_1; // @[Top.scala 129:22]
  wire [7:0] n147_I_0_2_2; // @[Top.scala 129:22]
  wire [7:0] n147_I_1_0_0; // @[Top.scala 129:22]
  wire [7:0] n147_I_1_0_1; // @[Top.scala 129:22]
  wire [7:0] n147_I_1_0_2; // @[Top.scala 129:22]
  wire [7:0] n147_I_1_1_0; // @[Top.scala 129:22]
  wire [7:0] n147_I_1_1_1; // @[Top.scala 129:22]
  wire [7:0] n147_I_1_1_2; // @[Top.scala 129:22]
  wire [7:0] n147_I_1_2_0; // @[Top.scala 129:22]
  wire [7:0] n147_I_1_2_1; // @[Top.scala 129:22]
  wire [7:0] n147_I_1_2_2; // @[Top.scala 129:22]
  wire [7:0] n147_O_0_0_0; // @[Top.scala 129:22]
  wire [7:0] n147_O_1_0_0; // @[Top.scala 129:22]
  wire  n148_valid_up; // @[Top.scala 132:22]
  wire  n148_valid_down; // @[Top.scala 132:22]
  wire [7:0] n148_I_0_0_0; // @[Top.scala 132:22]
  wire [7:0] n148_I_1_0_0; // @[Top.scala 132:22]
  wire [7:0] n148_O_0_0; // @[Top.scala 132:22]
  wire [7:0] n148_O_1_0; // @[Top.scala 132:22]
  wire  n149_valid_up; // @[Top.scala 135:22]
  wire  n149_valid_down; // @[Top.scala 135:22]
  wire [7:0] n149_I_0_0; // @[Top.scala 135:22]
  wire [7:0] n149_I_1_0; // @[Top.scala 135:22]
  wire [7:0] n149_O_0; // @[Top.scala 135:22]
  wire [7:0] n149_O_1; // @[Top.scala 135:22]
  wire  n150_clock; // @[Top.scala 138:22]
  wire  n150_reset; // @[Top.scala 138:22]
  wire  n150_valid_up; // @[Top.scala 138:22]
  wire  n150_valid_down; // @[Top.scala 138:22]
  wire [7:0] n150_I_0; // @[Top.scala 138:22]
  wire [7:0] n150_I_1; // @[Top.scala 138:22]
  wire [7:0] n150_O_0; // @[Top.scala 138:22]
  wire [7:0] n150_O_1; // @[Top.scala 138:22]
  wire  n151_clock; // @[Top.scala 141:22]
  wire  n151_reset; // @[Top.scala 141:22]
  wire  n151_valid_up; // @[Top.scala 141:22]
  wire  n151_valid_down; // @[Top.scala 141:22]
  wire [7:0] n151_I_0; // @[Top.scala 141:22]
  wire [7:0] n151_I_1; // @[Top.scala 141:22]
  wire [7:0] n151_O_0; // @[Top.scala 141:22]
  wire [7:0] n151_O_1; // @[Top.scala 141:22]
  wire  n152_clock; // @[Top.scala 144:22]
  wire  n152_reset; // @[Top.scala 144:22]
  wire  n152_valid_up; // @[Top.scala 144:22]
  wire  n152_valid_down; // @[Top.scala 144:22]
  wire [7:0] n152_I_0; // @[Top.scala 144:22]
  wire [7:0] n152_I_1; // @[Top.scala 144:22]
  wire [7:0] n152_O_0; // @[Top.scala 144:22]
  wire [7:0] n152_O_1; // @[Top.scala 144:22]
  FIFO n1 ( // @[Top.scala 46:20]
    .clock(n1_clock),
    .reset(n1_reset),
    .valid_up(n1_valid_up),
    .valid_down(n1_valid_down),
    .I_0(n1_I_0),
    .I_1(n1_I_1),
    .O_0(n1_O_0),
    .O_1(n1_O_1)
  );
  ShiftTS n2 ( // @[Top.scala 49:20]
    .clock(n2_clock),
    .reset(n2_reset),
    .valid_up(n2_valid_up),
    .valid_down(n2_valid_down),
    .I_0(n2_I_0),
    .I_1(n2_I_1),
    .O_0(n2_O_0),
    .O_1(n2_O_1)
  );
  ShiftTS n3 ( // @[Top.scala 52:20]
    .clock(n3_clock),
    .reset(n3_reset),
    .valid_up(n3_valid_up),
    .valid_down(n3_valid_down),
    .I_0(n3_I_0),
    .I_1(n3_I_1),
    .O_0(n3_O_0),
    .O_1(n3_O_1)
  );
  ShiftTS_2 n4 ( // @[Top.scala 55:20]
    .clock(n4_clock),
    .valid_up(n4_valid_up),
    .valid_down(n4_valid_down),
    .I_0(n4_I_0),
    .I_1(n4_I_1),
    .O_0(n4_O_0),
    .O_1(n4_O_1)
  );
  ShiftTS_2 n5 ( // @[Top.scala 58:20]
    .clock(n5_clock),
    .valid_up(n5_valid_up),
    .valid_down(n5_valid_down),
    .I_0(n5_I_0),
    .I_1(n5_I_1),
    .O_0(n5_O_0),
    .O_1(n5_O_1)
  );
  Map2T n6 ( // @[Top.scala 61:20]
    .valid_up(n6_valid_up),
    .valid_down(n6_valid_down),
    .I0_0(n6_I0_0),
    .I0_1(n6_I0_1),
    .I1_0(n6_I1_0),
    .I1_1(n6_I1_1),
    .O_0_0(n6_O_0_0),
    .O_0_1(n6_O_0_1),
    .O_1_0(n6_O_1_0),
    .O_1_1(n6_O_1_1)
  );
  Map2T_1 n13 ( // @[Top.scala 65:21]
    .valid_up(n13_valid_up),
    .valid_down(n13_valid_down),
    .I0_0_0(n13_I0_0_0),
    .I0_0_1(n13_I0_0_1),
    .I0_1_0(n13_I0_1_0),
    .I0_1_1(n13_I0_1_1),
    .I1_0(n13_I1_0),
    .I1_1(n13_I1_1),
    .O_0_0(n13_O_0_0),
    .O_0_1(n13_O_0_1),
    .O_0_2(n13_O_0_2),
    .O_1_0(n13_O_1_0),
    .O_1_1(n13_O_1_1),
    .O_1_2(n13_O_1_2)
  );
  MapT n22 ( // @[Top.scala 69:21]
    .valid_up(n22_valid_up),
    .valid_down(n22_valid_down),
    .I_0_0(n22_I_0_0),
    .I_0_1(n22_I_0_1),
    .I_0_2(n22_I_0_2),
    .I_1_0(n22_I_1_0),
    .I_1_1(n22_I_1_1),
    .I_1_2(n22_I_1_2),
    .O_0_0_0(n22_O_0_0_0),
    .O_0_0_1(n22_O_0_0_1),
    .O_0_0_2(n22_O_0_0_2),
    .O_1_0_0(n22_O_1_0_0),
    .O_1_0_1(n22_O_1_0_1),
    .O_1_0_2(n22_O_1_0_2)
  );
  MapT_1 n29 ( // @[Top.scala 72:21]
    .valid_up(n29_valid_up),
    .valid_down(n29_valid_down),
    .I_0_0_0(n29_I_0_0_0),
    .I_0_0_1(n29_I_0_0_1),
    .I_0_0_2(n29_I_0_0_2),
    .I_1_0_0(n29_I_1_0_0),
    .I_1_0_1(n29_I_1_0_1),
    .I_1_0_2(n29_I_1_0_2),
    .O_0_0(n29_O_0_0),
    .O_0_1(n29_O_0_1),
    .O_0_2(n29_O_0_2),
    .O_1_0(n29_O_1_0),
    .O_1_1(n29_O_1_1),
    .O_1_2(n29_O_1_2)
  );
  ShiftTS_2 n30 ( // @[Top.scala 75:21]
    .clock(n30_clock),
    .valid_up(n30_valid_up),
    .valid_down(n30_valid_down),
    .I_0(n30_I_0),
    .I_1(n30_I_1),
    .O_0(n30_O_0),
    .O_1(n30_O_1)
  );
  ShiftTS_2 n31 ( // @[Top.scala 78:21]
    .clock(n31_clock),
    .valid_up(n31_valid_up),
    .valid_down(n31_valid_down),
    .I_0(n31_I_0),
    .I_1(n31_I_1),
    .O_0(n31_O_0),
    .O_1(n31_O_1)
  );
  Map2T n32 ( // @[Top.scala 81:21]
    .valid_up(n32_valid_up),
    .valid_down(n32_valid_down),
    .I0_0(n32_I0_0),
    .I0_1(n32_I0_1),
    .I1_0(n32_I1_0),
    .I1_1(n32_I1_1),
    .O_0_0(n32_O_0_0),
    .O_0_1(n32_O_0_1),
    .O_1_0(n32_O_1_0),
    .O_1_1(n32_O_1_1)
  );
  Map2T_1 n39 ( // @[Top.scala 85:21]
    .valid_up(n39_valid_up),
    .valid_down(n39_valid_down),
    .I0_0_0(n39_I0_0_0),
    .I0_0_1(n39_I0_0_1),
    .I0_1_0(n39_I0_1_0),
    .I0_1_1(n39_I0_1_1),
    .I1_0(n39_I1_0),
    .I1_1(n39_I1_1),
    .O_0_0(n39_O_0_0),
    .O_0_1(n39_O_0_1),
    .O_0_2(n39_O_0_2),
    .O_1_0(n39_O_1_0),
    .O_1_1(n39_O_1_1),
    .O_1_2(n39_O_1_2)
  );
  MapT n48 ( // @[Top.scala 89:21]
    .valid_up(n48_valid_up),
    .valid_down(n48_valid_down),
    .I_0_0(n48_I_0_0),
    .I_0_1(n48_I_0_1),
    .I_0_2(n48_I_0_2),
    .I_1_0(n48_I_1_0),
    .I_1_1(n48_I_1_1),
    .I_1_2(n48_I_1_2),
    .O_0_0_0(n48_O_0_0_0),
    .O_0_0_1(n48_O_0_0_1),
    .O_0_0_2(n48_O_0_0_2),
    .O_1_0_0(n48_O_1_0_0),
    .O_1_0_1(n48_O_1_0_1),
    .O_1_0_2(n48_O_1_0_2)
  );
  MapT_1 n55 ( // @[Top.scala 92:21]
    .valid_up(n55_valid_up),
    .valid_down(n55_valid_down),
    .I_0_0_0(n55_I_0_0_0),
    .I_0_0_1(n55_I_0_0_1),
    .I_0_0_2(n55_I_0_0_2),
    .I_1_0_0(n55_I_1_0_0),
    .I_1_0_1(n55_I_1_0_1),
    .I_1_0_2(n55_I_1_0_2),
    .O_0_0(n55_O_0_0),
    .O_0_1(n55_O_0_1),
    .O_0_2(n55_O_0_2),
    .O_1_0(n55_O_1_0),
    .O_1_1(n55_O_1_1),
    .O_1_2(n55_O_1_2)
  );
  Map2T_4 n56 ( // @[Top.scala 95:21]
    .valid_up(n56_valid_up),
    .valid_down(n56_valid_down),
    .I0_0_0(n56_I0_0_0),
    .I0_0_1(n56_I0_0_1),
    .I0_0_2(n56_I0_0_2),
    .I0_1_0(n56_I0_1_0),
    .I0_1_1(n56_I0_1_1),
    .I0_1_2(n56_I0_1_2),
    .I1_0_0(n56_I1_0_0),
    .I1_0_1(n56_I1_0_1),
    .I1_0_2(n56_I1_0_2),
    .I1_1_0(n56_I1_1_0),
    .I1_1_1(n56_I1_1_1),
    .I1_1_2(n56_I1_1_2),
    .O_0_0_0(n56_O_0_0_0),
    .O_0_0_1(n56_O_0_0_1),
    .O_0_0_2(n56_O_0_0_2),
    .O_0_1_0(n56_O_0_1_0),
    .O_0_1_1(n56_O_0_1_1),
    .O_0_1_2(n56_O_0_1_2),
    .O_1_0_0(n56_O_1_0_0),
    .O_1_0_1(n56_O_1_0_1),
    .O_1_0_2(n56_O_1_0_2),
    .O_1_1_0(n56_O_1_1_0),
    .O_1_1_1(n56_O_1_1_1),
    .O_1_1_2(n56_O_1_1_2)
  );
  ShiftTS_2 n63 ( // @[Top.scala 99:21]
    .clock(n63_clock),
    .valid_up(n63_valid_up),
    .valid_down(n63_valid_down),
    .I_0(n63_I_0),
    .I_1(n63_I_1),
    .O_0(n63_O_0),
    .O_1(n63_O_1)
  );
  ShiftTS_2 n64 ( // @[Top.scala 102:21]
    .clock(n64_clock),
    .valid_up(n64_valid_up),
    .valid_down(n64_valid_down),
    .I_0(n64_I_0),
    .I_1(n64_I_1),
    .O_0(n64_O_0),
    .O_1(n64_O_1)
  );
  Map2T n65 ( // @[Top.scala 105:21]
    .valid_up(n65_valid_up),
    .valid_down(n65_valid_down),
    .I0_0(n65_I0_0),
    .I0_1(n65_I0_1),
    .I1_0(n65_I1_0),
    .I1_1(n65_I1_1),
    .O_0_0(n65_O_0_0),
    .O_0_1(n65_O_0_1),
    .O_1_0(n65_O_1_0),
    .O_1_1(n65_O_1_1)
  );
  Map2T_1 n72 ( // @[Top.scala 109:21]
    .valid_up(n72_valid_up),
    .valid_down(n72_valid_down),
    .I0_0_0(n72_I0_0_0),
    .I0_0_1(n72_I0_0_1),
    .I0_1_0(n72_I0_1_0),
    .I0_1_1(n72_I0_1_1),
    .I1_0(n72_I1_0),
    .I1_1(n72_I1_1),
    .O_0_0(n72_O_0_0),
    .O_0_1(n72_O_0_1),
    .O_0_2(n72_O_0_2),
    .O_1_0(n72_O_1_0),
    .O_1_1(n72_O_1_1),
    .O_1_2(n72_O_1_2)
  );
  MapT n81 ( // @[Top.scala 113:21]
    .valid_up(n81_valid_up),
    .valid_down(n81_valid_down),
    .I_0_0(n81_I_0_0),
    .I_0_1(n81_I_0_1),
    .I_0_2(n81_I_0_2),
    .I_1_0(n81_I_1_0),
    .I_1_1(n81_I_1_1),
    .I_1_2(n81_I_1_2),
    .O_0_0_0(n81_O_0_0_0),
    .O_0_0_1(n81_O_0_0_1),
    .O_0_0_2(n81_O_0_0_2),
    .O_1_0_0(n81_O_1_0_0),
    .O_1_0_1(n81_O_1_0_1),
    .O_1_0_2(n81_O_1_0_2)
  );
  MapT_1 n88 ( // @[Top.scala 116:21]
    .valid_up(n88_valid_up),
    .valid_down(n88_valid_down),
    .I_0_0_0(n88_I_0_0_0),
    .I_0_0_1(n88_I_0_0_1),
    .I_0_0_2(n88_I_0_0_2),
    .I_1_0_0(n88_I_1_0_0),
    .I_1_0_1(n88_I_1_0_1),
    .I_1_0_2(n88_I_1_0_2),
    .O_0_0(n88_O_0_0),
    .O_0_1(n88_O_0_1),
    .O_0_2(n88_O_0_2),
    .O_1_0(n88_O_1_0),
    .O_1_1(n88_O_1_1),
    .O_1_2(n88_O_1_2)
  );
  Map2T_7 n89 ( // @[Top.scala 119:21]
    .valid_up(n89_valid_up),
    .valid_down(n89_valid_down),
    .I0_0_0_0(n89_I0_0_0_0),
    .I0_0_0_1(n89_I0_0_0_1),
    .I0_0_0_2(n89_I0_0_0_2),
    .I0_0_1_0(n89_I0_0_1_0),
    .I0_0_1_1(n89_I0_0_1_1),
    .I0_0_1_2(n89_I0_0_1_2),
    .I0_1_0_0(n89_I0_1_0_0),
    .I0_1_0_1(n89_I0_1_0_1),
    .I0_1_0_2(n89_I0_1_0_2),
    .I0_1_1_0(n89_I0_1_1_0),
    .I0_1_1_1(n89_I0_1_1_1),
    .I0_1_1_2(n89_I0_1_1_2),
    .I1_0_0(n89_I1_0_0),
    .I1_0_1(n89_I1_0_1),
    .I1_0_2(n89_I1_0_2),
    .I1_1_0(n89_I1_1_0),
    .I1_1_1(n89_I1_1_1),
    .I1_1_2(n89_I1_1_2),
    .O_0_0_0(n89_O_0_0_0),
    .O_0_0_1(n89_O_0_0_1),
    .O_0_0_2(n89_O_0_0_2),
    .O_0_1_0(n89_O_0_1_0),
    .O_0_1_1(n89_O_0_1_1),
    .O_0_1_2(n89_O_0_1_2),
    .O_0_2_0(n89_O_0_2_0),
    .O_0_2_1(n89_O_0_2_1),
    .O_0_2_2(n89_O_0_2_2),
    .O_1_0_0(n89_O_1_0_0),
    .O_1_0_1(n89_O_1_0_1),
    .O_1_0_2(n89_O_1_0_2),
    .O_1_1_0(n89_O_1_1_0),
    .O_1_1_1(n89_O_1_1_1),
    .O_1_1_2(n89_O_1_1_2),
    .O_1_2_0(n89_O_1_2_0),
    .O_1_2_1(n89_O_1_2_1),
    .O_1_2_2(n89_O_1_2_2)
  );
  MapT_6 n98 ( // @[Top.scala 123:21]
    .valid_up(n98_valid_up),
    .valid_down(n98_valid_down),
    .I_0_0_0(n98_I_0_0_0),
    .I_0_0_1(n98_I_0_0_1),
    .I_0_0_2(n98_I_0_0_2),
    .I_0_1_0(n98_I_0_1_0),
    .I_0_1_1(n98_I_0_1_1),
    .I_0_1_2(n98_I_0_1_2),
    .I_0_2_0(n98_I_0_2_0),
    .I_0_2_1(n98_I_0_2_1),
    .I_0_2_2(n98_I_0_2_2),
    .I_1_0_0(n98_I_1_0_0),
    .I_1_0_1(n98_I_1_0_1),
    .I_1_0_2(n98_I_1_0_2),
    .I_1_1_0(n98_I_1_1_0),
    .I_1_1_1(n98_I_1_1_1),
    .I_1_1_2(n98_I_1_1_2),
    .I_1_2_0(n98_I_1_2_0),
    .I_1_2_1(n98_I_1_2_1),
    .I_1_2_2(n98_I_1_2_2),
    .O_0_0_0_0(n98_O_0_0_0_0),
    .O_0_0_0_1(n98_O_0_0_0_1),
    .O_0_0_0_2(n98_O_0_0_0_2),
    .O_0_0_1_0(n98_O_0_0_1_0),
    .O_0_0_1_1(n98_O_0_0_1_1),
    .O_0_0_1_2(n98_O_0_0_1_2),
    .O_0_0_2_0(n98_O_0_0_2_0),
    .O_0_0_2_1(n98_O_0_0_2_1),
    .O_0_0_2_2(n98_O_0_0_2_2),
    .O_1_0_0_0(n98_O_1_0_0_0),
    .O_1_0_0_1(n98_O_1_0_0_1),
    .O_1_0_0_2(n98_O_1_0_0_2),
    .O_1_0_1_0(n98_O_1_0_1_0),
    .O_1_0_1_1(n98_O_1_0_1_1),
    .O_1_0_1_2(n98_O_1_0_1_2),
    .O_1_0_2_0(n98_O_1_0_2_0),
    .O_1_0_2_1(n98_O_1_0_2_1),
    .O_1_0_2_2(n98_O_1_0_2_2)
  );
  MapT_7 n105 ( // @[Top.scala 126:22]
    .valid_up(n105_valid_up),
    .valid_down(n105_valid_down),
    .I_0_0_0_0(n105_I_0_0_0_0),
    .I_0_0_0_1(n105_I_0_0_0_1),
    .I_0_0_0_2(n105_I_0_0_0_2),
    .I_0_0_1_0(n105_I_0_0_1_0),
    .I_0_0_1_1(n105_I_0_0_1_1),
    .I_0_0_1_2(n105_I_0_0_1_2),
    .I_0_0_2_0(n105_I_0_0_2_0),
    .I_0_0_2_1(n105_I_0_0_2_1),
    .I_0_0_2_2(n105_I_0_0_2_2),
    .I_1_0_0_0(n105_I_1_0_0_0),
    .I_1_0_0_1(n105_I_1_0_0_1),
    .I_1_0_0_2(n105_I_1_0_0_2),
    .I_1_0_1_0(n105_I_1_0_1_0),
    .I_1_0_1_1(n105_I_1_0_1_1),
    .I_1_0_1_2(n105_I_1_0_1_2),
    .I_1_0_2_0(n105_I_1_0_2_0),
    .I_1_0_2_1(n105_I_1_0_2_1),
    .I_1_0_2_2(n105_I_1_0_2_2),
    .O_0_0_0(n105_O_0_0_0),
    .O_0_0_1(n105_O_0_0_1),
    .O_0_0_2(n105_O_0_0_2),
    .O_0_1_0(n105_O_0_1_0),
    .O_0_1_1(n105_O_0_1_1),
    .O_0_1_2(n105_O_0_1_2),
    .O_0_2_0(n105_O_0_2_0),
    .O_0_2_1(n105_O_0_2_1),
    .O_0_2_2(n105_O_0_2_2),
    .O_1_0_0(n105_O_1_0_0),
    .O_1_0_1(n105_O_1_0_1),
    .O_1_0_2(n105_O_1_0_2),
    .O_1_1_0(n105_O_1_1_0),
    .O_1_1_1(n105_O_1_1_1),
    .O_1_1_2(n105_O_1_1_2),
    .O_1_2_0(n105_O_1_2_0),
    .O_1_2_1(n105_O_1_2_1),
    .O_1_2_2(n105_O_1_2_2)
  );
  MapT_8 n147 ( // @[Top.scala 129:22]
    .clock(n147_clock),
    .reset(n147_reset),
    .valid_up(n147_valid_up),
    .valid_down(n147_valid_down),
    .I_0_0_0(n147_I_0_0_0),
    .I_0_0_1(n147_I_0_0_1),
    .I_0_0_2(n147_I_0_0_2),
    .I_0_1_0(n147_I_0_1_0),
    .I_0_1_1(n147_I_0_1_1),
    .I_0_1_2(n147_I_0_1_2),
    .I_0_2_0(n147_I_0_2_0),
    .I_0_2_1(n147_I_0_2_1),
    .I_0_2_2(n147_I_0_2_2),
    .I_1_0_0(n147_I_1_0_0),
    .I_1_0_1(n147_I_1_0_1),
    .I_1_0_2(n147_I_1_0_2),
    .I_1_1_0(n147_I_1_1_0),
    .I_1_1_1(n147_I_1_1_1),
    .I_1_1_2(n147_I_1_1_2),
    .I_1_2_0(n147_I_1_2_0),
    .I_1_2_1(n147_I_1_2_1),
    .I_1_2_2(n147_I_1_2_2),
    .O_0_0_0(n147_O_0_0_0),
    .O_1_0_0(n147_O_1_0_0)
  );
  Passthrough n148 ( // @[Top.scala 132:22]
    .valid_up(n148_valid_up),
    .valid_down(n148_valid_down),
    .I_0_0_0(n148_I_0_0_0),
    .I_1_0_0(n148_I_1_0_0),
    .O_0_0(n148_O_0_0),
    .O_1_0(n148_O_1_0)
  );
  Passthrough_1 n149 ( // @[Top.scala 135:22]
    .valid_up(n149_valid_up),
    .valid_down(n149_valid_down),
    .I_0_0(n149_I_0_0),
    .I_1_0(n149_I_1_0),
    .O_0(n149_O_0),
    .O_1(n149_O_1)
  );
  FIFO n150 ( // @[Top.scala 138:22]
    .clock(n150_clock),
    .reset(n150_reset),
    .valid_up(n150_valid_up),
    .valid_down(n150_valid_down),
    .I_0(n150_I_0),
    .I_1(n150_I_1),
    .O_0(n150_O_0),
    .O_1(n150_O_1)
  );
  FIFO n151 ( // @[Top.scala 141:22]
    .clock(n151_clock),
    .reset(n151_reset),
    .valid_up(n151_valid_up),
    .valid_down(n151_valid_down),
    .I_0(n151_I_0),
    .I_1(n151_I_1),
    .O_0(n151_O_0),
    .O_1(n151_O_1)
  );
  FIFO n152 ( // @[Top.scala 144:22]
    .clock(n152_clock),
    .reset(n152_reset),
    .valid_up(n152_valid_up),
    .valid_down(n152_valid_down),
    .I_0(n152_I_0),
    .I_1(n152_I_1),
    .O_0(n152_O_0),
    .O_1(n152_O_1)
  );
  assign valid_down = n152_valid_down; // @[Top.scala 148:16]
  assign O_0 = n152_O_0; // @[Top.scala 147:7]
  assign O_1 = n152_O_1; // @[Top.scala 147:7]
  assign n1_clock = clock;
  assign n1_reset = reset;
  assign n1_valid_up = valid_up; // @[Top.scala 48:17]
  assign n1_I_0 = I_0; // @[Top.scala 47:10]
  assign n1_I_1 = I_1; // @[Top.scala 47:10]
  assign n2_clock = clock;
  assign n2_reset = reset;
  assign n2_valid_up = n1_valid_down; // @[Top.scala 51:17]
  assign n2_I_0 = n1_O_0; // @[Top.scala 50:10]
  assign n2_I_1 = n1_O_1; // @[Top.scala 50:10]
  assign n3_clock = clock;
  assign n3_reset = reset;
  assign n3_valid_up = n2_valid_down; // @[Top.scala 54:17]
  assign n3_I_0 = n2_O_0; // @[Top.scala 53:10]
  assign n3_I_1 = n2_O_1; // @[Top.scala 53:10]
  assign n4_clock = clock;
  assign n4_valid_up = n3_valid_down; // @[Top.scala 57:17]
  assign n4_I_0 = n3_O_0; // @[Top.scala 56:10]
  assign n4_I_1 = n3_O_1; // @[Top.scala 56:10]
  assign n5_clock = clock;
  assign n5_valid_up = n4_valid_down; // @[Top.scala 60:17]
  assign n5_I_0 = n4_O_0; // @[Top.scala 59:10]
  assign n5_I_1 = n4_O_1; // @[Top.scala 59:10]
  assign n6_valid_up = n5_valid_down & n4_valid_down; // @[Top.scala 64:17]
  assign n6_I0_0 = n5_O_0; // @[Top.scala 62:11]
  assign n6_I0_1 = n5_O_1; // @[Top.scala 62:11]
  assign n6_I1_0 = n4_O_0; // @[Top.scala 63:11]
  assign n6_I1_1 = n4_O_1; // @[Top.scala 63:11]
  assign n13_valid_up = n6_valid_down & n3_valid_down; // @[Top.scala 68:18]
  assign n13_I0_0_0 = n6_O_0_0; // @[Top.scala 66:12]
  assign n13_I0_0_1 = n6_O_0_1; // @[Top.scala 66:12]
  assign n13_I0_1_0 = n6_O_1_0; // @[Top.scala 66:12]
  assign n13_I0_1_1 = n6_O_1_1; // @[Top.scala 66:12]
  assign n13_I1_0 = n3_O_0; // @[Top.scala 67:12]
  assign n13_I1_1 = n3_O_1; // @[Top.scala 67:12]
  assign n22_valid_up = n13_valid_down; // @[Top.scala 71:18]
  assign n22_I_0_0 = n13_O_0_0; // @[Top.scala 70:11]
  assign n22_I_0_1 = n13_O_0_1; // @[Top.scala 70:11]
  assign n22_I_0_2 = n13_O_0_2; // @[Top.scala 70:11]
  assign n22_I_1_0 = n13_O_1_0; // @[Top.scala 70:11]
  assign n22_I_1_1 = n13_O_1_1; // @[Top.scala 70:11]
  assign n22_I_1_2 = n13_O_1_2; // @[Top.scala 70:11]
  assign n29_valid_up = n22_valid_down; // @[Top.scala 74:18]
  assign n29_I_0_0_0 = n22_O_0_0_0; // @[Top.scala 73:11]
  assign n29_I_0_0_1 = n22_O_0_0_1; // @[Top.scala 73:11]
  assign n29_I_0_0_2 = n22_O_0_0_2; // @[Top.scala 73:11]
  assign n29_I_1_0_0 = n22_O_1_0_0; // @[Top.scala 73:11]
  assign n29_I_1_0_1 = n22_O_1_0_1; // @[Top.scala 73:11]
  assign n29_I_1_0_2 = n22_O_1_0_2; // @[Top.scala 73:11]
  assign n30_clock = clock;
  assign n30_valid_up = n2_valid_down; // @[Top.scala 77:18]
  assign n30_I_0 = n2_O_0; // @[Top.scala 76:11]
  assign n30_I_1 = n2_O_1; // @[Top.scala 76:11]
  assign n31_clock = clock;
  assign n31_valid_up = n30_valid_down; // @[Top.scala 80:18]
  assign n31_I_0 = n30_O_0; // @[Top.scala 79:11]
  assign n31_I_1 = n30_O_1; // @[Top.scala 79:11]
  assign n32_valid_up = n31_valid_down & n30_valid_down; // @[Top.scala 84:18]
  assign n32_I0_0 = n31_O_0; // @[Top.scala 82:12]
  assign n32_I0_1 = n31_O_1; // @[Top.scala 82:12]
  assign n32_I1_0 = n30_O_0; // @[Top.scala 83:12]
  assign n32_I1_1 = n30_O_1; // @[Top.scala 83:12]
  assign n39_valid_up = n32_valid_down & n2_valid_down; // @[Top.scala 88:18]
  assign n39_I0_0_0 = n32_O_0_0; // @[Top.scala 86:12]
  assign n39_I0_0_1 = n32_O_0_1; // @[Top.scala 86:12]
  assign n39_I0_1_0 = n32_O_1_0; // @[Top.scala 86:12]
  assign n39_I0_1_1 = n32_O_1_1; // @[Top.scala 86:12]
  assign n39_I1_0 = n2_O_0; // @[Top.scala 87:12]
  assign n39_I1_1 = n2_O_1; // @[Top.scala 87:12]
  assign n48_valid_up = n39_valid_down; // @[Top.scala 91:18]
  assign n48_I_0_0 = n39_O_0_0; // @[Top.scala 90:11]
  assign n48_I_0_1 = n39_O_0_1; // @[Top.scala 90:11]
  assign n48_I_0_2 = n39_O_0_2; // @[Top.scala 90:11]
  assign n48_I_1_0 = n39_O_1_0; // @[Top.scala 90:11]
  assign n48_I_1_1 = n39_O_1_1; // @[Top.scala 90:11]
  assign n48_I_1_2 = n39_O_1_2; // @[Top.scala 90:11]
  assign n55_valid_up = n48_valid_down; // @[Top.scala 94:18]
  assign n55_I_0_0_0 = n48_O_0_0_0; // @[Top.scala 93:11]
  assign n55_I_0_0_1 = n48_O_0_0_1; // @[Top.scala 93:11]
  assign n55_I_0_0_2 = n48_O_0_0_2; // @[Top.scala 93:11]
  assign n55_I_1_0_0 = n48_O_1_0_0; // @[Top.scala 93:11]
  assign n55_I_1_0_1 = n48_O_1_0_1; // @[Top.scala 93:11]
  assign n55_I_1_0_2 = n48_O_1_0_2; // @[Top.scala 93:11]
  assign n56_valid_up = n29_valid_down & n55_valid_down; // @[Top.scala 98:18]
  assign n56_I0_0_0 = n29_O_0_0; // @[Top.scala 96:12]
  assign n56_I0_0_1 = n29_O_0_1; // @[Top.scala 96:12]
  assign n56_I0_0_2 = n29_O_0_2; // @[Top.scala 96:12]
  assign n56_I0_1_0 = n29_O_1_0; // @[Top.scala 96:12]
  assign n56_I0_1_1 = n29_O_1_1; // @[Top.scala 96:12]
  assign n56_I0_1_2 = n29_O_1_2; // @[Top.scala 96:12]
  assign n56_I1_0_0 = n55_O_0_0; // @[Top.scala 97:12]
  assign n56_I1_0_1 = n55_O_0_1; // @[Top.scala 97:12]
  assign n56_I1_0_2 = n55_O_0_2; // @[Top.scala 97:12]
  assign n56_I1_1_0 = n55_O_1_0; // @[Top.scala 97:12]
  assign n56_I1_1_1 = n55_O_1_1; // @[Top.scala 97:12]
  assign n56_I1_1_2 = n55_O_1_2; // @[Top.scala 97:12]
  assign n63_clock = clock;
  assign n63_valid_up = n1_valid_down; // @[Top.scala 101:18]
  assign n63_I_0 = n1_O_0; // @[Top.scala 100:11]
  assign n63_I_1 = n1_O_1; // @[Top.scala 100:11]
  assign n64_clock = clock;
  assign n64_valid_up = n63_valid_down; // @[Top.scala 104:18]
  assign n64_I_0 = n63_O_0; // @[Top.scala 103:11]
  assign n64_I_1 = n63_O_1; // @[Top.scala 103:11]
  assign n65_valid_up = n64_valid_down & n63_valid_down; // @[Top.scala 108:18]
  assign n65_I0_0 = n64_O_0; // @[Top.scala 106:12]
  assign n65_I0_1 = n64_O_1; // @[Top.scala 106:12]
  assign n65_I1_0 = n63_O_0; // @[Top.scala 107:12]
  assign n65_I1_1 = n63_O_1; // @[Top.scala 107:12]
  assign n72_valid_up = n65_valid_down & n1_valid_down; // @[Top.scala 112:18]
  assign n72_I0_0_0 = n65_O_0_0; // @[Top.scala 110:12]
  assign n72_I0_0_1 = n65_O_0_1; // @[Top.scala 110:12]
  assign n72_I0_1_0 = n65_O_1_0; // @[Top.scala 110:12]
  assign n72_I0_1_1 = n65_O_1_1; // @[Top.scala 110:12]
  assign n72_I1_0 = n1_O_0; // @[Top.scala 111:12]
  assign n72_I1_1 = n1_O_1; // @[Top.scala 111:12]
  assign n81_valid_up = n72_valid_down; // @[Top.scala 115:18]
  assign n81_I_0_0 = n72_O_0_0; // @[Top.scala 114:11]
  assign n81_I_0_1 = n72_O_0_1; // @[Top.scala 114:11]
  assign n81_I_0_2 = n72_O_0_2; // @[Top.scala 114:11]
  assign n81_I_1_0 = n72_O_1_0; // @[Top.scala 114:11]
  assign n81_I_1_1 = n72_O_1_1; // @[Top.scala 114:11]
  assign n81_I_1_2 = n72_O_1_2; // @[Top.scala 114:11]
  assign n88_valid_up = n81_valid_down; // @[Top.scala 118:18]
  assign n88_I_0_0_0 = n81_O_0_0_0; // @[Top.scala 117:11]
  assign n88_I_0_0_1 = n81_O_0_0_1; // @[Top.scala 117:11]
  assign n88_I_0_0_2 = n81_O_0_0_2; // @[Top.scala 117:11]
  assign n88_I_1_0_0 = n81_O_1_0_0; // @[Top.scala 117:11]
  assign n88_I_1_0_1 = n81_O_1_0_1; // @[Top.scala 117:11]
  assign n88_I_1_0_2 = n81_O_1_0_2; // @[Top.scala 117:11]
  assign n89_valid_up = n56_valid_down & n88_valid_down; // @[Top.scala 122:18]
  assign n89_I0_0_0_0 = n56_O_0_0_0; // @[Top.scala 120:12]
  assign n89_I0_0_0_1 = n56_O_0_0_1; // @[Top.scala 120:12]
  assign n89_I0_0_0_2 = n56_O_0_0_2; // @[Top.scala 120:12]
  assign n89_I0_0_1_0 = n56_O_0_1_0; // @[Top.scala 120:12]
  assign n89_I0_0_1_1 = n56_O_0_1_1; // @[Top.scala 120:12]
  assign n89_I0_0_1_2 = n56_O_0_1_2; // @[Top.scala 120:12]
  assign n89_I0_1_0_0 = n56_O_1_0_0; // @[Top.scala 120:12]
  assign n89_I0_1_0_1 = n56_O_1_0_1; // @[Top.scala 120:12]
  assign n89_I0_1_0_2 = n56_O_1_0_2; // @[Top.scala 120:12]
  assign n89_I0_1_1_0 = n56_O_1_1_0; // @[Top.scala 120:12]
  assign n89_I0_1_1_1 = n56_O_1_1_1; // @[Top.scala 120:12]
  assign n89_I0_1_1_2 = n56_O_1_1_2; // @[Top.scala 120:12]
  assign n89_I1_0_0 = n88_O_0_0; // @[Top.scala 121:12]
  assign n89_I1_0_1 = n88_O_0_1; // @[Top.scala 121:12]
  assign n89_I1_0_2 = n88_O_0_2; // @[Top.scala 121:12]
  assign n89_I1_1_0 = n88_O_1_0; // @[Top.scala 121:12]
  assign n89_I1_1_1 = n88_O_1_1; // @[Top.scala 121:12]
  assign n89_I1_1_2 = n88_O_1_2; // @[Top.scala 121:12]
  assign n98_valid_up = n89_valid_down; // @[Top.scala 125:18]
  assign n98_I_0_0_0 = n89_O_0_0_0; // @[Top.scala 124:11]
  assign n98_I_0_0_1 = n89_O_0_0_1; // @[Top.scala 124:11]
  assign n98_I_0_0_2 = n89_O_0_0_2; // @[Top.scala 124:11]
  assign n98_I_0_1_0 = n89_O_0_1_0; // @[Top.scala 124:11]
  assign n98_I_0_1_1 = n89_O_0_1_1; // @[Top.scala 124:11]
  assign n98_I_0_1_2 = n89_O_0_1_2; // @[Top.scala 124:11]
  assign n98_I_0_2_0 = n89_O_0_2_0; // @[Top.scala 124:11]
  assign n98_I_0_2_1 = n89_O_0_2_1; // @[Top.scala 124:11]
  assign n98_I_0_2_2 = n89_O_0_2_2; // @[Top.scala 124:11]
  assign n98_I_1_0_0 = n89_O_1_0_0; // @[Top.scala 124:11]
  assign n98_I_1_0_1 = n89_O_1_0_1; // @[Top.scala 124:11]
  assign n98_I_1_0_2 = n89_O_1_0_2; // @[Top.scala 124:11]
  assign n98_I_1_1_0 = n89_O_1_1_0; // @[Top.scala 124:11]
  assign n98_I_1_1_1 = n89_O_1_1_1; // @[Top.scala 124:11]
  assign n98_I_1_1_2 = n89_O_1_1_2; // @[Top.scala 124:11]
  assign n98_I_1_2_0 = n89_O_1_2_0; // @[Top.scala 124:11]
  assign n98_I_1_2_1 = n89_O_1_2_1; // @[Top.scala 124:11]
  assign n98_I_1_2_2 = n89_O_1_2_2; // @[Top.scala 124:11]
  assign n105_valid_up = n98_valid_down; // @[Top.scala 128:19]
  assign n105_I_0_0_0_0 = n98_O_0_0_0_0; // @[Top.scala 127:12]
  assign n105_I_0_0_0_1 = n98_O_0_0_0_1; // @[Top.scala 127:12]
  assign n105_I_0_0_0_2 = n98_O_0_0_0_2; // @[Top.scala 127:12]
  assign n105_I_0_0_1_0 = n98_O_0_0_1_0; // @[Top.scala 127:12]
  assign n105_I_0_0_1_1 = n98_O_0_0_1_1; // @[Top.scala 127:12]
  assign n105_I_0_0_1_2 = n98_O_0_0_1_2; // @[Top.scala 127:12]
  assign n105_I_0_0_2_0 = n98_O_0_0_2_0; // @[Top.scala 127:12]
  assign n105_I_0_0_2_1 = n98_O_0_0_2_1; // @[Top.scala 127:12]
  assign n105_I_0_0_2_2 = n98_O_0_0_2_2; // @[Top.scala 127:12]
  assign n105_I_1_0_0_0 = n98_O_1_0_0_0; // @[Top.scala 127:12]
  assign n105_I_1_0_0_1 = n98_O_1_0_0_1; // @[Top.scala 127:12]
  assign n105_I_1_0_0_2 = n98_O_1_0_0_2; // @[Top.scala 127:12]
  assign n105_I_1_0_1_0 = n98_O_1_0_1_0; // @[Top.scala 127:12]
  assign n105_I_1_0_1_1 = n98_O_1_0_1_1; // @[Top.scala 127:12]
  assign n105_I_1_0_1_2 = n98_O_1_0_1_2; // @[Top.scala 127:12]
  assign n105_I_1_0_2_0 = n98_O_1_0_2_0; // @[Top.scala 127:12]
  assign n105_I_1_0_2_1 = n98_O_1_0_2_1; // @[Top.scala 127:12]
  assign n105_I_1_0_2_2 = n98_O_1_0_2_2; // @[Top.scala 127:12]
  assign n147_clock = clock;
  assign n147_reset = reset;
  assign n147_valid_up = n105_valid_down; // @[Top.scala 131:19]
  assign n147_I_0_0_0 = n105_O_0_0_0; // @[Top.scala 130:12]
  assign n147_I_0_0_1 = n105_O_0_0_1; // @[Top.scala 130:12]
  assign n147_I_0_0_2 = n105_O_0_0_2; // @[Top.scala 130:12]
  assign n147_I_0_1_0 = n105_O_0_1_0; // @[Top.scala 130:12]
  assign n147_I_0_1_1 = n105_O_0_1_1; // @[Top.scala 130:12]
  assign n147_I_0_1_2 = n105_O_0_1_2; // @[Top.scala 130:12]
  assign n147_I_0_2_0 = n105_O_0_2_0; // @[Top.scala 130:12]
  assign n147_I_0_2_1 = n105_O_0_2_1; // @[Top.scala 130:12]
  assign n147_I_0_2_2 = n105_O_0_2_2; // @[Top.scala 130:12]
  assign n147_I_1_0_0 = n105_O_1_0_0; // @[Top.scala 130:12]
  assign n147_I_1_0_1 = n105_O_1_0_1; // @[Top.scala 130:12]
  assign n147_I_1_0_2 = n105_O_1_0_2; // @[Top.scala 130:12]
  assign n147_I_1_1_0 = n105_O_1_1_0; // @[Top.scala 130:12]
  assign n147_I_1_1_1 = n105_O_1_1_1; // @[Top.scala 130:12]
  assign n147_I_1_1_2 = n105_O_1_1_2; // @[Top.scala 130:12]
  assign n147_I_1_2_0 = n105_O_1_2_0; // @[Top.scala 130:12]
  assign n147_I_1_2_1 = n105_O_1_2_1; // @[Top.scala 130:12]
  assign n147_I_1_2_2 = n105_O_1_2_2; // @[Top.scala 130:12]
  assign n148_valid_up = n147_valid_down; // @[Top.scala 134:19]
  assign n148_I_0_0_0 = n147_O_0_0_0; // @[Top.scala 133:12]
  assign n148_I_1_0_0 = n147_O_1_0_0; // @[Top.scala 133:12]
  assign n149_valid_up = n148_valid_down; // @[Top.scala 137:19]
  assign n149_I_0_0 = n148_O_0_0; // @[Top.scala 136:12]
  assign n149_I_1_0 = n148_O_1_0; // @[Top.scala 136:12]
  assign n150_clock = clock;
  assign n150_reset = reset;
  assign n150_valid_up = n149_valid_down; // @[Top.scala 140:19]
  assign n150_I_0 = n149_O_0; // @[Top.scala 139:12]
  assign n150_I_1 = n149_O_1; // @[Top.scala 139:12]
  assign n151_clock = clock;
  assign n151_reset = reset;
  assign n151_valid_up = n150_valid_down; // @[Top.scala 143:19]
  assign n151_I_0 = n150_O_0; // @[Top.scala 142:12]
  assign n151_I_1 = n150_O_1; // @[Top.scala 142:12]
  assign n152_clock = clock;
  assign n152_reset = reset;
  assign n152_valid_up = n151_valid_down; // @[Top.scala 146:19]
  assign n152_I_0 = n151_O_0; // @[Top.scala 145:12]
  assign n152_I_1 = n151_O_1; // @[Top.scala 145:12]
endmodule
