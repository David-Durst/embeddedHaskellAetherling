// Latency = 4
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(clock), // @[:@1296.4]
    .reset('b0), // @[:@1297.4]
    .io_in_x348_TREADY(dontcare), // @[:@1298.4]
    .io_in_x348_TDATA({I_0,I_1}), // @[:@1298.4]
    .io_in_x348_TID(8'h0),
    .io_in_x348_TDEST(8'h0),
    .io_in_x349_TVALID(valid_down), // @[:@1298.4]
    .io_in_x349_TDATA({O_0_0_0,O_1_0_0}), // @[:@1298.4]
    .io_in_x349_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x356_ctrchain cchain ( // @[:@2879.2]
    .clock(clock), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule


module SRAMVerilogSim
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule


module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 311:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 315:12:@24.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : io_wPort_0_data_0; // @[MemPrimitives.scala 315:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 316:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        ff <= io_wPort_0_data_0;
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh14); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh14); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_parentAck, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  _T_81; // @[Controllers.scala 86:43:@328.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_93; // @[Controllers.scala 92:52:@342.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_134; // @[Controllers.scala 129:57:@382.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  wire  _T_167; // @[package.scala 100:41:@414.4]
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign _T_81 = io_rst | done_0_io_output; // @[Controllers.scala 86:43:@328.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_93 = synchronize | io_rst; // @[Controllers.scala 92:52:@342.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_134 = _T_133 | io_parentAck; // @[Controllers.scala 129:57:@382.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign _T_167 = done_0_io_output & _T_166; // @[package.scala 100:41:@414.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_134 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = _T_81 | io_parentAck; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = _T_93 | io_parentAck; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = _T_167 | io_parentAck; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module SRAM( // @[:@507.2]
  input         clock, // @[:@508.4]
  input  [20:0] io_raddr, // @[:@510.4]
  output [7:0]  io_rdata, // @[:@510.4]
  input         io_backpressure // @[:@510.4]
);
  wire [7:0] SRAMVerilogSim_rdata; // @[SRAM.scala 185:23:@512.4]
  wire [7:0] SRAMVerilogSim_wdata; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_backpressure; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_wen; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_waddrEn; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_raddrEn; // @[SRAM.scala 185:23:@512.4]
  wire [20:0] SRAMVerilogSim_waddr; // @[SRAM.scala 185:23:@512.4]
  wire [20:0] SRAMVerilogSim_raddr; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_clk; // @[SRAM.scala 185:23:@512.4]
  SRAMVerilogSim #(.DWIDTH(8), .WORDS(2073600), .AWIDTH(21)) SRAMVerilogSim ( // @[SRAM.scala 185:23:@512.4]
    .rdata(SRAMVerilogSim_rdata),
    .wdata(SRAMVerilogSim_wdata),
    .backpressure(SRAMVerilogSim_backpressure),
    .wen(SRAMVerilogSim_wen),
    .waddrEn(SRAMVerilogSim_waddrEn),
    .raddrEn(SRAMVerilogSim_raddrEn),
    .waddr(SRAMVerilogSim_waddr),
    .raddr(SRAMVerilogSim_raddr),
    .clk(SRAMVerilogSim_clk)
  );
  assign io_rdata = SRAMVerilogSim_rdata; // @[SRAM.scala 195:16:@532.4]
  assign SRAMVerilogSim_wdata = 8'h0; // @[SRAM.scala 190:20:@526.4]
  assign SRAMVerilogSim_backpressure = io_backpressure; // @[SRAM.scala 191:27:@527.4]
  assign SRAMVerilogSim_wen = 1'h0; // @[SRAM.scala 188:18:@524.4]
  assign SRAMVerilogSim_waddrEn = 1'h1; // @[SRAM.scala 193:22:@529.4]
  assign SRAMVerilogSim_raddrEn = 1'h1; // @[SRAM.scala 192:22:@528.4]
  assign SRAMVerilogSim_waddr = 21'h0; // @[SRAM.scala 189:20:@525.4]
  assign SRAMVerilogSim_raddr = io_raddr; // @[SRAM.scala 187:20:@523.4]
  assign SRAMVerilogSim_clk = clock; // @[SRAM.scala 186:18:@522.4]
endmodule
module RetimeWrapper_5( // @[:@546.2]
  input         clock, // @[:@547.4]
  input         reset, // @[:@548.4]
  input         io_flow, // @[:@549.4]
  input  [20:0] io_in, // @[:@549.4]
  output [20:0] io_out // @[:@549.4]
);
  wire [20:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire [20:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire [20:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@551.4]
  RetimeShiftRegister #(.WIDTH(21), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@551.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@564.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@563.4]
  assign sr_init = 21'h0; // @[RetimeShiftRegister.scala 19:16:@562.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@561.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@560.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@558.4]
endmodule
module Mem1D( // @[:@566.2]
  input         clock, // @[:@567.4]
  input         reset, // @[:@568.4]
  input  [20:0] io_r_ofs_0, // @[:@569.4]
  input         io_r_backpressure, // @[:@569.4]
  output [7:0]  io_output // @[:@569.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 705:21:@573.4]
  wire [20:0] SRAM_io_raddr; // @[MemPrimitives.scala 705:21:@573.4]
  wire [7:0] SRAM_io_rdata; // @[MemPrimitives.scala 705:21:@573.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 705:21:@573.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@576.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@576.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@576.4]
  wire [20:0] RetimeWrapper_io_in; // @[package.scala 93:22:@576.4]
  wire [20:0] RetimeWrapper_io_out; // @[package.scala 93:22:@576.4]
  SRAM SRAM ( // @[MemPrimitives.scala 705:21:@573.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@576.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 712:17:@589.4]
  assign SRAM_clock = clock; // @[:@574.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 706:37:@583.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 711:30:@588.4]
  assign RetimeWrapper_clock = clock; // @[:@577.4]
  assign RetimeWrapper_reset = reset; // @[:@578.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@580.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@579.4]
endmodule
module StickySelects( // @[:@591.2]
  input   io_ins_0, // @[:@594.4]
  output  io_outs_0 // @[:@594.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 34:26:@596.4]
endmodule
module RetimeWrapper_6( // @[:@610.2]
  input   clock, // @[:@611.4]
  input   reset, // @[:@612.4]
  input   io_flow, // @[:@613.4]
  input   io_in, // @[:@613.4]
  output  io_out // @[:@613.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@615.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@615.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@628.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@627.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@626.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@625.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@624.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@622.4]
endmodule
module x350_outbuf_0( // @[:@630.2]
  input         clock, // @[:@631.4]
  input         reset, // @[:@632.4]
  input  [20:0] io_rPort_0_ofs_0, // @[:@633.4]
  input         io_rPort_0_en_0, // @[:@633.4]
  input         io_rPort_0_backpressure, // @[:@633.4]
  output [7:0]  io_rPort_0_output_0 // @[:@633.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@648.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@648.4]
  wire [20:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@648.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@648.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@648.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@674.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@674.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@688.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@688.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@688.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@688.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@688.4]
  wire  _T_76; // @[MemPrimitives.scala 123:41:@678.4]
  wire [22:0] _T_78; // @[Cat.scala 30:58:@680.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@648.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@674.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@688.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@678.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@680.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 148:13:@695.4]
  assign Mem1D_clock = clock; // @[:@649.4]
  assign Mem1D_reset = reset; // @[:@650.4]
  assign Mem1D_io_r_ofs_0 = _T_78[20:0]; // @[MemPrimitives.scala 127:28:@684.4]
  assign Mem1D_io_r_backpressure = _T_78[21]; // @[MemPrimitives.scala 128:32:@685.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 122:60:@677.4]
  assign RetimeWrapper_clock = clock; // @[:@689.4]
  assign RetimeWrapper_reset = reset; // @[:@690.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@692.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@691.4]
endmodule
module x607_sm( // @[:@839.2]
  input   clock, // @[:@840.4]
  input   reset, // @[:@841.4]
  input   io_enable, // @[:@842.4]
  output  io_done, // @[:@842.4]
  input   io_ctrDone, // @[:@842.4]
  output  io_ctrInc, // @[:@842.4]
  input   io_parentAck, // @[:@842.4]
  input   io_doneIn_0, // @[:@842.4]
  input   io_doneIn_1, // @[:@842.4]
  output  io_enableOut_0, // @[:@842.4]
  output  io_enableOut_1, // @[:@842.4]
  output  io_childAck_0, // @[:@842.4]
  output  io_childAck_1 // @[:@842.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@845.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@848.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@851.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@854.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@886.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1004.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1004.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1004.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1004.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1004.4]
  wire  allDone; // @[Controllers.scala 80:47:@857.4]
  wire  synchronize; // @[Controllers.scala 146:56:@911.4]
  wire  _T_127; // @[Controllers.scala 150:35:@913.4]
  wire  _T_129; // @[Controllers.scala 150:60:@914.4]
  wire  _T_130; // @[Controllers.scala 150:58:@915.4]
  wire  _T_132; // @[Controllers.scala 150:76:@916.4]
  wire  _T_133; // @[Controllers.scala 150:74:@917.4]
  wire  _T_135; // @[Controllers.scala 150:97:@918.4]
  wire  _T_136; // @[Controllers.scala 150:95:@919.4]
  wire  _T_152; // @[Controllers.scala 150:35:@937.4]
  wire  _T_154; // @[Controllers.scala 150:60:@938.4]
  wire  _T_155; // @[Controllers.scala 150:58:@939.4]
  wire  _T_157; // @[Controllers.scala 150:76:@940.4]
  wire  _T_158; // @[Controllers.scala 150:74:@941.4]
  wire  _T_161; // @[Controllers.scala 150:95:@943.4]
  wire  _T_179; // @[Controllers.scala 213:68:@965.4]
  wire  _T_181; // @[Controllers.scala 213:90:@967.4]
  wire  _T_183; // @[Controllers.scala 213:132:@969.4]
  wire  _T_184; // @[Controllers.scala 213:130:@970.4]
  wire  _T_185; // @[Controllers.scala 213:156:@971.4]
  wire  _T_187; // @[Controllers.scala 213:68:@974.4]
  wire  _T_189; // @[Controllers.scala 213:90:@976.4]
  wire  _T_196; // @[package.scala 100:49:@982.4]
  reg  _T_199; // @[package.scala 48:56:@983.4]
  reg [31:0] _RAND_0;
  wire  _T_200; // @[package.scala 100:41:@985.4]
  reg  _T_213; // @[package.scala 48:56:@1001.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@845.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@848.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@851.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@854.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@883.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@886.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@987.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1004.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@857.4]
  assign synchronize = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 146:56:@911.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 150:35:@913.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 150:60:@914.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 150:58:@915.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 150:76:@916.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 150:74:@917.4]
  assign _T_135 = io_ctrDone == 1'h0; // @[Controllers.scala 150:97:@918.4]
  assign _T_136 = _T_133 & _T_135; // @[Controllers.scala 150:95:@919.4]
  assign _T_152 = ~ iterDone_1_io_output; // @[Controllers.scala 150:35:@937.4]
  assign _T_154 = io_doneIn_1 == 1'h0; // @[Controllers.scala 150:60:@938.4]
  assign _T_155 = _T_152 & _T_154; // @[Controllers.scala 150:58:@939.4]
  assign _T_157 = done_1_io_output == 1'h0; // @[Controllers.scala 150:76:@940.4]
  assign _T_158 = _T_155 & _T_157; // @[Controllers.scala 150:74:@941.4]
  assign _T_161 = _T_158 & _T_135; // @[Controllers.scala 150:95:@943.4]
  assign _T_179 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@965.4]
  assign _T_181 = _T_179 & _T_127; // @[Controllers.scala 213:90:@967.4]
  assign _T_183 = ~ allDone; // @[Controllers.scala 213:132:@969.4]
  assign _T_184 = _T_181 & _T_183; // @[Controllers.scala 213:130:@970.4]
  assign _T_185 = ~ io_ctrDone; // @[Controllers.scala 213:156:@971.4]
  assign _T_187 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@974.4]
  assign _T_189 = _T_187 & _T_152; // @[Controllers.scala 213:90:@976.4]
  assign _T_196 = allDone == 1'h0; // @[package.scala 100:49:@982.4]
  assign _T_200 = allDone & _T_199; // @[package.scala 100:41:@985.4]
  assign io_done = RetimeWrapper_1_io_out; // @[Controllers.scala 245:13:@1011.4]
  assign io_ctrInc = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 143:17:@910.4]
  assign io_enableOut_0 = _T_184 & _T_185; // @[Controllers.scala 213:55:@973.4]
  assign io_enableOut_1 = _T_189 & _T_183; // @[Controllers.scala 213:55:@981.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@962.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@964.4]
  assign active_0_clock = clock; // @[:@846.4]
  assign active_0_reset = reset; // @[:@847.4]
  assign active_0_io_input_set = _T_136 & io_enable; // @[Controllers.scala 150:32:@922.4]
  assign active_0_io_input_reset = io_doneIn_0 | io_parentAck; // @[Controllers.scala 151:34:@926.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@860.4]
  assign active_1_clock = clock; // @[:@849.4]
  assign active_1_reset = reset; // @[:@850.4]
  assign active_1_io_input_set = _T_161 & io_enable; // @[Controllers.scala 150:32:@946.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_parentAck; // @[Controllers.scala 151:34:@950.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@861.4]
  assign done_0_clock = clock; // @[:@852.4]
  assign done_0_reset = reset; // @[:@853.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@936.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@872.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@862.4]
  assign done_1_clock = clock; // @[:@855.4]
  assign done_1_reset = reset; // @[:@856.4]
  assign done_1_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@960.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@881.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@863.4]
  assign iterDone_0_clock = clock; // @[:@884.4]
  assign iterDone_0_reset = reset; // @[:@885.4]
  assign iterDone_0_io_input_set = io_doneIn_0; // @[Controllers.scala 152:34:@932.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@899.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@889.4]
  assign iterDone_1_clock = clock; // @[:@887.4]
  assign iterDone_1_reset = reset; // @[:@888.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 152:34:@956.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@908.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@890.4]
  assign RetimeWrapper_clock = clock; // @[:@988.4]
  assign RetimeWrapper_reset = reset; // @[:@989.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@991.4]
  assign RetimeWrapper_io_in = _T_200 | io_parentAck; // @[package.scala 94:16:@990.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1005.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1006.4]
  assign RetimeWrapper_1_io_flow = io_enable; // @[package.scala 95:18:@1008.4]
  assign RetimeWrapper_1_io_in = allDone & _T_213; // @[package.scala 94:16:@1007.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_199 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_213 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_199 <= 1'h0;
    end else begin
      _T_199 <= _T_196;
    end
    if (reset) begin
      _T_213 <= 1'h0;
    end else begin
      _T_213 <= _T_196;
    end
  end
endmodule
module x528_outr_UnitPipe_sm( // @[:@1428.2]
  input   clock, // @[:@1429.4]
  input   reset, // @[:@1430.4]
  input   io_enable, // @[:@1431.4]
  output  io_done, // @[:@1431.4]
  input   io_parentAck, // @[:@1431.4]
  input   io_doneIn_0, // @[:@1431.4]
  input   io_doneIn_1, // @[:@1431.4]
  output  io_enableOut_0, // @[:@1431.4]
  output  io_enableOut_1, // @[:@1431.4]
  output  io_childAck_0, // @[:@1431.4]
  output  io_childAck_1, // @[:@1431.4]
  input   io_ctrCopyDone_0, // @[:@1431.4]
  input   io_ctrCopyDone_1 // @[:@1431.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@1434.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@1437.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@1440.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1443.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1475.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1681.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1681.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1681.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1681.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1681.4]
  wire  allDone; // @[Controllers.scala 80:47:@1446.4]
  wire  _T_127; // @[Controllers.scala 165:35:@1500.4]
  wire  _T_129; // @[Controllers.scala 165:60:@1501.4]
  wire  _T_130; // @[Controllers.scala 165:58:@1502.4]
  wire  _T_132; // @[Controllers.scala 165:76:@1503.4]
  wire  _T_133; // @[Controllers.scala 165:74:@1504.4]
  wire  _T_137; // @[Controllers.scala 165:109:@1507.4]
  wire  _T_140; // @[Controllers.scala 165:141:@1509.4]
  wire  _T_148; // @[package.scala 96:25:@1521.4 package.scala 96:25:@1522.4]
  wire  _T_152; // @[Controllers.scala 167:54:@1524.4]
  wire  _T_153; // @[Controllers.scala 167:52:@1525.4]
  wire  _T_160; // @[package.scala 96:25:@1535.4 package.scala 96:25:@1536.4]
  wire  _T_178; // @[package.scala 96:25:@1553.4 package.scala 96:25:@1554.4]
  wire  _T_182; // @[Controllers.scala 169:67:@1556.4]
  wire  _T_183; // @[Controllers.scala 169:86:@1557.4]
  wire  _T_195; // @[Controllers.scala 165:35:@1569.4]
  wire  _T_197; // @[Controllers.scala 165:60:@1570.4]
  wire  _T_198; // @[Controllers.scala 165:58:@1571.4]
  wire  _T_200; // @[Controllers.scala 165:76:@1572.4]
  wire  _T_201; // @[Controllers.scala 165:74:@1573.4]
  wire  _T_205; // @[Controllers.scala 165:109:@1576.4]
  wire  _T_208; // @[Controllers.scala 165:141:@1578.4]
  wire  _T_216; // @[package.scala 96:25:@1590.4 package.scala 96:25:@1591.4]
  wire  _T_220; // @[Controllers.scala 167:54:@1593.4]
  wire  _T_221; // @[Controllers.scala 167:52:@1594.4]
  wire  _T_228; // @[package.scala 96:25:@1604.4 package.scala 96:25:@1605.4]
  wire  _T_246; // @[package.scala 96:25:@1622.4 package.scala 96:25:@1623.4]
  wire  _T_250; // @[Controllers.scala 169:67:@1625.4]
  wire  _T_251; // @[Controllers.scala 169:86:@1626.4]
  wire  _T_265; // @[Controllers.scala 213:68:@1642.4]
  wire  _T_267; // @[Controllers.scala 213:90:@1644.4]
  wire  _T_269; // @[Controllers.scala 213:132:@1646.4]
  wire  _T_273; // @[Controllers.scala 213:68:@1651.4]
  wire  _T_275; // @[Controllers.scala 213:90:@1653.4]
  wire  _T_282; // @[package.scala 100:49:@1659.4]
  reg  _T_285; // @[package.scala 48:56:@1660.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@1662.4]
  reg  _T_299; // @[package.scala 48:56:@1678.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@1434.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@1437.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@1440.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1443.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1472.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1475.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1516.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1530.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1548.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1585.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1599.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1617.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1664.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1681.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1446.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1500.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1501.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@1502.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1503.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@1504.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@1507.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1509.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@1521.4 package.scala 96:25:@1522.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@1524.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@1525.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1535.4 package.scala 96:25:@1536.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1553.4 package.scala 96:25:@1554.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@1556.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@1557.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1569.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1570.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@1571.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1572.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@1573.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@1576.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1578.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1590.4 package.scala 96:25:@1591.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@1593.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@1594.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1604.4 package.scala 96:25:@1605.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1622.4 package.scala 96:25:@1623.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@1625.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@1626.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1642.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@1644.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@1646.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1651.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@1653.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@1659.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@1662.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@1688.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@1650.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@1658.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1639.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1641.4]
  assign active_0_clock = clock; // @[:@1435.4]
  assign active_0_reset = reset; // @[:@1436.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@1511.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1515.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1449.4]
  assign active_1_clock = clock; // @[:@1438.4]
  assign active_1_reset = reset; // @[:@1439.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@1580.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1584.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1450.4]
  assign done_0_clock = clock; // @[:@1441.4]
  assign done_0_reset = reset; // @[:@1442.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@1561.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1461.4 Controllers.scala 170:32:@1568.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1451.4]
  assign done_1_clock = clock; // @[:@1444.4]
  assign done_1_reset = reset; // @[:@1445.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@1630.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1470.4 Controllers.scala 170:32:@1637.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1452.4]
  assign iterDone_0_clock = clock; // @[:@1473.4]
  assign iterDone_0_reset = reset; // @[:@1474.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@1529.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@1488.4 Controllers.scala 168:36:@1545.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1478.4]
  assign iterDone_1_clock = clock; // @[:@1476.4]
  assign iterDone_1_reset = reset; // @[:@1477.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@1598.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@1497.4 Controllers.scala 168:36:@1614.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1479.4]
  assign RetimeWrapper_clock = clock; // @[:@1517.4]
  assign RetimeWrapper_reset = reset; // @[:@1518.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1520.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1519.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1531.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1532.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1534.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1533.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1549.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1550.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1552.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1551.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1586.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1587.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1589.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1588.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1600.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1601.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1603.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1602.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1618.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1619.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1621.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1620.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1665.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1666.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1668.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@1667.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1682.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1683.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@1685.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@1684.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module CompactingIncDincCtr( // @[:@1917.2]
  input   clock, // @[:@1918.4]
  input   reset, // @[:@1919.4]
  input   io_input_inc_en_0, // @[:@1920.4]
  input   io_input_dinc_en_0, // @[:@1920.4]
  output  io_output_full // @[:@1920.4]
);
  reg [31:0] cnt; // @[Counter.scala 170:20:@1922.4]
  reg [31:0] _RAND_0;
  wire [14:0] numPushed; // @[Counter.scala 172:47:@1923.4]
  wire [14:0] numPopped; // @[Counter.scala 173:48:@1924.4]
  wire [31:0] _GEN_0; // @[Counter.scala 174:14:@1925.4]
  wire [32:0] _T_37; // @[Counter.scala 174:14:@1925.4]
  wire [31:0] _T_38; // @[Counter.scala 174:14:@1926.4]
  wire [31:0] _T_39; // @[Counter.scala 174:14:@1927.4]
  wire [31:0] _GEN_1; // @[Counter.scala 174:26:@1928.4]
  wire [32:0] _T_40; // @[Counter.scala 174:26:@1928.4]
  wire [31:0] _T_41; // @[Counter.scala 174:26:@1929.4]
  wire [31:0] _T_42; // @[Counter.scala 174:26:@1930.4]
  assign numPushed = io_input_inc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 172:47:@1923.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 173:48:@1924.4]
  assign _GEN_0 = {{17{numPushed[14]}},numPushed}; // @[Counter.scala 174:14:@1925.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1925.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1926.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 174:14:@1927.4]
  assign _GEN_1 = {{17{numPopped[14]}},numPopped}; // @[Counter.scala 174:26:@1928.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1928.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1929.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 174:26:@1930.4]
  assign io_output_full = $signed(cnt) > $signed(32'sh1dff); // @[Counter.scala 180:18:@1944.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module x351_fifoinraw_0( // @[:@2067.2]
  input   clock, // @[:@2068.4]
  input   reset // @[:@2069.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 382:24:@2114.4]
  wire  elements_reset; // @[MemPrimitives.scala 382:24:@2114.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 382:24:@2114.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 382:24:@2114.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 382:24:@2114.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 382:24:@2114.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign elements_clock = clock; // @[:@2115.4]
  assign elements_reset = reset; // @[:@2116.4]
  assign elements_io_input_inc_en_0 = 1'h0; // @[MemPrimitives.scala 384:79:@2126.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 385:80:@2127.4]
endmodule
module x352_fifoinpacked_0( // @[:@2490.2]
  input   clock, // @[:@2491.4]
  input   reset, // @[:@2492.4]
  input   io_wPort_0_en_0, // @[:@2493.4]
  output  io_full, // @[:@2493.4]
  input   io_active_0_in, // @[:@2493.4]
  output  io_active_0_out // @[:@2493.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 382:24:@2537.4]
  wire  elements_reset; // @[MemPrimitives.scala 382:24:@2537.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 382:24:@2537.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 382:24:@2537.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 382:24:@2537.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 382:24:@2537.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 429:39:@2611.4]
  assign io_active_0_out = io_active_0_in; // @[MemPrimitives.scala 427:129:@2609.4]
  assign elements_clock = clock; // @[:@2538.4]
  assign elements_reset = reset; // @[:@2539.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 384:79:@2549.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 385:80:@2550.4]
endmodule
module FF_7( // @[:@3040.2]
  input         clock, // @[:@3041.4]
  input         reset, // @[:@3042.4]
  output [12:0] io_rPort_0_output_0, // @[:@3043.4]
  input  [12:0] io_wPort_0_data_0, // @[:@3043.4]
  input         io_wPort_0_reset, // @[:@3043.4]
  input         io_wPort_0_en_0 // @[:@3043.4]
);
  reg [12:0] ff; // @[MemPrimitives.scala 311:19:@3058.4]
  reg [31:0] _RAND_0;
  wire [12:0] _T_68; // @[MemPrimitives.scala 315:32:@3060.4]
  wire [12:0] _T_69; // @[MemPrimitives.scala 315:12:@3061.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 315:32:@3060.4]
  assign _T_69 = io_wPort_0_reset ? 13'h0 : _T_68; // @[MemPrimitives.scala 315:12:@3061.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 316:34:@3063.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 13'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 13'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_1( // @[:@3078.2]
  input         clock, // @[:@3079.4]
  input         reset, // @[:@3080.4]
  input         io_setup_saturate, // @[:@3081.4]
  input         io_input_reset, // @[:@3081.4]
  input         io_input_enable, // @[:@3081.4]
  output [12:0] io_output_count_0, // @[:@3081.4]
  output        io_output_oobs_0, // @[:@3081.4]
  output        io_output_done, // @[:@3081.4]
  output        io_output_saturated // @[:@3081.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3094.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3094.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3094.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3094.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3094.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3094.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3110.4]
  wire  _T_36; // @[Counter.scala 264:45:@3113.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3138.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3139.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3140.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3141.4]
  wire  _T_57; // @[Counter.scala 293:18:@3143.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3151.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3153.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3154.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3155.4]
  wire  _T_75; // @[Counter.scala 322:102:@3159.4]
  wire  _T_77; // @[Counter.scala 322:130:@3160.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3094.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3110.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3113.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3138.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3139.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3140.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3141.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh438); // @[Counter.scala 293:18:@3143.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3151.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3153.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3154.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3155.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3159.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh438); // @[Counter.scala 322:130:@3160.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3158.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3162.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3164.4]
  assign io_output_saturated = io_setup_saturate & _T_57; // @[Counter.scala 340:25:@3167.4]
  assign bases_0_clock = clock; // @[:@3095.4]
  assign bases_0_reset = reset; // @[:@3096.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3157.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3136.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3137.4]
  assign SRFF_clock = clock; // @[:@3111.4]
  assign SRFF_reset = reset; // @[:@3112.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3115.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3117.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3118.4]
endmodule
module SingleCounter_2( // @[:@3207.2]
  input         clock, // @[:@3208.4]
  input         reset, // @[:@3209.4]
  input         io_setup_saturate, // @[:@3210.4]
  input         io_input_reset, // @[:@3210.4]
  input         io_input_enable, // @[:@3210.4]
  output [12:0] io_output_count_0, // @[:@3210.4]
  output        io_output_oobs_0, // @[:@3210.4]
  output        io_output_done // @[:@3210.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3223.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3223.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3223.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3223.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3223.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3223.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3239.4]
  wire  _T_36; // @[Counter.scala 264:45:@3242.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3267.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3268.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3269.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3270.4]
  wire  _T_57; // @[Counter.scala 293:18:@3272.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3280.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3282.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3283.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3284.4]
  wire  _T_75; // @[Counter.scala 322:102:@3288.4]
  wire  _T_77; // @[Counter.scala 322:130:@3289.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3223.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3239.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3242.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3267.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh2); // @[Counter.scala 291:33:@3268.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh2); // @[Counter.scala 291:33:@3269.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3270.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh780); // @[Counter.scala 293:18:@3272.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3280.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3282.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3283.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3284.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3288.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh780); // @[Counter.scala 322:130:@3289.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3287.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3291.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3293.4]
  assign bases_0_clock = clock; // @[:@3224.4]
  assign bases_0_reset = reset; // @[:@3225.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3286.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3265.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3266.4]
  assign SRFF_clock = clock; // @[:@3240.4]
  assign SRFF_reset = reset; // @[:@3241.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3244.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3246.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3247.4]
endmodule
module x356_ctrchain( // @[:@3298.2]
  input         clock, // @[:@3299.4]
  input         reset, // @[:@3300.4]
  input         io_input_reset, // @[:@3301.4]
  input         io_input_enable, // @[:@3301.4]
  output [12:0] io_output_counts_1, // @[:@3301.4]
  output [12:0] io_output_counts_0, // @[:@3301.4]
  output        io_output_oobs_0, // @[:@3301.4]
  output        io_output_oobs_1, // @[:@3301.4]
  output        io_output_done // @[:@3301.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@3303.4]
  wire [12:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@3306.4]
  wire [12:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@3306.4]
  wire  isDone; // @[Counter.scala 541:51:@3323.4]
  reg  wasDone; // @[Counter.scala 542:24:@3324.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@3332.4]
  wire  _T_66; // @[Counter.scala 546:80:@3333.4]
  reg  doneLatch; // @[Counter.scala 550:26:@3338.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@3339.4]
  wire  _T_74; // @[Counter.scala 551:19:@3340.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@3303.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@3306.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@3323.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@3332.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@3333.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@3339.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@3340.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@3345.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@3342.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3344.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3347.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@3335.4]
  assign ctrs_0_clock = clock; // @[:@3304.4]
  assign ctrs_0_reset = reset; // @[:@3305.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 530:29:@3320.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3312.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@3319.4]
  assign ctrs_1_clock = clock; // @[:@3307.4]
  assign ctrs_1_reset = reset; // @[:@3308.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@3322.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3316.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@3317.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_21( // @[:@3387.2]
  input   clock, // @[:@3388.4]
  input   reset, // @[:@3389.4]
  input   io_flow, // @[:@3390.4]
  input   io_in, // @[:@3390.4]
  output  io_out // @[:@3390.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@3392.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3405.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3404.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3403.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3402.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3401.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3399.4]
endmodule
module RetimeWrapper_25( // @[:@3515.2]
  input   clock, // @[:@3516.4]
  input   reset, // @[:@3517.4]
  input   io_flow, // @[:@3518.4]
  input   io_in, // @[:@3518.4]
  output  io_out // @[:@3518.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@3520.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3533.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3532.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3531.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3530.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3529.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3527.4]
endmodule
module x374_inr_Foreach_sm( // @[:@3535.2]
  input   clock, // @[:@3536.4]
  input   reset, // @[:@3537.4]
  input   io_enable, // @[:@3538.4]
  output  io_done, // @[:@3538.4]
  output  io_doneLatch, // @[:@3538.4]
  input   io_ctrDone, // @[:@3538.4]
  output  io_datapathEn, // @[:@3538.4]
  output  io_ctrInc, // @[:@3538.4]
  output  io_ctrRst, // @[:@3538.4]
  input   io_parentAck, // @[:@3538.4]
  input   io_backpressure, // @[:@3538.4]
  input   io_break // @[:@3538.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3540.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3540.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3540.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3540.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3540.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3540.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3543.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3543.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3543.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3543.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3543.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3543.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3635.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3635.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3635.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3635.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3635.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3548.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3549.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3550.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3551.4]
  wire  _T_100; // @[package.scala 100:49:@3568.4]
  reg  _T_103; // @[package.scala 48:56:@3569.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3582.4 package.scala 96:25:@3583.4]
  wire  _T_110; // @[package.scala 100:49:@3584.4]
  reg  _T_113; // @[package.scala 48:56:@3585.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3587.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3592.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3593.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3596.4]
  wire  _T_124; // @[package.scala 96:25:@3604.4 package.scala 96:25:@3605.4]
  wire  _T_126; // @[package.scala 100:49:@3606.4]
  reg  _T_129; // @[package.scala 48:56:@3607.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3629.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3631.4]
  reg  _T_153; // @[package.scala 48:56:@3632.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3640.4 package.scala 96:25:@3641.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3642.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3643.4]
  SRFF active ( // @[Controllers.scala 261:22:@3540.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3543.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@3577.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3599.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3611.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3619.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@3635.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3548.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3549.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3550.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3551.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3568.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3582.4 package.scala 96:25:@3583.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3584.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3587.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3592.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3593.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3596.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3604.4 package.scala 96:25:@3605.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3606.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3631.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3640.4 package.scala 96:25:@3641.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3642.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3643.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3610.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3645.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3595.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3598.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3590.4]
  assign active_clock = clock; // @[:@3541.4]
  assign active_reset = reset; // @[:@3542.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3553.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3557.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3558.4]
  assign done_clock = clock; // @[:@3544.4]
  assign done_reset = reset; // @[:@3545.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3573.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3566.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3567.4]
  assign RetimeWrapper_clock = clock; // @[:@3578.4]
  assign RetimeWrapper_reset = reset; // @[:@3579.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3581.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3580.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3600.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3601.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3603.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3602.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3612.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3613.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3615.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3614.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3620.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3621.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3623.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3622.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3636.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3637.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3639.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3638.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SimBlackBoxesfix2fixBox( // @[:@3752.2]
  input  [31:0] io_a, // @[:@3755.4]
  output [31:0] io_b // @[:@3755.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@3768.4]
endmodule
module _( // @[:@3770.2]
  input  [31:0] io_b, // @[:@3773.4]
  output [31:0] io_result // @[:@3773.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3778.4]
  wire [31:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3778.4]
  SimBlackBoxesfix2fixBox SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3778.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3791.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3786.4]
endmodule
module SimBlackBoxesfix2fixBox_2( // @[:@3834.2]
  input  [31:0] io_a, // @[:@3837.4]
  output [32:0] io_b // @[:@3837.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@3847.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@3847.4]
  assign io_b = {_T_20,io_a}; // @[SimBlackBoxes.scala 99:40:@3852.4]
endmodule
module __2( // @[:@3854.2]
  input  [31:0] io_b, // @[:@3857.4]
  output [32:0] io_result // @[:@3857.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3862.4]
  wire [32:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3862.4]
  SimBlackBoxesfix2fixBox_2 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3862.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3875.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3870.4]
endmodule
module RetimeWrapper_29( // @[:@3932.2]
  input         clock, // @[:@3933.4]
  input         reset, // @[:@3934.4]
  input         io_flow, // @[:@3935.4]
  input  [31:0] io_in, // @[:@3935.4]
  output [31:0] io_out // @[:@3935.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3937.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3950.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3949.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3948.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3947.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3946.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3944.4]
endmodule
module fix2fixBox( // @[:@3952.2]
  input         clock, // @[:@3953.4]
  input         reset, // @[:@3954.4]
  input  [32:0] io_a, // @[:@3955.4]
  input         io_flow, // @[:@3955.4]
  output [31:0] io_b // @[:@3955.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3968.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3968.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3968.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3968.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3968.4]
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@3968.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@3975.4]
  assign RetimeWrapper_clock = clock; // @[:@3969.4]
  assign RetimeWrapper_reset = reset; // @[:@3970.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@3972.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@3971.4]
endmodule
module x577_sub( // @[:@3977.2]
  input         clock, // @[:@3978.4]
  input         reset, // @[:@3979.4]
  input  [31:0] io_a, // @[:@3980.4]
  input  [31:0] io_b, // @[:@3980.4]
  input         io_flow, // @[:@3980.4]
  output [31:0] io_result // @[:@3980.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@3988.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@3988.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@3995.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@3995.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@4014.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@4014.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@4014.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@4014.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@4014.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@3993.4 Math.scala 713:14:@3994.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@4000.4 Math.scala 713:14:@4001.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@4002.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@4003.4]
  __2 _ ( // @[Math.scala 709:24:@3988.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@3995.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 182:30:@4014.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@3993.4 Math.scala 713:14:@3994.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@4000.4 Math.scala 713:14:@4001.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@4002.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@4003.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@4022.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@3991.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@3998.4]
  assign fix2fixBox_clock = clock; // @[:@4015.4]
  assign fix2fixBox_reset = reset; // @[:@4016.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@4017.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@4020.4]
endmodule
module x362_sum( // @[:@4199.2]
  input         clock, // @[:@4200.4]
  input         reset, // @[:@4201.4]
  input  [31:0] io_a, // @[:@4202.4]
  input  [31:0] io_b, // @[:@4202.4]
  input         io_flow, // @[:@4202.4]
  output [31:0] io_result // @[:@4202.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@4210.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@4210.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@4217.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@4217.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4235.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4235.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4235.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4235.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4235.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@4215.4 Math.scala 713:14:@4216.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@4222.4 Math.scala 713:14:@4223.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@4224.4]
  __2 _ ( // @[Math.scala 709:24:@4210.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@4217.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 141:30:@4235.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@4215.4 Math.scala 713:14:@4216.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@4222.4 Math.scala 713:14:@4223.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4224.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4243.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@4213.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@4220.4]
  assign fix2fixBox_clock = clock; // @[:@4236.4]
  assign fix2fixBox_reset = reset; // @[:@4237.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4238.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4241.4]
endmodule
module x374_inr_Foreach_kernelx374_inr_Foreach_concrete1( // @[:@5179.2]
  input         clock, // @[:@5180.4]
  input         reset, // @[:@5181.4]
  output        io_in_x352_fifoinpacked_0_wPort_0_en_0, // @[:@5182.4]
  input         io_in_x352_fifoinpacked_0_full, // @[:@5182.4]
  output        io_in_x352_fifoinpacked_0_active_0_in, // @[:@5182.4]
  input         io_in_x352_fifoinpacked_0_active_0_out, // @[:@5182.4]
  input         io_sigsIn_backpressure, // @[:@5182.4]
  input         io_sigsIn_datapathEn, // @[:@5182.4]
  input         io_sigsIn_break, // @[:@5182.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_1, // @[:@5182.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@5182.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@5182.4]
  input         io_sigsIn_cchainOutputs_0_oobs_1, // @[:@5182.4]
  input         io_rr // @[:@5182.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@5216.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@5216.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@5228.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@5228.4]
  wire  x577_sub_1_clock; // @[Math.scala 191:24:@5255.4]
  wire  x577_sub_1_reset; // @[Math.scala 191:24:@5255.4]
  wire [31:0] x577_sub_1_io_a; // @[Math.scala 191:24:@5255.4]
  wire [31:0] x577_sub_1_io_b; // @[Math.scala 191:24:@5255.4]
  wire  x577_sub_1_io_flow; // @[Math.scala 191:24:@5255.4]
  wire [31:0] x577_sub_1_io_result; // @[Math.scala 191:24:@5255.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@5265.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@5265.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@5265.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@5265.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@5265.4]
  wire  x362_sum_1_clock; // @[Math.scala 150:24:@5274.4]
  wire  x362_sum_1_reset; // @[Math.scala 150:24:@5274.4]
  wire [31:0] x362_sum_1_io_a; // @[Math.scala 150:24:@5274.4]
  wire [31:0] x362_sum_1_io_b; // @[Math.scala 150:24:@5274.4]
  wire  x362_sum_1_io_flow; // @[Math.scala 150:24:@5274.4]
  wire [31:0] x362_sum_1_io_result; // @[Math.scala 150:24:@5274.4]
  wire  x363_sum_1_clock; // @[Math.scala 150:24:@5286.4]
  wire  x363_sum_1_reset; // @[Math.scala 150:24:@5286.4]
  wire [31:0] x363_sum_1_io_a; // @[Math.scala 150:24:@5286.4]
  wire [31:0] x363_sum_1_io_b; // @[Math.scala 150:24:@5286.4]
  wire  x363_sum_1_io_flow; // @[Math.scala 150:24:@5286.4]
  wire [31:0] x363_sum_1_io_result; // @[Math.scala 150:24:@5286.4]
  wire  x579_sum_1_clock; // @[Math.scala 150:24:@5301.4]
  wire  x579_sum_1_reset; // @[Math.scala 150:24:@5301.4]
  wire [31:0] x579_sum_1_io_a; // @[Math.scala 150:24:@5301.4]
  wire [31:0] x579_sum_1_io_b; // @[Math.scala 150:24:@5301.4]
  wire  x579_sum_1_io_flow; // @[Math.scala 150:24:@5301.4]
  wire [31:0] x579_sum_1_io_result; // @[Math.scala 150:24:@5301.4]
  wire  x367_sum_1_clock; // @[Math.scala 150:24:@5333.4]
  wire  x367_sum_1_reset; // @[Math.scala 150:24:@5333.4]
  wire [31:0] x367_sum_1_io_a; // @[Math.scala 150:24:@5333.4]
  wire [31:0] x367_sum_1_io_b; // @[Math.scala 150:24:@5333.4]
  wire  x367_sum_1_io_flow; // @[Math.scala 150:24:@5333.4]
  wire [31:0] x367_sum_1_io_result; // @[Math.scala 150:24:@5333.4]
  wire  x582_sum_1_clock; // @[Math.scala 150:24:@5348.4]
  wire  x582_sum_1_reset; // @[Math.scala 150:24:@5348.4]
  wire [31:0] x582_sum_1_io_a; // @[Math.scala 150:24:@5348.4]
  wire [31:0] x582_sum_1_io_b; // @[Math.scala 150:24:@5348.4]
  wire  x582_sum_1_io_flow; // @[Math.scala 150:24:@5348.4]
  wire [31:0] x582_sum_1_io_result; // @[Math.scala 150:24:@5348.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@5384.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@5384.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@5384.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@5384.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@5384.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@5393.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@5393.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@5393.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@5393.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@5393.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@5404.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@5404.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@5404.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@5404.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@5404.4]
  wire  _T_327; // @[sm_x374_inr_Foreach.scala 62:18:@5241.4]
  wire  _T_328; // @[sm_x374_inr_Foreach.scala 62:55:@5242.4]
  wire [31:0] b357_number; // @[Math.scala 712:22:@5221.4 Math.scala 713:14:@5222.4]
  wire [42:0] _GEN_0; // @[Math.scala 450:32:@5246.4]
  wire [42:0] _T_332; // @[Math.scala 450:32:@5246.4]
  wire [38:0] _GEN_1; // @[Math.scala 450:32:@5251.4]
  wire [38:0] _T_336; // @[Math.scala 450:32:@5251.4]
  wire [31:0] x363_sum_number; // @[Math.scala 154:22:@5292.4 Math.scala 155:14:@5293.4]
  wire [33:0] _GEN_2; // @[Math.scala 450:32:@5297.4]
  wire [33:0] _T_356; // @[Math.scala 450:32:@5297.4]
  wire [31:0] x367_sum_number; // @[Math.scala 154:22:@5339.4 Math.scala 155:14:@5340.4]
  wire [33:0] _GEN_3; // @[Math.scala 450:32:@5344.4]
  wire [33:0] _T_385; // @[Math.scala 450:32:@5344.4]
  wire  _T_419; // @[sm_x374_inr_Foreach.scala 103:131:@5401.4]
  wire  _T_423; // @[package.scala 96:25:@5409.4 package.scala 96:25:@5410.4]
  wire  _T_425; // @[implicits.scala 55:10:@5411.4]
  wire  _T_426; // @[sm_x374_inr_Foreach.scala 103:148:@5412.4]
  wire  _T_428; // @[sm_x374_inr_Foreach.scala 103:236:@5414.4]
  wire  _T_429; // @[sm_x374_inr_Foreach.scala 103:255:@5415.4]
  wire  x610_b359_D4; // @[package.scala 96:25:@5389.4 package.scala 96:25:@5390.4]
  wire  _T_432; // @[sm_x374_inr_Foreach.scala 103:291:@5417.4]
  wire  x611_b360_D4; // @[package.scala 96:25:@5398.4 package.scala 96:25:@5399.4]
  _ _ ( // @[Math.scala 709:24:@5216.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@5228.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x577_sub x577_sub_1 ( // @[Math.scala 191:24:@5255.4]
    .clock(x577_sub_1_clock),
    .reset(x577_sub_1_reset),
    .io_a(x577_sub_1_io_a),
    .io_b(x577_sub_1_io_b),
    .io_flow(x577_sub_1_io_flow),
    .io_result(x577_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@5265.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x362_sum x362_sum_1 ( // @[Math.scala 150:24:@5274.4]
    .clock(x362_sum_1_clock),
    .reset(x362_sum_1_reset),
    .io_a(x362_sum_1_io_a),
    .io_b(x362_sum_1_io_b),
    .io_flow(x362_sum_1_io_flow),
    .io_result(x362_sum_1_io_result)
  );
  x362_sum x363_sum_1 ( // @[Math.scala 150:24:@5286.4]
    .clock(x363_sum_1_clock),
    .reset(x363_sum_1_reset),
    .io_a(x363_sum_1_io_a),
    .io_b(x363_sum_1_io_b),
    .io_flow(x363_sum_1_io_flow),
    .io_result(x363_sum_1_io_result)
  );
  x362_sum x579_sum_1 ( // @[Math.scala 150:24:@5301.4]
    .clock(x579_sum_1_clock),
    .reset(x579_sum_1_reset),
    .io_a(x579_sum_1_io_a),
    .io_b(x579_sum_1_io_b),
    .io_flow(x579_sum_1_io_flow),
    .io_result(x579_sum_1_io_result)
  );
  x362_sum x367_sum_1 ( // @[Math.scala 150:24:@5333.4]
    .clock(x367_sum_1_clock),
    .reset(x367_sum_1_reset),
    .io_a(x367_sum_1_io_a),
    .io_b(x367_sum_1_io_b),
    .io_flow(x367_sum_1_io_flow),
    .io_result(x367_sum_1_io_result)
  );
  x362_sum x582_sum_1 ( // @[Math.scala 150:24:@5348.4]
    .clock(x582_sum_1_clock),
    .reset(x582_sum_1_reset),
    .io_a(x582_sum_1_io_a),
    .io_b(x582_sum_1_io_b),
    .io_flow(x582_sum_1_io_flow),
    .io_result(x582_sum_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@5384.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_2 ( // @[package.scala 93:22:@5393.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_3 ( // @[package.scala 93:22:@5404.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_327 = ~ io_in_x352_fifoinpacked_0_full; // @[sm_x374_inr_Foreach.scala 62:18:@5241.4]
  assign _T_328 = ~ io_in_x352_fifoinpacked_0_active_0_out; // @[sm_x374_inr_Foreach.scala 62:55:@5242.4]
  assign b357_number = __io_result; // @[Math.scala 712:22:@5221.4 Math.scala 713:14:@5222.4]
  assign _GEN_0 = {{11'd0}, b357_number}; // @[Math.scala 450:32:@5246.4]
  assign _T_332 = _GEN_0 << 11; // @[Math.scala 450:32:@5246.4]
  assign _GEN_1 = {{7'd0}, b357_number}; // @[Math.scala 450:32:@5251.4]
  assign _T_336 = _GEN_1 << 7; // @[Math.scala 450:32:@5251.4]
  assign x363_sum_number = x363_sum_1_io_result; // @[Math.scala 154:22:@5292.4 Math.scala 155:14:@5293.4]
  assign _GEN_2 = {{2'd0}, x363_sum_number}; // @[Math.scala 450:32:@5297.4]
  assign _T_356 = _GEN_2 << 2; // @[Math.scala 450:32:@5297.4]
  assign x367_sum_number = x367_sum_1_io_result; // @[Math.scala 154:22:@5339.4 Math.scala 155:14:@5340.4]
  assign _GEN_3 = {{2'd0}, x367_sum_number}; // @[Math.scala 450:32:@5344.4]
  assign _T_385 = _GEN_3 << 2; // @[Math.scala 450:32:@5344.4]
  assign _T_419 = ~ io_sigsIn_break; // @[sm_x374_inr_Foreach.scala 103:131:@5401.4]
  assign _T_423 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@5409.4 package.scala 96:25:@5410.4]
  assign _T_425 = io_rr ? _T_423 : 1'h0; // @[implicits.scala 55:10:@5411.4]
  assign _T_426 = _T_419 & _T_425; // @[sm_x374_inr_Foreach.scala 103:148:@5412.4]
  assign _T_428 = _T_426 & _T_419; // @[sm_x374_inr_Foreach.scala 103:236:@5414.4]
  assign _T_429 = _T_428 & io_sigsIn_backpressure; // @[sm_x374_inr_Foreach.scala 103:255:@5415.4]
  assign x610_b359_D4 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@5389.4 package.scala 96:25:@5390.4]
  assign _T_432 = _T_429 & x610_b359_D4; // @[sm_x374_inr_Foreach.scala 103:291:@5417.4]
  assign x611_b360_D4 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@5398.4 package.scala 96:25:@5399.4]
  assign io_in_x352_fifoinpacked_0_wPort_0_en_0 = _T_432 & x611_b360_D4; // @[MemInterfaceType.scala 93:57:@5421.4]
  assign io_in_x352_fifoinpacked_0_active_0_in = x610_b359_D4 & x611_b360_D4; // @[MemInterfaceType.scala 147:18:@5424.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@5219.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@5231.4]
  assign x577_sub_1_clock = clock; // @[:@5256.4]
  assign x577_sub_1_reset = reset; // @[:@5257.4]
  assign x577_sub_1_io_a = _T_332[31:0]; // @[Math.scala 192:17:@5258.4]
  assign x577_sub_1_io_b = _T_336[31:0]; // @[Math.scala 193:17:@5259.4]
  assign x577_sub_1_io_flow = _T_327 | _T_328; // @[Math.scala 194:20:@5260.4]
  assign RetimeWrapper_clock = clock; // @[:@5266.4]
  assign RetimeWrapper_reset = reset; // @[:@5267.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5269.4]
  assign RetimeWrapper_io_in = __1_io_result; // @[package.scala 94:16:@5268.4]
  assign x362_sum_1_clock = clock; // @[:@5275.4]
  assign x362_sum_1_reset = reset; // @[:@5276.4]
  assign x362_sum_1_io_a = x577_sub_1_io_result; // @[Math.scala 151:17:@5277.4]
  assign x362_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@5278.4]
  assign x362_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5279.4]
  assign x363_sum_1_clock = clock; // @[:@5287.4]
  assign x363_sum_1_reset = reset; // @[:@5288.4]
  assign x363_sum_1_io_a = x362_sum_1_io_result; // @[Math.scala 151:17:@5289.4]
  assign x363_sum_1_io_b = 32'h1; // @[Math.scala 152:17:@5290.4]
  assign x363_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5291.4]
  assign x579_sum_1_clock = clock; // @[:@5302.4]
  assign x579_sum_1_reset = reset; // @[:@5303.4]
  assign x579_sum_1_io_a = _T_356[31:0]; // @[Math.scala 151:17:@5304.4]
  assign x579_sum_1_io_b = x363_sum_1_io_result; // @[Math.scala 152:17:@5305.4]
  assign x579_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5306.4]
  assign x367_sum_1_clock = clock; // @[:@5334.4]
  assign x367_sum_1_reset = reset; // @[:@5335.4]
  assign x367_sum_1_io_a = x362_sum_1_io_result; // @[Math.scala 151:17:@5336.4]
  assign x367_sum_1_io_b = 32'h2; // @[Math.scala 152:17:@5337.4]
  assign x367_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5338.4]
  assign x582_sum_1_clock = clock; // @[:@5349.4]
  assign x582_sum_1_reset = reset; // @[:@5350.4]
  assign x582_sum_1_io_a = _T_385[31:0]; // @[Math.scala 151:17:@5351.4]
  assign x582_sum_1_io_b = x367_sum_1_io_result; // @[Math.scala 152:17:@5352.4]
  assign x582_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5353.4]
  assign RetimeWrapper_1_clock = clock; // @[:@5385.4]
  assign RetimeWrapper_1_reset = reset; // @[:@5386.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5388.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@5387.4]
  assign RetimeWrapper_2_clock = clock; // @[:@5394.4]
  assign RetimeWrapper_2_reset = reset; // @[:@5395.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5397.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@5396.4]
  assign RetimeWrapper_3_clock = clock; // @[:@5405.4]
  assign RetimeWrapper_3_reset = reset; // @[:@5406.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5408.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5407.4]
endmodule
module RetimeWrapper_44( // @[:@6542.2]
  input   clock, // @[:@6543.4]
  input   reset, // @[:@6544.4]
  input   io_flow, // @[:@6545.4]
  input   io_in, // @[:@6545.4]
  output  io_out // @[:@6545.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6547.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6547.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6547.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6547.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6547.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6547.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@6547.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6560.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6559.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6558.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6557.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6556.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6554.4]
endmodule
module RetimeWrapper_48( // @[:@6670.2]
  input   clock, // @[:@6671.4]
  input   reset, // @[:@6672.4]
  input   io_flow, // @[:@6673.4]
  input   io_in, // @[:@6673.4]
  output  io_out // @[:@6673.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6675.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6675.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6675.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6675.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6675.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6675.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(19)) sr ( // @[RetimeShiftRegister.scala 15:20:@6675.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6688.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6687.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6686.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6685.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6684.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6682.4]
endmodule
module x526_inr_Foreach_SAMPLER_BOX_sm( // @[:@6690.2]
  input   clock, // @[:@6691.4]
  input   reset, // @[:@6692.4]
  input   io_enable, // @[:@6693.4]
  output  io_done, // @[:@6693.4]
  output  io_doneLatch, // @[:@6693.4]
  input   io_ctrDone, // @[:@6693.4]
  output  io_datapathEn, // @[:@6693.4]
  output  io_ctrInc, // @[:@6693.4]
  output  io_ctrRst, // @[:@6693.4]
  input   io_parentAck, // @[:@6693.4]
  input   io_backpressure, // @[:@6693.4]
  input   io_break // @[:@6693.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@6695.4]
  wire  active_reset; // @[Controllers.scala 261:22:@6695.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@6695.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@6695.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@6695.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@6695.4]
  wire  done_clock; // @[Controllers.scala 262:20:@6698.4]
  wire  done_reset; // @[Controllers.scala 262:20:@6698.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@6698.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@6698.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@6698.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@6698.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6732.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6732.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6732.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@6732.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@6732.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6754.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6754.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6754.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6754.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6754.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6766.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6766.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6766.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6766.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6766.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6774.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6774.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6774.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6774.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6774.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@6790.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@6790.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@6790.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@6790.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@6790.4]
  wire  _T_80; // @[Controllers.scala 264:48:@6703.4]
  wire  _T_81; // @[Controllers.scala 264:46:@6704.4]
  wire  _T_82; // @[Controllers.scala 264:62:@6705.4]
  wire  _T_83; // @[Controllers.scala 264:60:@6706.4]
  wire  _T_100; // @[package.scala 100:49:@6723.4]
  reg  _T_103; // @[package.scala 48:56:@6724.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@6737.4 package.scala 96:25:@6738.4]
  wire  _T_110; // @[package.scala 100:49:@6739.4]
  reg  _T_113; // @[package.scala 48:56:@6740.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@6742.4]
  wire  _T_118; // @[Controllers.scala 283:41:@6747.4]
  wire  _T_119; // @[Controllers.scala 283:59:@6748.4]
  wire  _T_121; // @[Controllers.scala 284:37:@6751.4]
  wire  _T_124; // @[package.scala 96:25:@6759.4 package.scala 96:25:@6760.4]
  wire  _T_126; // @[package.scala 100:49:@6761.4]
  reg  _T_129; // @[package.scala 48:56:@6762.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@6784.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@6786.4]
  reg  _T_153; // @[package.scala 48:56:@6787.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@6795.4 package.scala 96:25:@6796.4]
  wire  _T_158; // @[Controllers.scala 292:61:@6797.4]
  wire  _T_159; // @[Controllers.scala 292:24:@6798.4]
  SRFF active ( // @[Controllers.scala 261:22:@6695.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@6698.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_44 RetimeWrapper ( // @[package.scala 93:22:@6732.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_1 ( // @[package.scala 93:22:@6754.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@6766.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@6774.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_48 RetimeWrapper_4 ( // @[package.scala 93:22:@6790.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@6703.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@6704.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@6705.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@6706.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@6723.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@6737.4 package.scala 96:25:@6738.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@6739.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@6742.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@6747.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@6748.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@6751.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6759.4 package.scala 96:25:@6760.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@6761.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@6786.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@6795.4 package.scala 96:25:@6796.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@6797.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@6798.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@6765.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@6800.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@6750.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@6753.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@6745.4]
  assign active_clock = clock; // @[:@6696.4]
  assign active_reset = reset; // @[:@6697.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@6708.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@6712.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@6713.4]
  assign done_clock = clock; // @[:@6699.4]
  assign done_reset = reset; // @[:@6700.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@6728.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@6721.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@6722.4]
  assign RetimeWrapper_clock = clock; // @[:@6733.4]
  assign RetimeWrapper_reset = reset; // @[:@6734.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@6736.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@6735.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6755.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6756.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@6758.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@6757.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6767.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6768.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@6770.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@6769.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6775.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6776.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@6778.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@6777.4]
  assign RetimeWrapper_4_clock = clock; // @[:@6791.4]
  assign RetimeWrapper_4_reset = reset; // @[:@6792.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@6794.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@6793.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module RetimeWrapper_52( // @[:@7001.2]
  input         clock, // @[:@7002.4]
  input         reset, // @[:@7003.4]
  input         io_flow, // @[:@7004.4]
  input  [15:0] io_in, // @[:@7004.4]
  output [15:0] io_out // @[:@7004.4]
);
  wire [15:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@7006.4]
  wire [15:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@7006.4]
  wire [15:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@7006.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@7006.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@7006.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@7006.4]
  RetimeShiftRegister #(.WIDTH(16), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@7006.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@7019.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@7018.4]
  assign sr_init = 16'h0; // @[RetimeShiftRegister.scala 19:16:@7017.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@7016.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@7015.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@7013.4]
endmodule
module SRAM_1( // @[:@7037.2]
  input        clock, // @[:@7038.4]
  input  [8:0] io_raddr, // @[:@7040.4]
  input        io_wen, // @[:@7040.4]
  input  [8:0] io_waddr, // @[:@7040.4]
  input  [7:0] io_wdata, // @[:@7040.4]
  output [7:0] io_rdata, // @[:@7040.4]
  input        io_backpressure // @[:@7040.4]
);
  wire [7:0] SRAMVerilogSim_rdata; // @[SRAM.scala 185:23:@7042.4]
  wire [7:0] SRAMVerilogSim_wdata; // @[SRAM.scala 185:23:@7042.4]
  wire  SRAMVerilogSim_backpressure; // @[SRAM.scala 185:23:@7042.4]
  wire  SRAMVerilogSim_wen; // @[SRAM.scala 185:23:@7042.4]
  wire  SRAMVerilogSim_waddrEn; // @[SRAM.scala 185:23:@7042.4]
  wire  SRAMVerilogSim_raddrEn; // @[SRAM.scala 185:23:@7042.4]
  wire [8:0] SRAMVerilogSim_waddr; // @[SRAM.scala 185:23:@7042.4]
  wire [8:0] SRAMVerilogSim_raddr; // @[SRAM.scala 185:23:@7042.4]
  wire  SRAMVerilogSim_clk; // @[SRAM.scala 185:23:@7042.4]
  SRAMVerilogSim #(.DWIDTH(8), .WORDS(480), .AWIDTH(9)) SRAMVerilogSim ( // @[SRAM.scala 185:23:@7042.4]
    .rdata(SRAMVerilogSim_rdata),
    .wdata(SRAMVerilogSim_wdata),
    .backpressure(SRAMVerilogSim_backpressure),
    .wen(SRAMVerilogSim_wen),
    .waddrEn(SRAMVerilogSim_waddrEn),
    .raddrEn(SRAMVerilogSim_raddrEn),
    .waddr(SRAMVerilogSim_waddr),
    .raddr(SRAMVerilogSim_raddr),
    .clk(SRAMVerilogSim_clk)
  );
  assign io_rdata = SRAMVerilogSim_rdata; // @[SRAM.scala 195:16:@7062.4]
  assign SRAMVerilogSim_wdata = io_wdata; // @[SRAM.scala 190:20:@7056.4]
  assign SRAMVerilogSim_backpressure = io_backpressure; // @[SRAM.scala 191:27:@7057.4]
  assign SRAMVerilogSim_wen = io_wen; // @[SRAM.scala 188:18:@7054.4]
  assign SRAMVerilogSim_waddrEn = 1'h1; // @[SRAM.scala 193:22:@7059.4]
  assign SRAMVerilogSim_raddrEn = 1'h1; // @[SRAM.scala 192:22:@7058.4]
  assign SRAMVerilogSim_waddr = io_waddr; // @[SRAM.scala 189:20:@7055.4]
  assign SRAMVerilogSim_raddr = io_raddr; // @[SRAM.scala 187:20:@7053.4]
  assign SRAMVerilogSim_clk = clock; // @[SRAM.scala 186:18:@7052.4]
endmodule
module RetimeWrapper_53( // @[:@7076.2]
  input        clock, // @[:@7077.4]
  input        reset, // @[:@7078.4]
  input        io_flow, // @[:@7079.4]
  input  [8:0] io_in, // @[:@7079.4]
  output [8:0] io_out // @[:@7079.4]
);
  wire [8:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@7081.4]
  wire [8:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@7081.4]
  wire [8:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@7081.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@7081.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@7081.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@7081.4]
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@7081.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@7094.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@7093.4]
  assign sr_init = 9'h0; // @[RetimeShiftRegister.scala 19:16:@7092.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@7091.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@7090.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@7088.4]
endmodule
module Mem1D_5( // @[:@7096.2]
  input        clock, // @[:@7097.4]
  input        reset, // @[:@7098.4]
  input  [8:0] io_r_ofs_0, // @[:@7099.4]
  input        io_r_backpressure, // @[:@7099.4]
  input  [8:0] io_w_ofs_0, // @[:@7099.4]
  input  [7:0] io_w_data_0, // @[:@7099.4]
  input        io_w_en_0, // @[:@7099.4]
  output [7:0] io_output // @[:@7099.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 705:21:@7103.4]
  wire [8:0] SRAM_io_raddr; // @[MemPrimitives.scala 705:21:@7103.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 705:21:@7103.4]
  wire [8:0] SRAM_io_waddr; // @[MemPrimitives.scala 705:21:@7103.4]
  wire [7:0] SRAM_io_wdata; // @[MemPrimitives.scala 705:21:@7103.4]
  wire [7:0] SRAM_io_rdata; // @[MemPrimitives.scala 705:21:@7103.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 705:21:@7103.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@7106.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@7106.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@7106.4]
  wire [8:0] RetimeWrapper_io_in; // @[package.scala 93:22:@7106.4]
  wire [8:0] RetimeWrapper_io_out; // @[package.scala 93:22:@7106.4]
  wire  wInBound; // @[MemPrimitives.scala 692:32:@7101.4]
  SRAM_1 SRAM ( // @[MemPrimitives.scala 705:21:@7103.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_53 RetimeWrapper ( // @[package.scala 93:22:@7106.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 9'h1e0; // @[MemPrimitives.scala 692:32:@7101.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 712:17:@7119.4]
  assign SRAM_clock = clock; // @[:@7104.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 706:37:@7113.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 709:22:@7116.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 708:22:@7114.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 710:22:@7117.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 711:30:@7118.4]
  assign RetimeWrapper_clock = clock; // @[:@7107.4]
  assign RetimeWrapper_reset = reset; // @[:@7108.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@7110.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@7109.4]
endmodule
module StickySelects_1( // @[:@8621.2]
  input   clock, // @[:@8622.4]
  input   reset, // @[:@8623.4]
  input   io_ins_0, // @[:@8624.4]
  input   io_ins_1, // @[:@8624.4]
  input   io_ins_2, // @[:@8624.4]
  input   io_ins_3, // @[:@8624.4]
  input   io_ins_4, // @[:@8624.4]
  input   io_ins_5, // @[:@8624.4]
  output  io_outs_0, // @[:@8624.4]
  output  io_outs_1, // @[:@8624.4]
  output  io_outs_2, // @[:@8624.4]
  output  io_outs_3, // @[:@8624.4]
  output  io_outs_4, // @[:@8624.4]
  output  io_outs_5 // @[:@8624.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@8626.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@8627.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@8628.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@8629.4]
  reg [31:0] _RAND_3;
  reg  _T_31; // @[StickySelects.scala 37:46:@8630.4]
  reg [31:0] _RAND_4;
  reg  _T_34; // @[StickySelects.scala 37:46:@8631.4]
  reg [31:0] _RAND_5;
  wire  _T_35; // @[StickySelects.scala 47:46:@8632.4]
  wire  _T_36; // @[StickySelects.scala 47:46:@8633.4]
  wire  _T_37; // @[StickySelects.scala 47:46:@8634.4]
  wire  _T_38; // @[StickySelects.scala 47:46:@8635.4]
  wire  _T_39; // @[StickySelects.scala 49:53:@8636.4]
  wire  _T_40; // @[StickySelects.scala 49:21:@8637.4]
  wire  _T_41; // @[StickySelects.scala 47:46:@8639.4]
  wire  _T_42; // @[StickySelects.scala 47:46:@8640.4]
  wire  _T_43; // @[StickySelects.scala 47:46:@8641.4]
  wire  _T_44; // @[StickySelects.scala 47:46:@8642.4]
  wire  _T_45; // @[StickySelects.scala 49:53:@8643.4]
  wire  _T_46; // @[StickySelects.scala 49:21:@8644.4]
  wire  _T_47; // @[StickySelects.scala 47:46:@8646.4]
  wire  _T_48; // @[StickySelects.scala 47:46:@8647.4]
  wire  _T_49; // @[StickySelects.scala 47:46:@8648.4]
  wire  _T_50; // @[StickySelects.scala 47:46:@8649.4]
  wire  _T_51; // @[StickySelects.scala 49:53:@8650.4]
  wire  _T_52; // @[StickySelects.scala 49:21:@8651.4]
  wire  _T_54; // @[StickySelects.scala 47:46:@8654.4]
  wire  _T_55; // @[StickySelects.scala 47:46:@8655.4]
  wire  _T_56; // @[StickySelects.scala 47:46:@8656.4]
  wire  _T_57; // @[StickySelects.scala 49:53:@8657.4]
  wire  _T_58; // @[StickySelects.scala 49:21:@8658.4]
  wire  _T_61; // @[StickySelects.scala 47:46:@8662.4]
  wire  _T_62; // @[StickySelects.scala 47:46:@8663.4]
  wire  _T_63; // @[StickySelects.scala 49:53:@8664.4]
  wire  _T_64; // @[StickySelects.scala 49:21:@8665.4]
  wire  _T_68; // @[StickySelects.scala 47:46:@8670.4]
  wire  _T_69; // @[StickySelects.scala 49:53:@8671.4]
  wire  _T_70; // @[StickySelects.scala 49:21:@8672.4]
  assign _T_35 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@8632.4]
  assign _T_36 = _T_35 | io_ins_3; // @[StickySelects.scala 47:46:@8633.4]
  assign _T_37 = _T_36 | io_ins_4; // @[StickySelects.scala 47:46:@8634.4]
  assign _T_38 = _T_37 | io_ins_5; // @[StickySelects.scala 47:46:@8635.4]
  assign _T_39 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@8636.4]
  assign _T_40 = _T_38 ? io_ins_0 : _T_39; // @[StickySelects.scala 49:21:@8637.4]
  assign _T_41 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@8639.4]
  assign _T_42 = _T_41 | io_ins_3; // @[StickySelects.scala 47:46:@8640.4]
  assign _T_43 = _T_42 | io_ins_4; // @[StickySelects.scala 47:46:@8641.4]
  assign _T_44 = _T_43 | io_ins_5; // @[StickySelects.scala 47:46:@8642.4]
  assign _T_45 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@8643.4]
  assign _T_46 = _T_44 ? io_ins_1 : _T_45; // @[StickySelects.scala 49:21:@8644.4]
  assign _T_47 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@8646.4]
  assign _T_48 = _T_47 | io_ins_3; // @[StickySelects.scala 47:46:@8647.4]
  assign _T_49 = _T_48 | io_ins_4; // @[StickySelects.scala 47:46:@8648.4]
  assign _T_50 = _T_49 | io_ins_5; // @[StickySelects.scala 47:46:@8649.4]
  assign _T_51 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@8650.4]
  assign _T_52 = _T_50 ? io_ins_2 : _T_51; // @[StickySelects.scala 49:21:@8651.4]
  assign _T_54 = _T_47 | io_ins_2; // @[StickySelects.scala 47:46:@8654.4]
  assign _T_55 = _T_54 | io_ins_4; // @[StickySelects.scala 47:46:@8655.4]
  assign _T_56 = _T_55 | io_ins_5; // @[StickySelects.scala 47:46:@8656.4]
  assign _T_57 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@8657.4]
  assign _T_58 = _T_56 ? io_ins_3 : _T_57; // @[StickySelects.scala 49:21:@8658.4]
  assign _T_61 = _T_54 | io_ins_3; // @[StickySelects.scala 47:46:@8662.4]
  assign _T_62 = _T_61 | io_ins_5; // @[StickySelects.scala 47:46:@8663.4]
  assign _T_63 = io_ins_4 | _T_31; // @[StickySelects.scala 49:53:@8664.4]
  assign _T_64 = _T_62 ? io_ins_4 : _T_63; // @[StickySelects.scala 49:21:@8665.4]
  assign _T_68 = _T_61 | io_ins_4; // @[StickySelects.scala 47:46:@8670.4]
  assign _T_69 = io_ins_5 | _T_34; // @[StickySelects.scala 49:53:@8671.4]
  assign _T_70 = _T_68 ? io_ins_5 : _T_69; // @[StickySelects.scala 49:21:@8672.4]
  assign io_outs_0 = _T_38 ? io_ins_0 : _T_39; // @[StickySelects.scala 53:57:@8674.4]
  assign io_outs_1 = _T_44 ? io_ins_1 : _T_45; // @[StickySelects.scala 53:57:@8675.4]
  assign io_outs_2 = _T_50 ? io_ins_2 : _T_51; // @[StickySelects.scala 53:57:@8676.4]
  assign io_outs_3 = _T_56 ? io_ins_3 : _T_57; // @[StickySelects.scala 53:57:@8677.4]
  assign io_outs_4 = _T_62 ? io_ins_4 : _T_63; // @[StickySelects.scala 53:57:@8678.4]
  assign io_outs_5 = _T_68 ? io_ins_5 : _T_69; // @[StickySelects.scala 53:57:@8679.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_31 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_38) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_39;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_44) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_45;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_50) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_51;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_56) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_57;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_62) begin
        _T_31 <= io_ins_4;
      end else begin
        _T_31 <= _T_63;
      end
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (_T_68) begin
        _T_34 <= io_ins_5;
      end else begin
        _T_34 <= _T_69;
      end
    end
  end
endmodule
module x385_lb_0( // @[:@12653.2]
  input        clock, // @[:@12654.4]
  input        reset, // @[:@12655.4]
  input  [2:0] io_rPort_11_banks_1, // @[:@12656.4]
  input  [2:0] io_rPort_11_banks_0, // @[:@12656.4]
  input  [8:0] io_rPort_11_ofs_0, // @[:@12656.4]
  input        io_rPort_11_en_0, // @[:@12656.4]
  input        io_rPort_11_backpressure, // @[:@12656.4]
  output [7:0] io_rPort_11_output_0, // @[:@12656.4]
  input  [2:0] io_rPort_10_banks_1, // @[:@12656.4]
  input  [2:0] io_rPort_10_banks_0, // @[:@12656.4]
  input  [8:0] io_rPort_10_ofs_0, // @[:@12656.4]
  input        io_rPort_10_en_0, // @[:@12656.4]
  input        io_rPort_10_backpressure, // @[:@12656.4]
  output [7:0] io_rPort_10_output_0, // @[:@12656.4]
  input  [2:0] io_rPort_9_banks_1, // @[:@12656.4]
  input  [2:0] io_rPort_9_banks_0, // @[:@12656.4]
  input  [8:0] io_rPort_9_ofs_0, // @[:@12656.4]
  input        io_rPort_9_en_0, // @[:@12656.4]
  input        io_rPort_9_backpressure, // @[:@12656.4]
  output [7:0] io_rPort_9_output_0, // @[:@12656.4]
  input  [2:0] io_rPort_8_banks_1, // @[:@12656.4]
  input  [2:0] io_rPort_8_banks_0, // @[:@12656.4]
  input  [8:0] io_rPort_8_ofs_0, // @[:@12656.4]
  input        io_rPort_8_en_0, // @[:@12656.4]
  input        io_rPort_8_backpressure, // @[:@12656.4]
  output [7:0] io_rPort_8_output_0, // @[:@12656.4]
  input  [2:0] io_rPort_7_banks_1, // @[:@12656.4]
  input  [2:0] io_rPort_7_banks_0, // @[:@12656.4]
  input  [8:0] io_rPort_7_ofs_0, // @[:@12656.4]
  input        io_rPort_7_en_0, // @[:@12656.4]
  input        io_rPort_7_backpressure, // @[:@12656.4]
  output [7:0] io_rPort_7_output_0, // @[:@12656.4]
  input  [2:0] io_rPort_6_banks_1, // @[:@12656.4]
  input  [2:0] io_rPort_6_banks_0, // @[:@12656.4]
  input  [8:0] io_rPort_6_ofs_0, // @[:@12656.4]
  input        io_rPort_6_en_0, // @[:@12656.4]
  input        io_rPort_6_backpressure, // @[:@12656.4]
  output [7:0] io_rPort_6_output_0, // @[:@12656.4]
  input  [2:0] io_rPort_5_banks_1, // @[:@12656.4]
  input  [2:0] io_rPort_5_banks_0, // @[:@12656.4]
  input  [8:0] io_rPort_5_ofs_0, // @[:@12656.4]
  input        io_rPort_5_en_0, // @[:@12656.4]
  input        io_rPort_5_backpressure, // @[:@12656.4]
  output [7:0] io_rPort_5_output_0, // @[:@12656.4]
  input  [2:0] io_rPort_4_banks_1, // @[:@12656.4]
  input  [2:0] io_rPort_4_banks_0, // @[:@12656.4]
  input  [8:0] io_rPort_4_ofs_0, // @[:@12656.4]
  input        io_rPort_4_en_0, // @[:@12656.4]
  input        io_rPort_4_backpressure, // @[:@12656.4]
  output [7:0] io_rPort_4_output_0, // @[:@12656.4]
  input  [2:0] io_rPort_3_banks_1, // @[:@12656.4]
  input  [2:0] io_rPort_3_banks_0, // @[:@12656.4]
  input  [8:0] io_rPort_3_ofs_0, // @[:@12656.4]
  input        io_rPort_3_en_0, // @[:@12656.4]
  input        io_rPort_3_backpressure, // @[:@12656.4]
  output [7:0] io_rPort_3_output_0, // @[:@12656.4]
  input  [2:0] io_rPort_2_banks_1, // @[:@12656.4]
  input  [2:0] io_rPort_2_banks_0, // @[:@12656.4]
  input  [8:0] io_rPort_2_ofs_0, // @[:@12656.4]
  input        io_rPort_2_en_0, // @[:@12656.4]
  input        io_rPort_2_backpressure, // @[:@12656.4]
  output [7:0] io_rPort_2_output_0, // @[:@12656.4]
  input  [2:0] io_rPort_1_banks_1, // @[:@12656.4]
  input  [2:0] io_rPort_1_banks_0, // @[:@12656.4]
  input  [8:0] io_rPort_1_ofs_0, // @[:@12656.4]
  input        io_rPort_1_en_0, // @[:@12656.4]
  input        io_rPort_1_backpressure, // @[:@12656.4]
  output [7:0] io_rPort_1_output_0, // @[:@12656.4]
  input  [2:0] io_rPort_0_banks_1, // @[:@12656.4]
  input  [2:0] io_rPort_0_banks_0, // @[:@12656.4]
  input  [8:0] io_rPort_0_ofs_0, // @[:@12656.4]
  input        io_rPort_0_en_0, // @[:@12656.4]
  input        io_rPort_0_backpressure, // @[:@12656.4]
  output [7:0] io_rPort_0_output_0, // @[:@12656.4]
  input  [2:0] io_wPort_1_banks_1, // @[:@12656.4]
  input  [2:0] io_wPort_1_banks_0, // @[:@12656.4]
  input  [8:0] io_wPort_1_ofs_0, // @[:@12656.4]
  input  [7:0] io_wPort_1_data_0, // @[:@12656.4]
  input        io_wPort_1_en_0, // @[:@12656.4]
  input  [2:0] io_wPort_0_banks_1, // @[:@12656.4]
  input  [2:0] io_wPort_0_banks_0, // @[:@12656.4]
  input  [8:0] io_wPort_0_ofs_0, // @[:@12656.4]
  input  [7:0] io_wPort_0_data_0, // @[:@12656.4]
  input        io_wPort_0_en_0 // @[:@12656.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@12747.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@12747.4]
  wire [8:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12747.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12747.4]
  wire [8:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12747.4]
  wire [7:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@12747.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@12747.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@12747.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@12763.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@12763.4]
  wire [8:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12763.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12763.4]
  wire [8:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12763.4]
  wire [7:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@12763.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@12763.4]
  wire [7:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@12763.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@12779.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@12779.4]
  wire [8:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12779.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12779.4]
  wire [8:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12779.4]
  wire [7:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@12779.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@12779.4]
  wire [7:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@12779.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@12795.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@12795.4]
  wire [8:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12795.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12795.4]
  wire [8:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12795.4]
  wire [7:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@12795.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@12795.4]
  wire [7:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@12795.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@12811.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@12811.4]
  wire [8:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12811.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12811.4]
  wire [8:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12811.4]
  wire [7:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@12811.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@12811.4]
  wire [7:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@12811.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@12827.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@12827.4]
  wire [8:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12827.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12827.4]
  wire [8:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12827.4]
  wire [7:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@12827.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@12827.4]
  wire [7:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@12827.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@12843.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@12843.4]
  wire [8:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12843.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12843.4]
  wire [8:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12843.4]
  wire [7:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@12843.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@12843.4]
  wire [7:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@12843.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@12859.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@12859.4]
  wire [8:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12859.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12859.4]
  wire [8:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12859.4]
  wire [7:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@12859.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@12859.4]
  wire [7:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@12859.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@12875.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@12875.4]
  wire [8:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12875.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12875.4]
  wire [8:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12875.4]
  wire [7:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@12875.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@12875.4]
  wire [7:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@12875.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@12891.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@12891.4]
  wire [8:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12891.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12891.4]
  wire [8:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12891.4]
  wire [7:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@12891.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@12891.4]
  wire [7:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@12891.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@12907.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@12907.4]
  wire [8:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12907.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12907.4]
  wire [8:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12907.4]
  wire [7:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@12907.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@12907.4]
  wire [7:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@12907.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@12923.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@12923.4]
  wire [8:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12923.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12923.4]
  wire [8:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12923.4]
  wire [7:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@12923.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@12923.4]
  wire [7:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@12923.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@12939.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@12939.4]
  wire [8:0] Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12939.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12939.4]
  wire [8:0] Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12939.4]
  wire [7:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@12939.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@12939.4]
  wire [7:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@12939.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@12955.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@12955.4]
  wire [8:0] Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12955.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12955.4]
  wire [8:0] Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12955.4]
  wire [7:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@12955.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@12955.4]
  wire [7:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@12955.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@12971.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@12971.4]
  wire [8:0] Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12971.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12971.4]
  wire [8:0] Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12971.4]
  wire [7:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@12971.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@12971.4]
  wire [7:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@12971.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@12987.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@12987.4]
  wire [8:0] Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12987.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12987.4]
  wire [8:0] Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12987.4]
  wire [7:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@12987.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@12987.4]
  wire [7:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@12987.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 121:29:@13219.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 121:29:@13219.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@13219.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 121:29:@13219.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 121:29:@13219.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 121:29:@13219.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 121:29:@13219.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 121:29:@13219.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@13219.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 121:29:@13219.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 121:29:@13219.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 121:29:@13219.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 121:29:@13219.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 121:29:@13219.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 121:29:@13281.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 121:29:@13281.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@13281.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 121:29:@13281.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 121:29:@13281.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 121:29:@13281.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 121:29:@13281.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 121:29:@13281.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@13281.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 121:29:@13281.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 121:29:@13281.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 121:29:@13281.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 121:29:@13281.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 121:29:@13281.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 121:29:@13343.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 121:29:@13343.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@13343.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 121:29:@13343.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 121:29:@13343.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 121:29:@13343.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 121:29:@13343.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 121:29:@13343.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@13343.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 121:29:@13343.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 121:29:@13343.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 121:29:@13343.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 121:29:@13343.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 121:29:@13343.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 121:29:@13405.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 121:29:@13405.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@13405.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 121:29:@13405.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 121:29:@13405.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 121:29:@13405.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 121:29:@13405.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 121:29:@13405.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@13405.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 121:29:@13405.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 121:29:@13405.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 121:29:@13405.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 121:29:@13405.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 121:29:@13405.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 121:29:@13467.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 121:29:@13467.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@13467.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 121:29:@13467.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 121:29:@13467.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 121:29:@13467.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 121:29:@13467.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 121:29:@13467.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@13467.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 121:29:@13467.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 121:29:@13467.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 121:29:@13467.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 121:29:@13467.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 121:29:@13467.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 121:29:@13529.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 121:29:@13529.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@13529.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 121:29:@13529.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 121:29:@13529.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 121:29:@13529.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 121:29:@13529.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 121:29:@13529.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@13529.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 121:29:@13529.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 121:29:@13529.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 121:29:@13529.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 121:29:@13529.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 121:29:@13529.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 121:29:@13591.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 121:29:@13591.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@13591.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 121:29:@13591.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 121:29:@13591.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 121:29:@13591.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 121:29:@13591.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 121:29:@13591.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@13591.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 121:29:@13591.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 121:29:@13591.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 121:29:@13591.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 121:29:@13591.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 121:29:@13591.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 121:29:@13653.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 121:29:@13653.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@13653.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 121:29:@13653.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 121:29:@13653.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 121:29:@13653.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 121:29:@13653.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 121:29:@13653.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@13653.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 121:29:@13653.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 121:29:@13653.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 121:29:@13653.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 121:29:@13653.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 121:29:@13653.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 121:29:@13715.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 121:29:@13777.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 121:29:@13777.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@13777.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 121:29:@13777.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 121:29:@13777.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 121:29:@13777.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 121:29:@13777.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 121:29:@13777.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@13777.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 121:29:@13777.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 121:29:@13777.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 121:29:@13777.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 121:29:@13777.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 121:29:@13777.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 121:29:@13839.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 121:29:@13839.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@13839.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 121:29:@13839.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 121:29:@13839.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 121:29:@13839.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 121:29:@13839.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 121:29:@13839.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@13839.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 121:29:@13839.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 121:29:@13839.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 121:29:@13839.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 121:29:@13839.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 121:29:@13839.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 121:29:@13901.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 121:29:@13901.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@13901.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 121:29:@13901.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 121:29:@13901.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 121:29:@13901.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 121:29:@13901.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 121:29:@13901.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@13901.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 121:29:@13901.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 121:29:@13901.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 121:29:@13901.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 121:29:@13901.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 121:29:@13901.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_12_io_ins_4; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_12_io_ins_5; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_12_io_outs_4; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_12_io_outs_5; // @[MemPrimitives.scala 121:29:@13963.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 121:29:@14025.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 121:29:@14025.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 121:29:@14025.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 121:29:@14025.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 121:29:@14025.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 121:29:@14025.4]
  wire  StickySelects_13_io_ins_4; // @[MemPrimitives.scala 121:29:@14025.4]
  wire  StickySelects_13_io_ins_5; // @[MemPrimitives.scala 121:29:@14025.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 121:29:@14025.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 121:29:@14025.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 121:29:@14025.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 121:29:@14025.4]
  wire  StickySelects_13_io_outs_4; // @[MemPrimitives.scala 121:29:@14025.4]
  wire  StickySelects_13_io_outs_5; // @[MemPrimitives.scala 121:29:@14025.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 121:29:@14087.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 121:29:@14087.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 121:29:@14087.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 121:29:@14087.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 121:29:@14087.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 121:29:@14087.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 121:29:@14087.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 121:29:@14087.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 121:29:@14087.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 121:29:@14087.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 121:29:@14087.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 121:29:@14087.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 121:29:@14087.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 121:29:@14087.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 121:29:@14149.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 121:29:@14149.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 121:29:@14149.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 121:29:@14149.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 121:29:@14149.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 121:29:@14149.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 121:29:@14149.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 121:29:@14149.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 121:29:@14149.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 121:29:@14149.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 121:29:@14149.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 121:29:@14149.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 121:29:@14149.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 121:29:@14149.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@14212.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@14212.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@14212.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@14212.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@14212.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@14220.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@14220.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@14220.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@14220.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@14220.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@14228.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@14228.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@14228.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@14228.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@14228.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@14236.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@14236.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@14236.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@14236.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@14236.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@14244.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@14244.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@14244.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@14244.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@14244.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@14252.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@14252.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@14252.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@14252.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@14252.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@14260.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@14260.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@14260.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@14260.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@14260.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@14268.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@14268.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@14268.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@14268.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@14268.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@14308.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@14308.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@14308.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@14308.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@14308.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@14316.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@14316.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@14316.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@14316.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@14316.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@14324.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@14324.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@14324.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@14324.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@14324.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@14332.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@14332.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@14332.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@14332.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@14332.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@14340.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@14340.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@14340.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@14340.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@14340.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@14348.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@14348.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@14348.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@14348.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@14348.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@14356.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@14356.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@14356.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@14356.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@14356.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@14364.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@14364.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@14364.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@14364.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@14364.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@14404.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@14404.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@14404.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@14404.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@14404.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@14412.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@14412.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@14412.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@14412.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@14412.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@14420.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@14420.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@14420.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@14420.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@14420.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@14428.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@14428.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@14428.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@14428.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@14428.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@14436.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@14436.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@14436.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@14436.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@14436.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@14444.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@14444.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@14444.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@14444.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@14444.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@14452.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@14452.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@14452.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@14452.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@14452.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@14460.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@14460.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@14460.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@14460.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@14460.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@14500.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@14500.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@14500.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@14500.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@14500.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@14508.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@14508.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@14508.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@14508.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@14508.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@14516.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@14516.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@14516.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@14516.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@14516.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@14524.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@14524.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@14524.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@14524.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@14524.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@14532.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@14532.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@14532.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@14532.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@14532.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@14540.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@14540.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@14540.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@14540.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@14540.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@14548.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@14548.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@14548.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@14548.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@14548.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@14556.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@14556.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@14556.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@14556.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@14556.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@14596.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@14596.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@14596.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@14596.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@14596.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@14604.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@14604.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@14604.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@14604.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@14604.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@14612.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@14612.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@14612.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@14612.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@14612.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@14620.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@14620.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@14620.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@14620.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@14620.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@14628.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@14628.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@14628.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@14628.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@14628.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@14636.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@14636.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@14636.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@14636.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@14636.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@14644.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@14644.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@14644.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@14644.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@14644.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@14652.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@14652.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@14652.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@14652.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@14652.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@14692.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@14692.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@14692.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@14692.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@14692.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@14700.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@14700.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@14700.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@14700.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@14700.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@14708.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@14708.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@14708.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@14708.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@14708.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@14716.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@14716.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@14716.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@14716.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@14716.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@14724.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@14724.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@14724.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@14724.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@14724.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@14732.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@14732.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@14732.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@14732.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@14732.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@14740.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@14740.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@14740.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@14740.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@14740.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@14748.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@14748.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@14748.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@14748.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@14748.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@14788.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@14788.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@14788.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@14788.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@14788.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@14796.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@14796.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@14796.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@14796.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@14796.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@14804.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@14804.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@14804.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@14804.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@14804.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@14812.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@14812.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@14812.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@14812.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@14812.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@14820.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@14820.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@14820.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@14820.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@14820.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@14828.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@14828.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@14828.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@14828.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@14828.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@14836.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@14836.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@14836.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@14836.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@14836.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@14844.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@14844.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@14844.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@14844.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@14844.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@14884.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@14884.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@14884.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@14884.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@14884.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@14892.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@14892.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@14892.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@14892.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@14892.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@14900.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@14900.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@14900.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@14900.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@14900.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@14908.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@14908.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@14908.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@14908.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@14908.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@14916.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@14916.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@14916.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@14916.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@14916.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@14924.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@14924.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@14924.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@14924.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@14924.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@14932.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@14932.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@14932.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@14932.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@14932.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@14940.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@14940.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@14940.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@14940.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@14940.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@14980.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@14980.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@14980.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@14980.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@14980.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@14988.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@14988.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@14988.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@14988.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@14988.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@14996.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@14996.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@14996.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@14996.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@14996.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@15004.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@15004.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@15004.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@15004.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@15004.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@15012.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@15012.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@15012.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@15012.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@15012.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@15020.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@15020.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@15020.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@15020.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@15020.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@15028.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@15028.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@15028.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@15028.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@15028.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@15036.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@15036.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@15036.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@15036.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@15036.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@15076.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@15076.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@15076.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@15076.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@15076.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@15084.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@15084.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@15084.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@15084.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@15084.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@15092.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@15092.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@15092.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@15092.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@15092.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@15100.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@15100.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@15100.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@15100.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@15100.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@15108.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@15108.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@15108.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@15108.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@15108.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@15116.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@15116.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@15116.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@15116.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@15116.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@15124.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@15124.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@15124.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@15124.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@15124.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@15132.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@15132.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@15132.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@15132.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@15132.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@15172.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@15172.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@15172.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@15172.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@15172.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@15180.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@15180.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@15180.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@15180.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@15180.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@15188.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@15188.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@15188.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@15188.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@15188.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@15196.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@15196.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@15196.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@15196.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@15196.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@15204.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@15204.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@15204.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@15204.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@15204.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@15212.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@15212.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@15212.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@15212.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@15212.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@15220.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@15220.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@15220.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@15220.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@15220.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@15228.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@15228.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@15228.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@15228.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@15228.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@15268.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@15268.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@15268.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@15268.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@15268.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@15276.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@15276.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@15276.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@15276.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@15276.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@15284.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@15284.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@15284.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@15284.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@15284.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@15292.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@15292.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@15292.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@15292.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@15292.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@15300.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@15300.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@15300.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@15300.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@15300.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@15308.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@15308.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@15308.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@15308.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@15308.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@15316.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@15316.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@15316.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@15316.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@15316.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@15324.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@15324.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@15324.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@15324.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@15324.4]
  wire  _T_444; // @[MemPrimitives.scala 82:210:@13003.4]
  wire  _T_446; // @[MemPrimitives.scala 82:210:@13004.4]
  wire  _T_447; // @[MemPrimitives.scala 82:228:@13005.4]
  wire  _T_448; // @[MemPrimitives.scala 83:102:@13006.4]
  wire [17:0] _T_450; // @[Cat.scala 30:58:@13008.4]
  wire  _T_455; // @[MemPrimitives.scala 82:210:@13015.4]
  wire  _T_457; // @[MemPrimitives.scala 82:210:@13016.4]
  wire  _T_458; // @[MemPrimitives.scala 82:228:@13017.4]
  wire  _T_459; // @[MemPrimitives.scala 83:102:@13018.4]
  wire [17:0] _T_461; // @[Cat.scala 30:58:@13020.4]
  wire  _T_468; // @[MemPrimitives.scala 82:210:@13028.4]
  wire  _T_469; // @[MemPrimitives.scala 82:228:@13029.4]
  wire  _T_470; // @[MemPrimitives.scala 83:102:@13030.4]
  wire [17:0] _T_472; // @[Cat.scala 30:58:@13032.4]
  wire  _T_479; // @[MemPrimitives.scala 82:210:@13040.4]
  wire  _T_480; // @[MemPrimitives.scala 82:228:@13041.4]
  wire  _T_481; // @[MemPrimitives.scala 83:102:@13042.4]
  wire [17:0] _T_483; // @[Cat.scala 30:58:@13044.4]
  wire  _T_488; // @[MemPrimitives.scala 82:210:@13051.4]
  wire  _T_491; // @[MemPrimitives.scala 82:228:@13053.4]
  wire  _T_492; // @[MemPrimitives.scala 83:102:@13054.4]
  wire [17:0] _T_494; // @[Cat.scala 30:58:@13056.4]
  wire  _T_499; // @[MemPrimitives.scala 82:210:@13063.4]
  wire  _T_502; // @[MemPrimitives.scala 82:228:@13065.4]
  wire  _T_503; // @[MemPrimitives.scala 83:102:@13066.4]
  wire [17:0] _T_505; // @[Cat.scala 30:58:@13068.4]
  wire  _T_513; // @[MemPrimitives.scala 82:228:@13077.4]
  wire  _T_514; // @[MemPrimitives.scala 83:102:@13078.4]
  wire [17:0] _T_516; // @[Cat.scala 30:58:@13080.4]
  wire  _T_524; // @[MemPrimitives.scala 82:228:@13089.4]
  wire  _T_525; // @[MemPrimitives.scala 83:102:@13090.4]
  wire [17:0] _T_527; // @[Cat.scala 30:58:@13092.4]
  wire  _T_532; // @[MemPrimitives.scala 82:210:@13099.4]
  wire  _T_535; // @[MemPrimitives.scala 82:228:@13101.4]
  wire  _T_536; // @[MemPrimitives.scala 83:102:@13102.4]
  wire [17:0] _T_538; // @[Cat.scala 30:58:@13104.4]
  wire  _T_543; // @[MemPrimitives.scala 82:210:@13111.4]
  wire  _T_546; // @[MemPrimitives.scala 82:228:@13113.4]
  wire  _T_547; // @[MemPrimitives.scala 83:102:@13114.4]
  wire [17:0] _T_549; // @[Cat.scala 30:58:@13116.4]
  wire  _T_557; // @[MemPrimitives.scala 82:228:@13125.4]
  wire  _T_558; // @[MemPrimitives.scala 83:102:@13126.4]
  wire [17:0] _T_560; // @[Cat.scala 30:58:@13128.4]
  wire  _T_568; // @[MemPrimitives.scala 82:228:@13137.4]
  wire  _T_569; // @[MemPrimitives.scala 83:102:@13138.4]
  wire [17:0] _T_571; // @[Cat.scala 30:58:@13140.4]
  wire  _T_576; // @[MemPrimitives.scala 82:210:@13147.4]
  wire  _T_579; // @[MemPrimitives.scala 82:228:@13149.4]
  wire  _T_580; // @[MemPrimitives.scala 83:102:@13150.4]
  wire [17:0] _T_582; // @[Cat.scala 30:58:@13152.4]
  wire  _T_587; // @[MemPrimitives.scala 82:210:@13159.4]
  wire  _T_590; // @[MemPrimitives.scala 82:228:@13161.4]
  wire  _T_591; // @[MemPrimitives.scala 83:102:@13162.4]
  wire [17:0] _T_593; // @[Cat.scala 30:58:@13164.4]
  wire  _T_601; // @[MemPrimitives.scala 82:228:@13173.4]
  wire  _T_602; // @[MemPrimitives.scala 83:102:@13174.4]
  wire [17:0] _T_604; // @[Cat.scala 30:58:@13176.4]
  wire  _T_612; // @[MemPrimitives.scala 82:228:@13185.4]
  wire  _T_613; // @[MemPrimitives.scala 83:102:@13186.4]
  wire [17:0] _T_615; // @[Cat.scala 30:58:@13188.4]
  wire  _T_620; // @[MemPrimitives.scala 110:210:@13195.4]
  wire  _T_622; // @[MemPrimitives.scala 110:210:@13196.4]
  wire  _T_623; // @[MemPrimitives.scala 110:228:@13197.4]
  wire  _T_626; // @[MemPrimitives.scala 110:210:@13199.4]
  wire  _T_628; // @[MemPrimitives.scala 110:210:@13200.4]
  wire  _T_629; // @[MemPrimitives.scala 110:228:@13201.4]
  wire  _T_632; // @[MemPrimitives.scala 110:210:@13203.4]
  wire  _T_634; // @[MemPrimitives.scala 110:210:@13204.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@13205.4]
  wire  _T_638; // @[MemPrimitives.scala 110:210:@13207.4]
  wire  _T_640; // @[MemPrimitives.scala 110:210:@13208.4]
  wire  _T_641; // @[MemPrimitives.scala 110:228:@13209.4]
  wire  _T_644; // @[MemPrimitives.scala 110:210:@13211.4]
  wire  _T_646; // @[MemPrimitives.scala 110:210:@13212.4]
  wire  _T_647; // @[MemPrimitives.scala 110:228:@13213.4]
  wire  _T_650; // @[MemPrimitives.scala 110:210:@13215.4]
  wire  _T_652; // @[MemPrimitives.scala 110:210:@13216.4]
  wire  _T_653; // @[MemPrimitives.scala 110:228:@13217.4]
  wire  _T_655; // @[MemPrimitives.scala 123:41:@13228.4]
  wire  _T_656; // @[MemPrimitives.scala 123:41:@13229.4]
  wire  _T_657; // @[MemPrimitives.scala 123:41:@13230.4]
  wire  _T_658; // @[MemPrimitives.scala 123:41:@13231.4]
  wire  _T_659; // @[MemPrimitives.scala 123:41:@13232.4]
  wire  _T_660; // @[MemPrimitives.scala 123:41:@13233.4]
  wire [10:0] _T_662; // @[Cat.scala 30:58:@13235.4]
  wire [10:0] _T_664; // @[Cat.scala 30:58:@13237.4]
  wire [10:0] _T_666; // @[Cat.scala 30:58:@13239.4]
  wire [10:0] _T_668; // @[Cat.scala 30:58:@13241.4]
  wire [10:0] _T_670; // @[Cat.scala 30:58:@13243.4]
  wire [10:0] _T_672; // @[Cat.scala 30:58:@13245.4]
  wire [10:0] _T_673; // @[Mux.scala 31:69:@13246.4]
  wire [10:0] _T_674; // @[Mux.scala 31:69:@13247.4]
  wire [10:0] _T_675; // @[Mux.scala 31:69:@13248.4]
  wire [10:0] _T_676; // @[Mux.scala 31:69:@13249.4]
  wire [10:0] _T_677; // @[Mux.scala 31:69:@13250.4]
  wire  _T_682; // @[MemPrimitives.scala 110:210:@13257.4]
  wire  _T_684; // @[MemPrimitives.scala 110:210:@13258.4]
  wire  _T_685; // @[MemPrimitives.scala 110:228:@13259.4]
  wire  _T_688; // @[MemPrimitives.scala 110:210:@13261.4]
  wire  _T_690; // @[MemPrimitives.scala 110:210:@13262.4]
  wire  _T_691; // @[MemPrimitives.scala 110:228:@13263.4]
  wire  _T_694; // @[MemPrimitives.scala 110:210:@13265.4]
  wire  _T_696; // @[MemPrimitives.scala 110:210:@13266.4]
  wire  _T_697; // @[MemPrimitives.scala 110:228:@13267.4]
  wire  _T_700; // @[MemPrimitives.scala 110:210:@13269.4]
  wire  _T_702; // @[MemPrimitives.scala 110:210:@13270.4]
  wire  _T_703; // @[MemPrimitives.scala 110:228:@13271.4]
  wire  _T_706; // @[MemPrimitives.scala 110:210:@13273.4]
  wire  _T_708; // @[MemPrimitives.scala 110:210:@13274.4]
  wire  _T_709; // @[MemPrimitives.scala 110:228:@13275.4]
  wire  _T_712; // @[MemPrimitives.scala 110:210:@13277.4]
  wire  _T_714; // @[MemPrimitives.scala 110:210:@13278.4]
  wire  _T_715; // @[MemPrimitives.scala 110:228:@13279.4]
  wire  _T_717; // @[MemPrimitives.scala 123:41:@13290.4]
  wire  _T_718; // @[MemPrimitives.scala 123:41:@13291.4]
  wire  _T_719; // @[MemPrimitives.scala 123:41:@13292.4]
  wire  _T_720; // @[MemPrimitives.scala 123:41:@13293.4]
  wire  _T_721; // @[MemPrimitives.scala 123:41:@13294.4]
  wire  _T_722; // @[MemPrimitives.scala 123:41:@13295.4]
  wire [10:0] _T_724; // @[Cat.scala 30:58:@13297.4]
  wire [10:0] _T_726; // @[Cat.scala 30:58:@13299.4]
  wire [10:0] _T_728; // @[Cat.scala 30:58:@13301.4]
  wire [10:0] _T_730; // @[Cat.scala 30:58:@13303.4]
  wire [10:0] _T_732; // @[Cat.scala 30:58:@13305.4]
  wire [10:0] _T_734; // @[Cat.scala 30:58:@13307.4]
  wire [10:0] _T_735; // @[Mux.scala 31:69:@13308.4]
  wire [10:0] _T_736; // @[Mux.scala 31:69:@13309.4]
  wire [10:0] _T_737; // @[Mux.scala 31:69:@13310.4]
  wire [10:0] _T_738; // @[Mux.scala 31:69:@13311.4]
  wire [10:0] _T_739; // @[Mux.scala 31:69:@13312.4]
  wire  _T_746; // @[MemPrimitives.scala 110:210:@13320.4]
  wire  _T_747; // @[MemPrimitives.scala 110:228:@13321.4]
  wire  _T_752; // @[MemPrimitives.scala 110:210:@13324.4]
  wire  _T_753; // @[MemPrimitives.scala 110:228:@13325.4]
  wire  _T_758; // @[MemPrimitives.scala 110:210:@13328.4]
  wire  _T_759; // @[MemPrimitives.scala 110:228:@13329.4]
  wire  _T_764; // @[MemPrimitives.scala 110:210:@13332.4]
  wire  _T_765; // @[MemPrimitives.scala 110:228:@13333.4]
  wire  _T_770; // @[MemPrimitives.scala 110:210:@13336.4]
  wire  _T_771; // @[MemPrimitives.scala 110:228:@13337.4]
  wire  _T_776; // @[MemPrimitives.scala 110:210:@13340.4]
  wire  _T_777; // @[MemPrimitives.scala 110:228:@13341.4]
  wire  _T_779; // @[MemPrimitives.scala 123:41:@13352.4]
  wire  _T_780; // @[MemPrimitives.scala 123:41:@13353.4]
  wire  _T_781; // @[MemPrimitives.scala 123:41:@13354.4]
  wire  _T_782; // @[MemPrimitives.scala 123:41:@13355.4]
  wire  _T_783; // @[MemPrimitives.scala 123:41:@13356.4]
  wire  _T_784; // @[MemPrimitives.scala 123:41:@13357.4]
  wire [10:0] _T_786; // @[Cat.scala 30:58:@13359.4]
  wire [10:0] _T_788; // @[Cat.scala 30:58:@13361.4]
  wire [10:0] _T_790; // @[Cat.scala 30:58:@13363.4]
  wire [10:0] _T_792; // @[Cat.scala 30:58:@13365.4]
  wire [10:0] _T_794; // @[Cat.scala 30:58:@13367.4]
  wire [10:0] _T_796; // @[Cat.scala 30:58:@13369.4]
  wire [10:0] _T_797; // @[Mux.scala 31:69:@13370.4]
  wire [10:0] _T_798; // @[Mux.scala 31:69:@13371.4]
  wire [10:0] _T_799; // @[Mux.scala 31:69:@13372.4]
  wire [10:0] _T_800; // @[Mux.scala 31:69:@13373.4]
  wire [10:0] _T_801; // @[Mux.scala 31:69:@13374.4]
  wire  _T_808; // @[MemPrimitives.scala 110:210:@13382.4]
  wire  _T_809; // @[MemPrimitives.scala 110:228:@13383.4]
  wire  _T_814; // @[MemPrimitives.scala 110:210:@13386.4]
  wire  _T_815; // @[MemPrimitives.scala 110:228:@13387.4]
  wire  _T_820; // @[MemPrimitives.scala 110:210:@13390.4]
  wire  _T_821; // @[MemPrimitives.scala 110:228:@13391.4]
  wire  _T_826; // @[MemPrimitives.scala 110:210:@13394.4]
  wire  _T_827; // @[MemPrimitives.scala 110:228:@13395.4]
  wire  _T_832; // @[MemPrimitives.scala 110:210:@13398.4]
  wire  _T_833; // @[MemPrimitives.scala 110:228:@13399.4]
  wire  _T_838; // @[MemPrimitives.scala 110:210:@13402.4]
  wire  _T_839; // @[MemPrimitives.scala 110:228:@13403.4]
  wire  _T_841; // @[MemPrimitives.scala 123:41:@13414.4]
  wire  _T_842; // @[MemPrimitives.scala 123:41:@13415.4]
  wire  _T_843; // @[MemPrimitives.scala 123:41:@13416.4]
  wire  _T_844; // @[MemPrimitives.scala 123:41:@13417.4]
  wire  _T_845; // @[MemPrimitives.scala 123:41:@13418.4]
  wire  _T_846; // @[MemPrimitives.scala 123:41:@13419.4]
  wire [10:0] _T_848; // @[Cat.scala 30:58:@13421.4]
  wire [10:0] _T_850; // @[Cat.scala 30:58:@13423.4]
  wire [10:0] _T_852; // @[Cat.scala 30:58:@13425.4]
  wire [10:0] _T_854; // @[Cat.scala 30:58:@13427.4]
  wire [10:0] _T_856; // @[Cat.scala 30:58:@13429.4]
  wire [10:0] _T_858; // @[Cat.scala 30:58:@13431.4]
  wire [10:0] _T_859; // @[Mux.scala 31:69:@13432.4]
  wire [10:0] _T_860; // @[Mux.scala 31:69:@13433.4]
  wire [10:0] _T_861; // @[Mux.scala 31:69:@13434.4]
  wire [10:0] _T_862; // @[Mux.scala 31:69:@13435.4]
  wire [10:0] _T_863; // @[Mux.scala 31:69:@13436.4]
  wire  _T_868; // @[MemPrimitives.scala 110:210:@13443.4]
  wire  _T_871; // @[MemPrimitives.scala 110:228:@13445.4]
  wire  _T_874; // @[MemPrimitives.scala 110:210:@13447.4]
  wire  _T_877; // @[MemPrimitives.scala 110:228:@13449.4]
  wire  _T_880; // @[MemPrimitives.scala 110:210:@13451.4]
  wire  _T_883; // @[MemPrimitives.scala 110:228:@13453.4]
  wire  _T_886; // @[MemPrimitives.scala 110:210:@13455.4]
  wire  _T_889; // @[MemPrimitives.scala 110:228:@13457.4]
  wire  _T_892; // @[MemPrimitives.scala 110:210:@13459.4]
  wire  _T_895; // @[MemPrimitives.scala 110:228:@13461.4]
  wire  _T_898; // @[MemPrimitives.scala 110:210:@13463.4]
  wire  _T_901; // @[MemPrimitives.scala 110:228:@13465.4]
  wire  _T_903; // @[MemPrimitives.scala 123:41:@13476.4]
  wire  _T_904; // @[MemPrimitives.scala 123:41:@13477.4]
  wire  _T_905; // @[MemPrimitives.scala 123:41:@13478.4]
  wire  _T_906; // @[MemPrimitives.scala 123:41:@13479.4]
  wire  _T_907; // @[MemPrimitives.scala 123:41:@13480.4]
  wire  _T_908; // @[MemPrimitives.scala 123:41:@13481.4]
  wire [10:0] _T_910; // @[Cat.scala 30:58:@13483.4]
  wire [10:0] _T_912; // @[Cat.scala 30:58:@13485.4]
  wire [10:0] _T_914; // @[Cat.scala 30:58:@13487.4]
  wire [10:0] _T_916; // @[Cat.scala 30:58:@13489.4]
  wire [10:0] _T_918; // @[Cat.scala 30:58:@13491.4]
  wire [10:0] _T_920; // @[Cat.scala 30:58:@13493.4]
  wire [10:0] _T_921; // @[Mux.scala 31:69:@13494.4]
  wire [10:0] _T_922; // @[Mux.scala 31:69:@13495.4]
  wire [10:0] _T_923; // @[Mux.scala 31:69:@13496.4]
  wire [10:0] _T_924; // @[Mux.scala 31:69:@13497.4]
  wire [10:0] _T_925; // @[Mux.scala 31:69:@13498.4]
  wire  _T_930; // @[MemPrimitives.scala 110:210:@13505.4]
  wire  _T_933; // @[MemPrimitives.scala 110:228:@13507.4]
  wire  _T_936; // @[MemPrimitives.scala 110:210:@13509.4]
  wire  _T_939; // @[MemPrimitives.scala 110:228:@13511.4]
  wire  _T_942; // @[MemPrimitives.scala 110:210:@13513.4]
  wire  _T_945; // @[MemPrimitives.scala 110:228:@13515.4]
  wire  _T_948; // @[MemPrimitives.scala 110:210:@13517.4]
  wire  _T_951; // @[MemPrimitives.scala 110:228:@13519.4]
  wire  _T_954; // @[MemPrimitives.scala 110:210:@13521.4]
  wire  _T_957; // @[MemPrimitives.scala 110:228:@13523.4]
  wire  _T_960; // @[MemPrimitives.scala 110:210:@13525.4]
  wire  _T_963; // @[MemPrimitives.scala 110:228:@13527.4]
  wire  _T_965; // @[MemPrimitives.scala 123:41:@13538.4]
  wire  _T_966; // @[MemPrimitives.scala 123:41:@13539.4]
  wire  _T_967; // @[MemPrimitives.scala 123:41:@13540.4]
  wire  _T_968; // @[MemPrimitives.scala 123:41:@13541.4]
  wire  _T_969; // @[MemPrimitives.scala 123:41:@13542.4]
  wire  _T_970; // @[MemPrimitives.scala 123:41:@13543.4]
  wire [10:0] _T_972; // @[Cat.scala 30:58:@13545.4]
  wire [10:0] _T_974; // @[Cat.scala 30:58:@13547.4]
  wire [10:0] _T_976; // @[Cat.scala 30:58:@13549.4]
  wire [10:0] _T_978; // @[Cat.scala 30:58:@13551.4]
  wire [10:0] _T_980; // @[Cat.scala 30:58:@13553.4]
  wire [10:0] _T_982; // @[Cat.scala 30:58:@13555.4]
  wire [10:0] _T_983; // @[Mux.scala 31:69:@13556.4]
  wire [10:0] _T_984; // @[Mux.scala 31:69:@13557.4]
  wire [10:0] _T_985; // @[Mux.scala 31:69:@13558.4]
  wire [10:0] _T_986; // @[Mux.scala 31:69:@13559.4]
  wire [10:0] _T_987; // @[Mux.scala 31:69:@13560.4]
  wire  _T_995; // @[MemPrimitives.scala 110:228:@13569.4]
  wire  _T_1001; // @[MemPrimitives.scala 110:228:@13573.4]
  wire  _T_1007; // @[MemPrimitives.scala 110:228:@13577.4]
  wire  _T_1013; // @[MemPrimitives.scala 110:228:@13581.4]
  wire  _T_1019; // @[MemPrimitives.scala 110:228:@13585.4]
  wire  _T_1025; // @[MemPrimitives.scala 110:228:@13589.4]
  wire  _T_1027; // @[MemPrimitives.scala 123:41:@13600.4]
  wire  _T_1028; // @[MemPrimitives.scala 123:41:@13601.4]
  wire  _T_1029; // @[MemPrimitives.scala 123:41:@13602.4]
  wire  _T_1030; // @[MemPrimitives.scala 123:41:@13603.4]
  wire  _T_1031; // @[MemPrimitives.scala 123:41:@13604.4]
  wire  _T_1032; // @[MemPrimitives.scala 123:41:@13605.4]
  wire [10:0] _T_1034; // @[Cat.scala 30:58:@13607.4]
  wire [10:0] _T_1036; // @[Cat.scala 30:58:@13609.4]
  wire [10:0] _T_1038; // @[Cat.scala 30:58:@13611.4]
  wire [10:0] _T_1040; // @[Cat.scala 30:58:@13613.4]
  wire [10:0] _T_1042; // @[Cat.scala 30:58:@13615.4]
  wire [10:0] _T_1044; // @[Cat.scala 30:58:@13617.4]
  wire [10:0] _T_1045; // @[Mux.scala 31:69:@13618.4]
  wire [10:0] _T_1046; // @[Mux.scala 31:69:@13619.4]
  wire [10:0] _T_1047; // @[Mux.scala 31:69:@13620.4]
  wire [10:0] _T_1048; // @[Mux.scala 31:69:@13621.4]
  wire [10:0] _T_1049; // @[Mux.scala 31:69:@13622.4]
  wire  _T_1057; // @[MemPrimitives.scala 110:228:@13631.4]
  wire  _T_1063; // @[MemPrimitives.scala 110:228:@13635.4]
  wire  _T_1069; // @[MemPrimitives.scala 110:228:@13639.4]
  wire  _T_1075; // @[MemPrimitives.scala 110:228:@13643.4]
  wire  _T_1081; // @[MemPrimitives.scala 110:228:@13647.4]
  wire  _T_1087; // @[MemPrimitives.scala 110:228:@13651.4]
  wire  _T_1089; // @[MemPrimitives.scala 123:41:@13662.4]
  wire  _T_1090; // @[MemPrimitives.scala 123:41:@13663.4]
  wire  _T_1091; // @[MemPrimitives.scala 123:41:@13664.4]
  wire  _T_1092; // @[MemPrimitives.scala 123:41:@13665.4]
  wire  _T_1093; // @[MemPrimitives.scala 123:41:@13666.4]
  wire  _T_1094; // @[MemPrimitives.scala 123:41:@13667.4]
  wire [10:0] _T_1096; // @[Cat.scala 30:58:@13669.4]
  wire [10:0] _T_1098; // @[Cat.scala 30:58:@13671.4]
  wire [10:0] _T_1100; // @[Cat.scala 30:58:@13673.4]
  wire [10:0] _T_1102; // @[Cat.scala 30:58:@13675.4]
  wire [10:0] _T_1104; // @[Cat.scala 30:58:@13677.4]
  wire [10:0] _T_1106; // @[Cat.scala 30:58:@13679.4]
  wire [10:0] _T_1107; // @[Mux.scala 31:69:@13680.4]
  wire [10:0] _T_1108; // @[Mux.scala 31:69:@13681.4]
  wire [10:0] _T_1109; // @[Mux.scala 31:69:@13682.4]
  wire [10:0] _T_1110; // @[Mux.scala 31:69:@13683.4]
  wire [10:0] _T_1111; // @[Mux.scala 31:69:@13684.4]
  wire  _T_1116; // @[MemPrimitives.scala 110:210:@13691.4]
  wire  _T_1119; // @[MemPrimitives.scala 110:228:@13693.4]
  wire  _T_1122; // @[MemPrimitives.scala 110:210:@13695.4]
  wire  _T_1125; // @[MemPrimitives.scala 110:228:@13697.4]
  wire  _T_1128; // @[MemPrimitives.scala 110:210:@13699.4]
  wire  _T_1131; // @[MemPrimitives.scala 110:228:@13701.4]
  wire  _T_1134; // @[MemPrimitives.scala 110:210:@13703.4]
  wire  _T_1137; // @[MemPrimitives.scala 110:228:@13705.4]
  wire  _T_1140; // @[MemPrimitives.scala 110:210:@13707.4]
  wire  _T_1143; // @[MemPrimitives.scala 110:228:@13709.4]
  wire  _T_1146; // @[MemPrimitives.scala 110:210:@13711.4]
  wire  _T_1149; // @[MemPrimitives.scala 110:228:@13713.4]
  wire  _T_1151; // @[MemPrimitives.scala 123:41:@13724.4]
  wire  _T_1152; // @[MemPrimitives.scala 123:41:@13725.4]
  wire  _T_1153; // @[MemPrimitives.scala 123:41:@13726.4]
  wire  _T_1154; // @[MemPrimitives.scala 123:41:@13727.4]
  wire  _T_1155; // @[MemPrimitives.scala 123:41:@13728.4]
  wire  _T_1156; // @[MemPrimitives.scala 123:41:@13729.4]
  wire [10:0] _T_1158; // @[Cat.scala 30:58:@13731.4]
  wire [10:0] _T_1160; // @[Cat.scala 30:58:@13733.4]
  wire [10:0] _T_1162; // @[Cat.scala 30:58:@13735.4]
  wire [10:0] _T_1164; // @[Cat.scala 30:58:@13737.4]
  wire [10:0] _T_1166; // @[Cat.scala 30:58:@13739.4]
  wire [10:0] _T_1168; // @[Cat.scala 30:58:@13741.4]
  wire [10:0] _T_1169; // @[Mux.scala 31:69:@13742.4]
  wire [10:0] _T_1170; // @[Mux.scala 31:69:@13743.4]
  wire [10:0] _T_1171; // @[Mux.scala 31:69:@13744.4]
  wire [10:0] _T_1172; // @[Mux.scala 31:69:@13745.4]
  wire [10:0] _T_1173; // @[Mux.scala 31:69:@13746.4]
  wire  _T_1178; // @[MemPrimitives.scala 110:210:@13753.4]
  wire  _T_1181; // @[MemPrimitives.scala 110:228:@13755.4]
  wire  _T_1184; // @[MemPrimitives.scala 110:210:@13757.4]
  wire  _T_1187; // @[MemPrimitives.scala 110:228:@13759.4]
  wire  _T_1190; // @[MemPrimitives.scala 110:210:@13761.4]
  wire  _T_1193; // @[MemPrimitives.scala 110:228:@13763.4]
  wire  _T_1196; // @[MemPrimitives.scala 110:210:@13765.4]
  wire  _T_1199; // @[MemPrimitives.scala 110:228:@13767.4]
  wire  _T_1202; // @[MemPrimitives.scala 110:210:@13769.4]
  wire  _T_1205; // @[MemPrimitives.scala 110:228:@13771.4]
  wire  _T_1208; // @[MemPrimitives.scala 110:210:@13773.4]
  wire  _T_1211; // @[MemPrimitives.scala 110:228:@13775.4]
  wire  _T_1213; // @[MemPrimitives.scala 123:41:@13786.4]
  wire  _T_1214; // @[MemPrimitives.scala 123:41:@13787.4]
  wire  _T_1215; // @[MemPrimitives.scala 123:41:@13788.4]
  wire  _T_1216; // @[MemPrimitives.scala 123:41:@13789.4]
  wire  _T_1217; // @[MemPrimitives.scala 123:41:@13790.4]
  wire  _T_1218; // @[MemPrimitives.scala 123:41:@13791.4]
  wire [10:0] _T_1220; // @[Cat.scala 30:58:@13793.4]
  wire [10:0] _T_1222; // @[Cat.scala 30:58:@13795.4]
  wire [10:0] _T_1224; // @[Cat.scala 30:58:@13797.4]
  wire [10:0] _T_1226; // @[Cat.scala 30:58:@13799.4]
  wire [10:0] _T_1228; // @[Cat.scala 30:58:@13801.4]
  wire [10:0] _T_1230; // @[Cat.scala 30:58:@13803.4]
  wire [10:0] _T_1231; // @[Mux.scala 31:69:@13804.4]
  wire [10:0] _T_1232; // @[Mux.scala 31:69:@13805.4]
  wire [10:0] _T_1233; // @[Mux.scala 31:69:@13806.4]
  wire [10:0] _T_1234; // @[Mux.scala 31:69:@13807.4]
  wire [10:0] _T_1235; // @[Mux.scala 31:69:@13808.4]
  wire  _T_1243; // @[MemPrimitives.scala 110:228:@13817.4]
  wire  _T_1249; // @[MemPrimitives.scala 110:228:@13821.4]
  wire  _T_1255; // @[MemPrimitives.scala 110:228:@13825.4]
  wire  _T_1261; // @[MemPrimitives.scala 110:228:@13829.4]
  wire  _T_1267; // @[MemPrimitives.scala 110:228:@13833.4]
  wire  _T_1273; // @[MemPrimitives.scala 110:228:@13837.4]
  wire  _T_1275; // @[MemPrimitives.scala 123:41:@13848.4]
  wire  _T_1276; // @[MemPrimitives.scala 123:41:@13849.4]
  wire  _T_1277; // @[MemPrimitives.scala 123:41:@13850.4]
  wire  _T_1278; // @[MemPrimitives.scala 123:41:@13851.4]
  wire  _T_1279; // @[MemPrimitives.scala 123:41:@13852.4]
  wire  _T_1280; // @[MemPrimitives.scala 123:41:@13853.4]
  wire [10:0] _T_1282; // @[Cat.scala 30:58:@13855.4]
  wire [10:0] _T_1284; // @[Cat.scala 30:58:@13857.4]
  wire [10:0] _T_1286; // @[Cat.scala 30:58:@13859.4]
  wire [10:0] _T_1288; // @[Cat.scala 30:58:@13861.4]
  wire [10:0] _T_1290; // @[Cat.scala 30:58:@13863.4]
  wire [10:0] _T_1292; // @[Cat.scala 30:58:@13865.4]
  wire [10:0] _T_1293; // @[Mux.scala 31:69:@13866.4]
  wire [10:0] _T_1294; // @[Mux.scala 31:69:@13867.4]
  wire [10:0] _T_1295; // @[Mux.scala 31:69:@13868.4]
  wire [10:0] _T_1296; // @[Mux.scala 31:69:@13869.4]
  wire [10:0] _T_1297; // @[Mux.scala 31:69:@13870.4]
  wire  _T_1305; // @[MemPrimitives.scala 110:228:@13879.4]
  wire  _T_1311; // @[MemPrimitives.scala 110:228:@13883.4]
  wire  _T_1317; // @[MemPrimitives.scala 110:228:@13887.4]
  wire  _T_1323; // @[MemPrimitives.scala 110:228:@13891.4]
  wire  _T_1329; // @[MemPrimitives.scala 110:228:@13895.4]
  wire  _T_1335; // @[MemPrimitives.scala 110:228:@13899.4]
  wire  _T_1337; // @[MemPrimitives.scala 123:41:@13910.4]
  wire  _T_1338; // @[MemPrimitives.scala 123:41:@13911.4]
  wire  _T_1339; // @[MemPrimitives.scala 123:41:@13912.4]
  wire  _T_1340; // @[MemPrimitives.scala 123:41:@13913.4]
  wire  _T_1341; // @[MemPrimitives.scala 123:41:@13914.4]
  wire  _T_1342; // @[MemPrimitives.scala 123:41:@13915.4]
  wire [10:0] _T_1344; // @[Cat.scala 30:58:@13917.4]
  wire [10:0] _T_1346; // @[Cat.scala 30:58:@13919.4]
  wire [10:0] _T_1348; // @[Cat.scala 30:58:@13921.4]
  wire [10:0] _T_1350; // @[Cat.scala 30:58:@13923.4]
  wire [10:0] _T_1352; // @[Cat.scala 30:58:@13925.4]
  wire [10:0] _T_1354; // @[Cat.scala 30:58:@13927.4]
  wire [10:0] _T_1355; // @[Mux.scala 31:69:@13928.4]
  wire [10:0] _T_1356; // @[Mux.scala 31:69:@13929.4]
  wire [10:0] _T_1357; // @[Mux.scala 31:69:@13930.4]
  wire [10:0] _T_1358; // @[Mux.scala 31:69:@13931.4]
  wire [10:0] _T_1359; // @[Mux.scala 31:69:@13932.4]
  wire  _T_1364; // @[MemPrimitives.scala 110:210:@13939.4]
  wire  _T_1367; // @[MemPrimitives.scala 110:228:@13941.4]
  wire  _T_1370; // @[MemPrimitives.scala 110:210:@13943.4]
  wire  _T_1373; // @[MemPrimitives.scala 110:228:@13945.4]
  wire  _T_1376; // @[MemPrimitives.scala 110:210:@13947.4]
  wire  _T_1379; // @[MemPrimitives.scala 110:228:@13949.4]
  wire  _T_1382; // @[MemPrimitives.scala 110:210:@13951.4]
  wire  _T_1385; // @[MemPrimitives.scala 110:228:@13953.4]
  wire  _T_1388; // @[MemPrimitives.scala 110:210:@13955.4]
  wire  _T_1391; // @[MemPrimitives.scala 110:228:@13957.4]
  wire  _T_1394; // @[MemPrimitives.scala 110:210:@13959.4]
  wire  _T_1397; // @[MemPrimitives.scala 110:228:@13961.4]
  wire  _T_1399; // @[MemPrimitives.scala 123:41:@13972.4]
  wire  _T_1400; // @[MemPrimitives.scala 123:41:@13973.4]
  wire  _T_1401; // @[MemPrimitives.scala 123:41:@13974.4]
  wire  _T_1402; // @[MemPrimitives.scala 123:41:@13975.4]
  wire  _T_1403; // @[MemPrimitives.scala 123:41:@13976.4]
  wire  _T_1404; // @[MemPrimitives.scala 123:41:@13977.4]
  wire [10:0] _T_1406; // @[Cat.scala 30:58:@13979.4]
  wire [10:0] _T_1408; // @[Cat.scala 30:58:@13981.4]
  wire [10:0] _T_1410; // @[Cat.scala 30:58:@13983.4]
  wire [10:0] _T_1412; // @[Cat.scala 30:58:@13985.4]
  wire [10:0] _T_1414; // @[Cat.scala 30:58:@13987.4]
  wire [10:0] _T_1416; // @[Cat.scala 30:58:@13989.4]
  wire [10:0] _T_1417; // @[Mux.scala 31:69:@13990.4]
  wire [10:0] _T_1418; // @[Mux.scala 31:69:@13991.4]
  wire [10:0] _T_1419; // @[Mux.scala 31:69:@13992.4]
  wire [10:0] _T_1420; // @[Mux.scala 31:69:@13993.4]
  wire [10:0] _T_1421; // @[Mux.scala 31:69:@13994.4]
  wire  _T_1426; // @[MemPrimitives.scala 110:210:@14001.4]
  wire  _T_1429; // @[MemPrimitives.scala 110:228:@14003.4]
  wire  _T_1432; // @[MemPrimitives.scala 110:210:@14005.4]
  wire  _T_1435; // @[MemPrimitives.scala 110:228:@14007.4]
  wire  _T_1438; // @[MemPrimitives.scala 110:210:@14009.4]
  wire  _T_1441; // @[MemPrimitives.scala 110:228:@14011.4]
  wire  _T_1444; // @[MemPrimitives.scala 110:210:@14013.4]
  wire  _T_1447; // @[MemPrimitives.scala 110:228:@14015.4]
  wire  _T_1450; // @[MemPrimitives.scala 110:210:@14017.4]
  wire  _T_1453; // @[MemPrimitives.scala 110:228:@14019.4]
  wire  _T_1456; // @[MemPrimitives.scala 110:210:@14021.4]
  wire  _T_1459; // @[MemPrimitives.scala 110:228:@14023.4]
  wire  _T_1461; // @[MemPrimitives.scala 123:41:@14034.4]
  wire  _T_1462; // @[MemPrimitives.scala 123:41:@14035.4]
  wire  _T_1463; // @[MemPrimitives.scala 123:41:@14036.4]
  wire  _T_1464; // @[MemPrimitives.scala 123:41:@14037.4]
  wire  _T_1465; // @[MemPrimitives.scala 123:41:@14038.4]
  wire  _T_1466; // @[MemPrimitives.scala 123:41:@14039.4]
  wire [10:0] _T_1468; // @[Cat.scala 30:58:@14041.4]
  wire [10:0] _T_1470; // @[Cat.scala 30:58:@14043.4]
  wire [10:0] _T_1472; // @[Cat.scala 30:58:@14045.4]
  wire [10:0] _T_1474; // @[Cat.scala 30:58:@14047.4]
  wire [10:0] _T_1476; // @[Cat.scala 30:58:@14049.4]
  wire [10:0] _T_1478; // @[Cat.scala 30:58:@14051.4]
  wire [10:0] _T_1479; // @[Mux.scala 31:69:@14052.4]
  wire [10:0] _T_1480; // @[Mux.scala 31:69:@14053.4]
  wire [10:0] _T_1481; // @[Mux.scala 31:69:@14054.4]
  wire [10:0] _T_1482; // @[Mux.scala 31:69:@14055.4]
  wire [10:0] _T_1483; // @[Mux.scala 31:69:@14056.4]
  wire  _T_1491; // @[MemPrimitives.scala 110:228:@14065.4]
  wire  _T_1497; // @[MemPrimitives.scala 110:228:@14069.4]
  wire  _T_1503; // @[MemPrimitives.scala 110:228:@14073.4]
  wire  _T_1509; // @[MemPrimitives.scala 110:228:@14077.4]
  wire  _T_1515; // @[MemPrimitives.scala 110:228:@14081.4]
  wire  _T_1521; // @[MemPrimitives.scala 110:228:@14085.4]
  wire  _T_1523; // @[MemPrimitives.scala 123:41:@14096.4]
  wire  _T_1524; // @[MemPrimitives.scala 123:41:@14097.4]
  wire  _T_1525; // @[MemPrimitives.scala 123:41:@14098.4]
  wire  _T_1526; // @[MemPrimitives.scala 123:41:@14099.4]
  wire  _T_1527; // @[MemPrimitives.scala 123:41:@14100.4]
  wire  _T_1528; // @[MemPrimitives.scala 123:41:@14101.4]
  wire [10:0] _T_1530; // @[Cat.scala 30:58:@14103.4]
  wire [10:0] _T_1532; // @[Cat.scala 30:58:@14105.4]
  wire [10:0] _T_1534; // @[Cat.scala 30:58:@14107.4]
  wire [10:0] _T_1536; // @[Cat.scala 30:58:@14109.4]
  wire [10:0] _T_1538; // @[Cat.scala 30:58:@14111.4]
  wire [10:0] _T_1540; // @[Cat.scala 30:58:@14113.4]
  wire [10:0] _T_1541; // @[Mux.scala 31:69:@14114.4]
  wire [10:0] _T_1542; // @[Mux.scala 31:69:@14115.4]
  wire [10:0] _T_1543; // @[Mux.scala 31:69:@14116.4]
  wire [10:0] _T_1544; // @[Mux.scala 31:69:@14117.4]
  wire [10:0] _T_1545; // @[Mux.scala 31:69:@14118.4]
  wire  _T_1553; // @[MemPrimitives.scala 110:228:@14127.4]
  wire  _T_1559; // @[MemPrimitives.scala 110:228:@14131.4]
  wire  _T_1565; // @[MemPrimitives.scala 110:228:@14135.4]
  wire  _T_1571; // @[MemPrimitives.scala 110:228:@14139.4]
  wire  _T_1577; // @[MemPrimitives.scala 110:228:@14143.4]
  wire  _T_1583; // @[MemPrimitives.scala 110:228:@14147.4]
  wire  _T_1585; // @[MemPrimitives.scala 123:41:@14158.4]
  wire  _T_1586; // @[MemPrimitives.scala 123:41:@14159.4]
  wire  _T_1587; // @[MemPrimitives.scala 123:41:@14160.4]
  wire  _T_1588; // @[MemPrimitives.scala 123:41:@14161.4]
  wire  _T_1589; // @[MemPrimitives.scala 123:41:@14162.4]
  wire  _T_1590; // @[MemPrimitives.scala 123:41:@14163.4]
  wire [10:0] _T_1592; // @[Cat.scala 30:58:@14165.4]
  wire [10:0] _T_1594; // @[Cat.scala 30:58:@14167.4]
  wire [10:0] _T_1596; // @[Cat.scala 30:58:@14169.4]
  wire [10:0] _T_1598; // @[Cat.scala 30:58:@14171.4]
  wire [10:0] _T_1600; // @[Cat.scala 30:58:@14173.4]
  wire [10:0] _T_1602; // @[Cat.scala 30:58:@14175.4]
  wire [10:0] _T_1603; // @[Mux.scala 31:69:@14176.4]
  wire [10:0] _T_1604; // @[Mux.scala 31:69:@14177.4]
  wire [10:0] _T_1605; // @[Mux.scala 31:69:@14178.4]
  wire [10:0] _T_1606; // @[Mux.scala 31:69:@14179.4]
  wire [10:0] _T_1607; // @[Mux.scala 31:69:@14180.4]
  wire  _T_1671; // @[package.scala 96:25:@14265.4 package.scala 96:25:@14266.4]
  wire [7:0] _T_1675; // @[Mux.scala 31:69:@14275.4]
  wire  _T_1668; // @[package.scala 96:25:@14257.4 package.scala 96:25:@14258.4]
  wire [7:0] _T_1676; // @[Mux.scala 31:69:@14276.4]
  wire  _T_1665; // @[package.scala 96:25:@14249.4 package.scala 96:25:@14250.4]
  wire [7:0] _T_1677; // @[Mux.scala 31:69:@14277.4]
  wire  _T_1662; // @[package.scala 96:25:@14241.4 package.scala 96:25:@14242.4]
  wire [7:0] _T_1678; // @[Mux.scala 31:69:@14278.4]
  wire  _T_1659; // @[package.scala 96:25:@14233.4 package.scala 96:25:@14234.4]
  wire [7:0] _T_1679; // @[Mux.scala 31:69:@14279.4]
  wire  _T_1656; // @[package.scala 96:25:@14225.4 package.scala 96:25:@14226.4]
  wire [7:0] _T_1680; // @[Mux.scala 31:69:@14280.4]
  wire  _T_1653; // @[package.scala 96:25:@14217.4 package.scala 96:25:@14218.4]
  wire  _T_1742; // @[package.scala 96:25:@14361.4 package.scala 96:25:@14362.4]
  wire [7:0] _T_1746; // @[Mux.scala 31:69:@14371.4]
  wire  _T_1739; // @[package.scala 96:25:@14353.4 package.scala 96:25:@14354.4]
  wire [7:0] _T_1747; // @[Mux.scala 31:69:@14372.4]
  wire  _T_1736; // @[package.scala 96:25:@14345.4 package.scala 96:25:@14346.4]
  wire [7:0] _T_1748; // @[Mux.scala 31:69:@14373.4]
  wire  _T_1733; // @[package.scala 96:25:@14337.4 package.scala 96:25:@14338.4]
  wire [7:0] _T_1749; // @[Mux.scala 31:69:@14374.4]
  wire  _T_1730; // @[package.scala 96:25:@14329.4 package.scala 96:25:@14330.4]
  wire [7:0] _T_1750; // @[Mux.scala 31:69:@14375.4]
  wire  _T_1727; // @[package.scala 96:25:@14321.4 package.scala 96:25:@14322.4]
  wire [7:0] _T_1751; // @[Mux.scala 31:69:@14376.4]
  wire  _T_1724; // @[package.scala 96:25:@14313.4 package.scala 96:25:@14314.4]
  wire  _T_1813; // @[package.scala 96:25:@14457.4 package.scala 96:25:@14458.4]
  wire [7:0] _T_1817; // @[Mux.scala 31:69:@14467.4]
  wire  _T_1810; // @[package.scala 96:25:@14449.4 package.scala 96:25:@14450.4]
  wire [7:0] _T_1818; // @[Mux.scala 31:69:@14468.4]
  wire  _T_1807; // @[package.scala 96:25:@14441.4 package.scala 96:25:@14442.4]
  wire [7:0] _T_1819; // @[Mux.scala 31:69:@14469.4]
  wire  _T_1804; // @[package.scala 96:25:@14433.4 package.scala 96:25:@14434.4]
  wire [7:0] _T_1820; // @[Mux.scala 31:69:@14470.4]
  wire  _T_1801; // @[package.scala 96:25:@14425.4 package.scala 96:25:@14426.4]
  wire [7:0] _T_1821; // @[Mux.scala 31:69:@14471.4]
  wire  _T_1798; // @[package.scala 96:25:@14417.4 package.scala 96:25:@14418.4]
  wire [7:0] _T_1822; // @[Mux.scala 31:69:@14472.4]
  wire  _T_1795; // @[package.scala 96:25:@14409.4 package.scala 96:25:@14410.4]
  wire  _T_1884; // @[package.scala 96:25:@14553.4 package.scala 96:25:@14554.4]
  wire [7:0] _T_1888; // @[Mux.scala 31:69:@14563.4]
  wire  _T_1881; // @[package.scala 96:25:@14545.4 package.scala 96:25:@14546.4]
  wire [7:0] _T_1889; // @[Mux.scala 31:69:@14564.4]
  wire  _T_1878; // @[package.scala 96:25:@14537.4 package.scala 96:25:@14538.4]
  wire [7:0] _T_1890; // @[Mux.scala 31:69:@14565.4]
  wire  _T_1875; // @[package.scala 96:25:@14529.4 package.scala 96:25:@14530.4]
  wire [7:0] _T_1891; // @[Mux.scala 31:69:@14566.4]
  wire  _T_1872; // @[package.scala 96:25:@14521.4 package.scala 96:25:@14522.4]
  wire [7:0] _T_1892; // @[Mux.scala 31:69:@14567.4]
  wire  _T_1869; // @[package.scala 96:25:@14513.4 package.scala 96:25:@14514.4]
  wire [7:0] _T_1893; // @[Mux.scala 31:69:@14568.4]
  wire  _T_1866; // @[package.scala 96:25:@14505.4 package.scala 96:25:@14506.4]
  wire  _T_1955; // @[package.scala 96:25:@14649.4 package.scala 96:25:@14650.4]
  wire [7:0] _T_1959; // @[Mux.scala 31:69:@14659.4]
  wire  _T_1952; // @[package.scala 96:25:@14641.4 package.scala 96:25:@14642.4]
  wire [7:0] _T_1960; // @[Mux.scala 31:69:@14660.4]
  wire  _T_1949; // @[package.scala 96:25:@14633.4 package.scala 96:25:@14634.4]
  wire [7:0] _T_1961; // @[Mux.scala 31:69:@14661.4]
  wire  _T_1946; // @[package.scala 96:25:@14625.4 package.scala 96:25:@14626.4]
  wire [7:0] _T_1962; // @[Mux.scala 31:69:@14662.4]
  wire  _T_1943; // @[package.scala 96:25:@14617.4 package.scala 96:25:@14618.4]
  wire [7:0] _T_1963; // @[Mux.scala 31:69:@14663.4]
  wire  _T_1940; // @[package.scala 96:25:@14609.4 package.scala 96:25:@14610.4]
  wire [7:0] _T_1964; // @[Mux.scala 31:69:@14664.4]
  wire  _T_1937; // @[package.scala 96:25:@14601.4 package.scala 96:25:@14602.4]
  wire  _T_2026; // @[package.scala 96:25:@14745.4 package.scala 96:25:@14746.4]
  wire [7:0] _T_2030; // @[Mux.scala 31:69:@14755.4]
  wire  _T_2023; // @[package.scala 96:25:@14737.4 package.scala 96:25:@14738.4]
  wire [7:0] _T_2031; // @[Mux.scala 31:69:@14756.4]
  wire  _T_2020; // @[package.scala 96:25:@14729.4 package.scala 96:25:@14730.4]
  wire [7:0] _T_2032; // @[Mux.scala 31:69:@14757.4]
  wire  _T_2017; // @[package.scala 96:25:@14721.4 package.scala 96:25:@14722.4]
  wire [7:0] _T_2033; // @[Mux.scala 31:69:@14758.4]
  wire  _T_2014; // @[package.scala 96:25:@14713.4 package.scala 96:25:@14714.4]
  wire [7:0] _T_2034; // @[Mux.scala 31:69:@14759.4]
  wire  _T_2011; // @[package.scala 96:25:@14705.4 package.scala 96:25:@14706.4]
  wire [7:0] _T_2035; // @[Mux.scala 31:69:@14760.4]
  wire  _T_2008; // @[package.scala 96:25:@14697.4 package.scala 96:25:@14698.4]
  wire  _T_2097; // @[package.scala 96:25:@14841.4 package.scala 96:25:@14842.4]
  wire [7:0] _T_2101; // @[Mux.scala 31:69:@14851.4]
  wire  _T_2094; // @[package.scala 96:25:@14833.4 package.scala 96:25:@14834.4]
  wire [7:0] _T_2102; // @[Mux.scala 31:69:@14852.4]
  wire  _T_2091; // @[package.scala 96:25:@14825.4 package.scala 96:25:@14826.4]
  wire [7:0] _T_2103; // @[Mux.scala 31:69:@14853.4]
  wire  _T_2088; // @[package.scala 96:25:@14817.4 package.scala 96:25:@14818.4]
  wire [7:0] _T_2104; // @[Mux.scala 31:69:@14854.4]
  wire  _T_2085; // @[package.scala 96:25:@14809.4 package.scala 96:25:@14810.4]
  wire [7:0] _T_2105; // @[Mux.scala 31:69:@14855.4]
  wire  _T_2082; // @[package.scala 96:25:@14801.4 package.scala 96:25:@14802.4]
  wire [7:0] _T_2106; // @[Mux.scala 31:69:@14856.4]
  wire  _T_2079; // @[package.scala 96:25:@14793.4 package.scala 96:25:@14794.4]
  wire  _T_2168; // @[package.scala 96:25:@14937.4 package.scala 96:25:@14938.4]
  wire [7:0] _T_2172; // @[Mux.scala 31:69:@14947.4]
  wire  _T_2165; // @[package.scala 96:25:@14929.4 package.scala 96:25:@14930.4]
  wire [7:0] _T_2173; // @[Mux.scala 31:69:@14948.4]
  wire  _T_2162; // @[package.scala 96:25:@14921.4 package.scala 96:25:@14922.4]
  wire [7:0] _T_2174; // @[Mux.scala 31:69:@14949.4]
  wire  _T_2159; // @[package.scala 96:25:@14913.4 package.scala 96:25:@14914.4]
  wire [7:0] _T_2175; // @[Mux.scala 31:69:@14950.4]
  wire  _T_2156; // @[package.scala 96:25:@14905.4 package.scala 96:25:@14906.4]
  wire [7:0] _T_2176; // @[Mux.scala 31:69:@14951.4]
  wire  _T_2153; // @[package.scala 96:25:@14897.4 package.scala 96:25:@14898.4]
  wire [7:0] _T_2177; // @[Mux.scala 31:69:@14952.4]
  wire  _T_2150; // @[package.scala 96:25:@14889.4 package.scala 96:25:@14890.4]
  wire  _T_2239; // @[package.scala 96:25:@15033.4 package.scala 96:25:@15034.4]
  wire [7:0] _T_2243; // @[Mux.scala 31:69:@15043.4]
  wire  _T_2236; // @[package.scala 96:25:@15025.4 package.scala 96:25:@15026.4]
  wire [7:0] _T_2244; // @[Mux.scala 31:69:@15044.4]
  wire  _T_2233; // @[package.scala 96:25:@15017.4 package.scala 96:25:@15018.4]
  wire [7:0] _T_2245; // @[Mux.scala 31:69:@15045.4]
  wire  _T_2230; // @[package.scala 96:25:@15009.4 package.scala 96:25:@15010.4]
  wire [7:0] _T_2246; // @[Mux.scala 31:69:@15046.4]
  wire  _T_2227; // @[package.scala 96:25:@15001.4 package.scala 96:25:@15002.4]
  wire [7:0] _T_2247; // @[Mux.scala 31:69:@15047.4]
  wire  _T_2224; // @[package.scala 96:25:@14993.4 package.scala 96:25:@14994.4]
  wire [7:0] _T_2248; // @[Mux.scala 31:69:@15048.4]
  wire  _T_2221; // @[package.scala 96:25:@14985.4 package.scala 96:25:@14986.4]
  wire  _T_2310; // @[package.scala 96:25:@15129.4 package.scala 96:25:@15130.4]
  wire [7:0] _T_2314; // @[Mux.scala 31:69:@15139.4]
  wire  _T_2307; // @[package.scala 96:25:@15121.4 package.scala 96:25:@15122.4]
  wire [7:0] _T_2315; // @[Mux.scala 31:69:@15140.4]
  wire  _T_2304; // @[package.scala 96:25:@15113.4 package.scala 96:25:@15114.4]
  wire [7:0] _T_2316; // @[Mux.scala 31:69:@15141.4]
  wire  _T_2301; // @[package.scala 96:25:@15105.4 package.scala 96:25:@15106.4]
  wire [7:0] _T_2317; // @[Mux.scala 31:69:@15142.4]
  wire  _T_2298; // @[package.scala 96:25:@15097.4 package.scala 96:25:@15098.4]
  wire [7:0] _T_2318; // @[Mux.scala 31:69:@15143.4]
  wire  _T_2295; // @[package.scala 96:25:@15089.4 package.scala 96:25:@15090.4]
  wire [7:0] _T_2319; // @[Mux.scala 31:69:@15144.4]
  wire  _T_2292; // @[package.scala 96:25:@15081.4 package.scala 96:25:@15082.4]
  wire  _T_2381; // @[package.scala 96:25:@15225.4 package.scala 96:25:@15226.4]
  wire [7:0] _T_2385; // @[Mux.scala 31:69:@15235.4]
  wire  _T_2378; // @[package.scala 96:25:@15217.4 package.scala 96:25:@15218.4]
  wire [7:0] _T_2386; // @[Mux.scala 31:69:@15236.4]
  wire  _T_2375; // @[package.scala 96:25:@15209.4 package.scala 96:25:@15210.4]
  wire [7:0] _T_2387; // @[Mux.scala 31:69:@15237.4]
  wire  _T_2372; // @[package.scala 96:25:@15201.4 package.scala 96:25:@15202.4]
  wire [7:0] _T_2388; // @[Mux.scala 31:69:@15238.4]
  wire  _T_2369; // @[package.scala 96:25:@15193.4 package.scala 96:25:@15194.4]
  wire [7:0] _T_2389; // @[Mux.scala 31:69:@15239.4]
  wire  _T_2366; // @[package.scala 96:25:@15185.4 package.scala 96:25:@15186.4]
  wire [7:0] _T_2390; // @[Mux.scala 31:69:@15240.4]
  wire  _T_2363; // @[package.scala 96:25:@15177.4 package.scala 96:25:@15178.4]
  wire  _T_2452; // @[package.scala 96:25:@15321.4 package.scala 96:25:@15322.4]
  wire [7:0] _T_2456; // @[Mux.scala 31:69:@15331.4]
  wire  _T_2449; // @[package.scala 96:25:@15313.4 package.scala 96:25:@15314.4]
  wire [7:0] _T_2457; // @[Mux.scala 31:69:@15332.4]
  wire  _T_2446; // @[package.scala 96:25:@15305.4 package.scala 96:25:@15306.4]
  wire [7:0] _T_2458; // @[Mux.scala 31:69:@15333.4]
  wire  _T_2443; // @[package.scala 96:25:@15297.4 package.scala 96:25:@15298.4]
  wire [7:0] _T_2459; // @[Mux.scala 31:69:@15334.4]
  wire  _T_2440; // @[package.scala 96:25:@15289.4 package.scala 96:25:@15290.4]
  wire [7:0] _T_2460; // @[Mux.scala 31:69:@15335.4]
  wire  _T_2437; // @[package.scala 96:25:@15281.4 package.scala 96:25:@15282.4]
  wire [7:0] _T_2461; // @[Mux.scala 31:69:@15336.4]
  wire  _T_2434; // @[package.scala 96:25:@15273.4 package.scala 96:25:@15274.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@12747.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@12763.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@12779.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@12795.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@12811.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@12827.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@12843.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@12859.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@12875.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@12891.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@12907.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@12923.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_5 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@12939.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_5 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@12955.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_5 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@12971.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_5 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@12987.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects_1 StickySelects ( // @[MemPrimitives.scala 121:29:@13219.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5)
  );
  StickySelects_1 StickySelects_1 ( // @[MemPrimitives.scala 121:29:@13281.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5)
  );
  StickySelects_1 StickySelects_2 ( // @[MemPrimitives.scala 121:29:@13343.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5)
  );
  StickySelects_1 StickySelects_3 ( // @[MemPrimitives.scala 121:29:@13405.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5)
  );
  StickySelects_1 StickySelects_4 ( // @[MemPrimitives.scala 121:29:@13467.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5)
  );
  StickySelects_1 StickySelects_5 ( // @[MemPrimitives.scala 121:29:@13529.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5)
  );
  StickySelects_1 StickySelects_6 ( // @[MemPrimitives.scala 121:29:@13591.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5)
  );
  StickySelects_1 StickySelects_7 ( // @[MemPrimitives.scala 121:29:@13653.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5)
  );
  StickySelects_1 StickySelects_8 ( // @[MemPrimitives.scala 121:29:@13715.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5)
  );
  StickySelects_1 StickySelects_9 ( // @[MemPrimitives.scala 121:29:@13777.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5)
  );
  StickySelects_1 StickySelects_10 ( // @[MemPrimitives.scala 121:29:@13839.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5)
  );
  StickySelects_1 StickySelects_11 ( // @[MemPrimitives.scala 121:29:@13901.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5)
  );
  StickySelects_1 StickySelects_12 ( // @[MemPrimitives.scala 121:29:@13963.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_ins_4(StickySelects_12_io_ins_4),
    .io_ins_5(StickySelects_12_io_ins_5),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3),
    .io_outs_4(StickySelects_12_io_outs_4),
    .io_outs_5(StickySelects_12_io_outs_5)
  );
  StickySelects_1 StickySelects_13 ( // @[MemPrimitives.scala 121:29:@14025.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_ins_4(StickySelects_13_io_ins_4),
    .io_ins_5(StickySelects_13_io_ins_5),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3),
    .io_outs_4(StickySelects_13_io_outs_4),
    .io_outs_5(StickySelects_13_io_outs_5)
  );
  StickySelects_1 StickySelects_14 ( // @[MemPrimitives.scala 121:29:@14087.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5)
  );
  StickySelects_1 StickySelects_15 ( // @[MemPrimitives.scala 121:29:@14149.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@14212.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@14220.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@14228.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@14236.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@14244.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@14252.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@14260.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@14268.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@14308.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@14316.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@14324.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@14332.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@14340.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@14348.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@14356.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@14364.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@14404.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@14412.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@14420.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@14428.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@14436.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@14444.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@14452.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@14460.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@14500.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@14508.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@14516.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@14524.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@14532.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@14540.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@14548.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@14556.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@14596.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@14604.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@14612.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@14620.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@14628.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@14636.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@14644.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@14652.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@14692.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@14700.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@14708.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@14716.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@14724.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@14732.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@14740.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@14748.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_48 ( // @[package.scala 93:22:@14788.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@14796.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_50 ( // @[package.scala 93:22:@14804.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@14812.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@14820.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_53 ( // @[package.scala 93:22:@14828.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@14836.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_55 ( // @[package.scala 93:22:@14844.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@14884.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_57 ( // @[package.scala 93:22:@14892.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@14900.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_59 ( // @[package.scala 93:22:@14908.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_60 ( // @[package.scala 93:22:@14916.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_61 ( // @[package.scala 93:22:@14924.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_62 ( // @[package.scala 93:22:@14932.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_63 ( // @[package.scala 93:22:@14940.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_64 ( // @[package.scala 93:22:@14980.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_65 ( // @[package.scala 93:22:@14988.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_66 ( // @[package.scala 93:22:@14996.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_67 ( // @[package.scala 93:22:@15004.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_68 ( // @[package.scala 93:22:@15012.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_69 ( // @[package.scala 93:22:@15020.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_70 ( // @[package.scala 93:22:@15028.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_71 ( // @[package.scala 93:22:@15036.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_72 ( // @[package.scala 93:22:@15076.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_73 ( // @[package.scala 93:22:@15084.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_74 ( // @[package.scala 93:22:@15092.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_75 ( // @[package.scala 93:22:@15100.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_76 ( // @[package.scala 93:22:@15108.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_77 ( // @[package.scala 93:22:@15116.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_78 ( // @[package.scala 93:22:@15124.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_79 ( // @[package.scala 93:22:@15132.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_80 ( // @[package.scala 93:22:@15172.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_81 ( // @[package.scala 93:22:@15180.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_82 ( // @[package.scala 93:22:@15188.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_83 ( // @[package.scala 93:22:@15196.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_84 ( // @[package.scala 93:22:@15204.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_85 ( // @[package.scala 93:22:@15212.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_86 ( // @[package.scala 93:22:@15220.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_87 ( // @[package.scala 93:22:@15228.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_88 ( // @[package.scala 93:22:@15268.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_89 ( // @[package.scala 93:22:@15276.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_90 ( // @[package.scala 93:22:@15284.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_91 ( // @[package.scala 93:22:@15292.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_92 ( // @[package.scala 93:22:@15300.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_93 ( // @[package.scala 93:22:@15308.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_94 ( // @[package.scala 93:22:@15316.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_95 ( // @[package.scala 93:22:@15324.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  assign _T_444 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@13003.4]
  assign _T_446 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@13004.4]
  assign _T_447 = _T_444 & _T_446; // @[MemPrimitives.scala 82:228:@13005.4]
  assign _T_448 = io_wPort_0_en_0 & _T_447; // @[MemPrimitives.scala 83:102:@13006.4]
  assign _T_450 = {_T_448,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13008.4]
  assign _T_455 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@13015.4]
  assign _T_457 = io_wPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@13016.4]
  assign _T_458 = _T_455 & _T_457; // @[MemPrimitives.scala 82:228:@13017.4]
  assign _T_459 = io_wPort_1_en_0 & _T_458; // @[MemPrimitives.scala 83:102:@13018.4]
  assign _T_461 = {_T_459,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13020.4]
  assign _T_468 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@13028.4]
  assign _T_469 = _T_444 & _T_468; // @[MemPrimitives.scala 82:228:@13029.4]
  assign _T_470 = io_wPort_0_en_0 & _T_469; // @[MemPrimitives.scala 83:102:@13030.4]
  assign _T_472 = {_T_470,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13032.4]
  assign _T_479 = io_wPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@13040.4]
  assign _T_480 = _T_455 & _T_479; // @[MemPrimitives.scala 82:228:@13041.4]
  assign _T_481 = io_wPort_1_en_0 & _T_480; // @[MemPrimitives.scala 83:102:@13042.4]
  assign _T_483 = {_T_481,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13044.4]
  assign _T_488 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@13051.4]
  assign _T_491 = _T_488 & _T_446; // @[MemPrimitives.scala 82:228:@13053.4]
  assign _T_492 = io_wPort_0_en_0 & _T_491; // @[MemPrimitives.scala 83:102:@13054.4]
  assign _T_494 = {_T_492,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13056.4]
  assign _T_499 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@13063.4]
  assign _T_502 = _T_499 & _T_457; // @[MemPrimitives.scala 82:228:@13065.4]
  assign _T_503 = io_wPort_1_en_0 & _T_502; // @[MemPrimitives.scala 83:102:@13066.4]
  assign _T_505 = {_T_503,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13068.4]
  assign _T_513 = _T_488 & _T_468; // @[MemPrimitives.scala 82:228:@13077.4]
  assign _T_514 = io_wPort_0_en_0 & _T_513; // @[MemPrimitives.scala 83:102:@13078.4]
  assign _T_516 = {_T_514,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13080.4]
  assign _T_524 = _T_499 & _T_479; // @[MemPrimitives.scala 82:228:@13089.4]
  assign _T_525 = io_wPort_1_en_0 & _T_524; // @[MemPrimitives.scala 83:102:@13090.4]
  assign _T_527 = {_T_525,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13092.4]
  assign _T_532 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@13099.4]
  assign _T_535 = _T_532 & _T_446; // @[MemPrimitives.scala 82:228:@13101.4]
  assign _T_536 = io_wPort_0_en_0 & _T_535; // @[MemPrimitives.scala 83:102:@13102.4]
  assign _T_538 = {_T_536,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13104.4]
  assign _T_543 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@13111.4]
  assign _T_546 = _T_543 & _T_457; // @[MemPrimitives.scala 82:228:@13113.4]
  assign _T_547 = io_wPort_1_en_0 & _T_546; // @[MemPrimitives.scala 83:102:@13114.4]
  assign _T_549 = {_T_547,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13116.4]
  assign _T_557 = _T_532 & _T_468; // @[MemPrimitives.scala 82:228:@13125.4]
  assign _T_558 = io_wPort_0_en_0 & _T_557; // @[MemPrimitives.scala 83:102:@13126.4]
  assign _T_560 = {_T_558,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13128.4]
  assign _T_568 = _T_543 & _T_479; // @[MemPrimitives.scala 82:228:@13137.4]
  assign _T_569 = io_wPort_1_en_0 & _T_568; // @[MemPrimitives.scala 83:102:@13138.4]
  assign _T_571 = {_T_569,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13140.4]
  assign _T_576 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@13147.4]
  assign _T_579 = _T_576 & _T_446; // @[MemPrimitives.scala 82:228:@13149.4]
  assign _T_580 = io_wPort_0_en_0 & _T_579; // @[MemPrimitives.scala 83:102:@13150.4]
  assign _T_582 = {_T_580,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13152.4]
  assign _T_587 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@13159.4]
  assign _T_590 = _T_587 & _T_457; // @[MemPrimitives.scala 82:228:@13161.4]
  assign _T_591 = io_wPort_1_en_0 & _T_590; // @[MemPrimitives.scala 83:102:@13162.4]
  assign _T_593 = {_T_591,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13164.4]
  assign _T_601 = _T_576 & _T_468; // @[MemPrimitives.scala 82:228:@13173.4]
  assign _T_602 = io_wPort_0_en_0 & _T_601; // @[MemPrimitives.scala 83:102:@13174.4]
  assign _T_604 = {_T_602,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13176.4]
  assign _T_612 = _T_587 & _T_479; // @[MemPrimitives.scala 82:228:@13185.4]
  assign _T_613 = io_wPort_1_en_0 & _T_612; // @[MemPrimitives.scala 83:102:@13186.4]
  assign _T_615 = {_T_613,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13188.4]
  assign _T_620 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13195.4]
  assign _T_622 = io_rPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13196.4]
  assign _T_623 = _T_620 & _T_622; // @[MemPrimitives.scala 110:228:@13197.4]
  assign _T_626 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13199.4]
  assign _T_628 = io_rPort_2_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13200.4]
  assign _T_629 = _T_626 & _T_628; // @[MemPrimitives.scala 110:228:@13201.4]
  assign _T_632 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13203.4]
  assign _T_634 = io_rPort_4_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13204.4]
  assign _T_635 = _T_632 & _T_634; // @[MemPrimitives.scala 110:228:@13205.4]
  assign _T_638 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13207.4]
  assign _T_640 = io_rPort_5_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13208.4]
  assign _T_641 = _T_638 & _T_640; // @[MemPrimitives.scala 110:228:@13209.4]
  assign _T_644 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13211.4]
  assign _T_646 = io_rPort_10_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13212.4]
  assign _T_647 = _T_644 & _T_646; // @[MemPrimitives.scala 110:228:@13213.4]
  assign _T_650 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13215.4]
  assign _T_652 = io_rPort_11_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13216.4]
  assign _T_653 = _T_650 & _T_652; // @[MemPrimitives.scala 110:228:@13217.4]
  assign _T_655 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@13228.4]
  assign _T_656 = StickySelects_io_outs_1; // @[MemPrimitives.scala 123:41:@13229.4]
  assign _T_657 = StickySelects_io_outs_2; // @[MemPrimitives.scala 123:41:@13230.4]
  assign _T_658 = StickySelects_io_outs_3; // @[MemPrimitives.scala 123:41:@13231.4]
  assign _T_659 = StickySelects_io_outs_4; // @[MemPrimitives.scala 123:41:@13232.4]
  assign _T_660 = StickySelects_io_outs_5; // @[MemPrimitives.scala 123:41:@13233.4]
  assign _T_662 = {_T_655,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13235.4]
  assign _T_664 = {_T_656,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13237.4]
  assign _T_666 = {_T_657,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13239.4]
  assign _T_668 = {_T_658,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13241.4]
  assign _T_670 = {_T_659,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13243.4]
  assign _T_672 = {_T_660,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13245.4]
  assign _T_673 = _T_659 ? _T_670 : _T_672; // @[Mux.scala 31:69:@13246.4]
  assign _T_674 = _T_658 ? _T_668 : _T_673; // @[Mux.scala 31:69:@13247.4]
  assign _T_675 = _T_657 ? _T_666 : _T_674; // @[Mux.scala 31:69:@13248.4]
  assign _T_676 = _T_656 ? _T_664 : _T_675; // @[Mux.scala 31:69:@13249.4]
  assign _T_677 = _T_655 ? _T_662 : _T_676; // @[Mux.scala 31:69:@13250.4]
  assign _T_682 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13257.4]
  assign _T_684 = io_rPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13258.4]
  assign _T_685 = _T_682 & _T_684; // @[MemPrimitives.scala 110:228:@13259.4]
  assign _T_688 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13261.4]
  assign _T_690 = io_rPort_3_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13262.4]
  assign _T_691 = _T_688 & _T_690; // @[MemPrimitives.scala 110:228:@13263.4]
  assign _T_694 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13265.4]
  assign _T_696 = io_rPort_6_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13266.4]
  assign _T_697 = _T_694 & _T_696; // @[MemPrimitives.scala 110:228:@13267.4]
  assign _T_700 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13269.4]
  assign _T_702 = io_rPort_7_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13270.4]
  assign _T_703 = _T_700 & _T_702; // @[MemPrimitives.scala 110:228:@13271.4]
  assign _T_706 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13273.4]
  assign _T_708 = io_rPort_8_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13274.4]
  assign _T_709 = _T_706 & _T_708; // @[MemPrimitives.scala 110:228:@13275.4]
  assign _T_712 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13277.4]
  assign _T_714 = io_rPort_9_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13278.4]
  assign _T_715 = _T_712 & _T_714; // @[MemPrimitives.scala 110:228:@13279.4]
  assign _T_717 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@13290.4]
  assign _T_718 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 123:41:@13291.4]
  assign _T_719 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 123:41:@13292.4]
  assign _T_720 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 123:41:@13293.4]
  assign _T_721 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 123:41:@13294.4]
  assign _T_722 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 123:41:@13295.4]
  assign _T_724 = {_T_717,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13297.4]
  assign _T_726 = {_T_718,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13299.4]
  assign _T_728 = {_T_719,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13301.4]
  assign _T_730 = {_T_720,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13303.4]
  assign _T_732 = {_T_721,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13305.4]
  assign _T_734 = {_T_722,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13307.4]
  assign _T_735 = _T_721 ? _T_732 : _T_734; // @[Mux.scala 31:69:@13308.4]
  assign _T_736 = _T_720 ? _T_730 : _T_735; // @[Mux.scala 31:69:@13309.4]
  assign _T_737 = _T_719 ? _T_728 : _T_736; // @[Mux.scala 31:69:@13310.4]
  assign _T_738 = _T_718 ? _T_726 : _T_737; // @[Mux.scala 31:69:@13311.4]
  assign _T_739 = _T_717 ? _T_724 : _T_738; // @[Mux.scala 31:69:@13312.4]
  assign _T_746 = io_rPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13320.4]
  assign _T_747 = _T_620 & _T_746; // @[MemPrimitives.scala 110:228:@13321.4]
  assign _T_752 = io_rPort_2_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13324.4]
  assign _T_753 = _T_626 & _T_752; // @[MemPrimitives.scala 110:228:@13325.4]
  assign _T_758 = io_rPort_4_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13328.4]
  assign _T_759 = _T_632 & _T_758; // @[MemPrimitives.scala 110:228:@13329.4]
  assign _T_764 = io_rPort_5_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13332.4]
  assign _T_765 = _T_638 & _T_764; // @[MemPrimitives.scala 110:228:@13333.4]
  assign _T_770 = io_rPort_10_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13336.4]
  assign _T_771 = _T_644 & _T_770; // @[MemPrimitives.scala 110:228:@13337.4]
  assign _T_776 = io_rPort_11_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13340.4]
  assign _T_777 = _T_650 & _T_776; // @[MemPrimitives.scala 110:228:@13341.4]
  assign _T_779 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@13352.4]
  assign _T_780 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 123:41:@13353.4]
  assign _T_781 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 123:41:@13354.4]
  assign _T_782 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 123:41:@13355.4]
  assign _T_783 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 123:41:@13356.4]
  assign _T_784 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 123:41:@13357.4]
  assign _T_786 = {_T_779,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13359.4]
  assign _T_788 = {_T_780,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13361.4]
  assign _T_790 = {_T_781,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13363.4]
  assign _T_792 = {_T_782,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13365.4]
  assign _T_794 = {_T_783,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13367.4]
  assign _T_796 = {_T_784,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13369.4]
  assign _T_797 = _T_783 ? _T_794 : _T_796; // @[Mux.scala 31:69:@13370.4]
  assign _T_798 = _T_782 ? _T_792 : _T_797; // @[Mux.scala 31:69:@13371.4]
  assign _T_799 = _T_781 ? _T_790 : _T_798; // @[Mux.scala 31:69:@13372.4]
  assign _T_800 = _T_780 ? _T_788 : _T_799; // @[Mux.scala 31:69:@13373.4]
  assign _T_801 = _T_779 ? _T_786 : _T_800; // @[Mux.scala 31:69:@13374.4]
  assign _T_808 = io_rPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13382.4]
  assign _T_809 = _T_682 & _T_808; // @[MemPrimitives.scala 110:228:@13383.4]
  assign _T_814 = io_rPort_3_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13386.4]
  assign _T_815 = _T_688 & _T_814; // @[MemPrimitives.scala 110:228:@13387.4]
  assign _T_820 = io_rPort_6_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13390.4]
  assign _T_821 = _T_694 & _T_820; // @[MemPrimitives.scala 110:228:@13391.4]
  assign _T_826 = io_rPort_7_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13394.4]
  assign _T_827 = _T_700 & _T_826; // @[MemPrimitives.scala 110:228:@13395.4]
  assign _T_832 = io_rPort_8_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13398.4]
  assign _T_833 = _T_706 & _T_832; // @[MemPrimitives.scala 110:228:@13399.4]
  assign _T_838 = io_rPort_9_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13402.4]
  assign _T_839 = _T_712 & _T_838; // @[MemPrimitives.scala 110:228:@13403.4]
  assign _T_841 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@13414.4]
  assign _T_842 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 123:41:@13415.4]
  assign _T_843 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 123:41:@13416.4]
  assign _T_844 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 123:41:@13417.4]
  assign _T_845 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 123:41:@13418.4]
  assign _T_846 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 123:41:@13419.4]
  assign _T_848 = {_T_841,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13421.4]
  assign _T_850 = {_T_842,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13423.4]
  assign _T_852 = {_T_843,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13425.4]
  assign _T_854 = {_T_844,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13427.4]
  assign _T_856 = {_T_845,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13429.4]
  assign _T_858 = {_T_846,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13431.4]
  assign _T_859 = _T_845 ? _T_856 : _T_858; // @[Mux.scala 31:69:@13432.4]
  assign _T_860 = _T_844 ? _T_854 : _T_859; // @[Mux.scala 31:69:@13433.4]
  assign _T_861 = _T_843 ? _T_852 : _T_860; // @[Mux.scala 31:69:@13434.4]
  assign _T_862 = _T_842 ? _T_850 : _T_861; // @[Mux.scala 31:69:@13435.4]
  assign _T_863 = _T_841 ? _T_848 : _T_862; // @[Mux.scala 31:69:@13436.4]
  assign _T_868 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13443.4]
  assign _T_871 = _T_868 & _T_622; // @[MemPrimitives.scala 110:228:@13445.4]
  assign _T_874 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13447.4]
  assign _T_877 = _T_874 & _T_628; // @[MemPrimitives.scala 110:228:@13449.4]
  assign _T_880 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13451.4]
  assign _T_883 = _T_880 & _T_634; // @[MemPrimitives.scala 110:228:@13453.4]
  assign _T_886 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13455.4]
  assign _T_889 = _T_886 & _T_640; // @[MemPrimitives.scala 110:228:@13457.4]
  assign _T_892 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13459.4]
  assign _T_895 = _T_892 & _T_646; // @[MemPrimitives.scala 110:228:@13461.4]
  assign _T_898 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13463.4]
  assign _T_901 = _T_898 & _T_652; // @[MemPrimitives.scala 110:228:@13465.4]
  assign _T_903 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@13476.4]
  assign _T_904 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 123:41:@13477.4]
  assign _T_905 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 123:41:@13478.4]
  assign _T_906 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 123:41:@13479.4]
  assign _T_907 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 123:41:@13480.4]
  assign _T_908 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 123:41:@13481.4]
  assign _T_910 = {_T_903,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13483.4]
  assign _T_912 = {_T_904,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13485.4]
  assign _T_914 = {_T_905,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13487.4]
  assign _T_916 = {_T_906,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13489.4]
  assign _T_918 = {_T_907,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13491.4]
  assign _T_920 = {_T_908,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13493.4]
  assign _T_921 = _T_907 ? _T_918 : _T_920; // @[Mux.scala 31:69:@13494.4]
  assign _T_922 = _T_906 ? _T_916 : _T_921; // @[Mux.scala 31:69:@13495.4]
  assign _T_923 = _T_905 ? _T_914 : _T_922; // @[Mux.scala 31:69:@13496.4]
  assign _T_924 = _T_904 ? _T_912 : _T_923; // @[Mux.scala 31:69:@13497.4]
  assign _T_925 = _T_903 ? _T_910 : _T_924; // @[Mux.scala 31:69:@13498.4]
  assign _T_930 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13505.4]
  assign _T_933 = _T_930 & _T_684; // @[MemPrimitives.scala 110:228:@13507.4]
  assign _T_936 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13509.4]
  assign _T_939 = _T_936 & _T_690; // @[MemPrimitives.scala 110:228:@13511.4]
  assign _T_942 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13513.4]
  assign _T_945 = _T_942 & _T_696; // @[MemPrimitives.scala 110:228:@13515.4]
  assign _T_948 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13517.4]
  assign _T_951 = _T_948 & _T_702; // @[MemPrimitives.scala 110:228:@13519.4]
  assign _T_954 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13521.4]
  assign _T_957 = _T_954 & _T_708; // @[MemPrimitives.scala 110:228:@13523.4]
  assign _T_960 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13525.4]
  assign _T_963 = _T_960 & _T_714; // @[MemPrimitives.scala 110:228:@13527.4]
  assign _T_965 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@13538.4]
  assign _T_966 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 123:41:@13539.4]
  assign _T_967 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 123:41:@13540.4]
  assign _T_968 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 123:41:@13541.4]
  assign _T_969 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 123:41:@13542.4]
  assign _T_970 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 123:41:@13543.4]
  assign _T_972 = {_T_965,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13545.4]
  assign _T_974 = {_T_966,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13547.4]
  assign _T_976 = {_T_967,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13549.4]
  assign _T_978 = {_T_968,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13551.4]
  assign _T_980 = {_T_969,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13553.4]
  assign _T_982 = {_T_970,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13555.4]
  assign _T_983 = _T_969 ? _T_980 : _T_982; // @[Mux.scala 31:69:@13556.4]
  assign _T_984 = _T_968 ? _T_978 : _T_983; // @[Mux.scala 31:69:@13557.4]
  assign _T_985 = _T_967 ? _T_976 : _T_984; // @[Mux.scala 31:69:@13558.4]
  assign _T_986 = _T_966 ? _T_974 : _T_985; // @[Mux.scala 31:69:@13559.4]
  assign _T_987 = _T_965 ? _T_972 : _T_986; // @[Mux.scala 31:69:@13560.4]
  assign _T_995 = _T_868 & _T_746; // @[MemPrimitives.scala 110:228:@13569.4]
  assign _T_1001 = _T_874 & _T_752; // @[MemPrimitives.scala 110:228:@13573.4]
  assign _T_1007 = _T_880 & _T_758; // @[MemPrimitives.scala 110:228:@13577.4]
  assign _T_1013 = _T_886 & _T_764; // @[MemPrimitives.scala 110:228:@13581.4]
  assign _T_1019 = _T_892 & _T_770; // @[MemPrimitives.scala 110:228:@13585.4]
  assign _T_1025 = _T_898 & _T_776; // @[MemPrimitives.scala 110:228:@13589.4]
  assign _T_1027 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@13600.4]
  assign _T_1028 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 123:41:@13601.4]
  assign _T_1029 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 123:41:@13602.4]
  assign _T_1030 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 123:41:@13603.4]
  assign _T_1031 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 123:41:@13604.4]
  assign _T_1032 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 123:41:@13605.4]
  assign _T_1034 = {_T_1027,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13607.4]
  assign _T_1036 = {_T_1028,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13609.4]
  assign _T_1038 = {_T_1029,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13611.4]
  assign _T_1040 = {_T_1030,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13613.4]
  assign _T_1042 = {_T_1031,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13615.4]
  assign _T_1044 = {_T_1032,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13617.4]
  assign _T_1045 = _T_1031 ? _T_1042 : _T_1044; // @[Mux.scala 31:69:@13618.4]
  assign _T_1046 = _T_1030 ? _T_1040 : _T_1045; // @[Mux.scala 31:69:@13619.4]
  assign _T_1047 = _T_1029 ? _T_1038 : _T_1046; // @[Mux.scala 31:69:@13620.4]
  assign _T_1048 = _T_1028 ? _T_1036 : _T_1047; // @[Mux.scala 31:69:@13621.4]
  assign _T_1049 = _T_1027 ? _T_1034 : _T_1048; // @[Mux.scala 31:69:@13622.4]
  assign _T_1057 = _T_930 & _T_808; // @[MemPrimitives.scala 110:228:@13631.4]
  assign _T_1063 = _T_936 & _T_814; // @[MemPrimitives.scala 110:228:@13635.4]
  assign _T_1069 = _T_942 & _T_820; // @[MemPrimitives.scala 110:228:@13639.4]
  assign _T_1075 = _T_948 & _T_826; // @[MemPrimitives.scala 110:228:@13643.4]
  assign _T_1081 = _T_954 & _T_832; // @[MemPrimitives.scala 110:228:@13647.4]
  assign _T_1087 = _T_960 & _T_838; // @[MemPrimitives.scala 110:228:@13651.4]
  assign _T_1089 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@13662.4]
  assign _T_1090 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 123:41:@13663.4]
  assign _T_1091 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 123:41:@13664.4]
  assign _T_1092 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 123:41:@13665.4]
  assign _T_1093 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 123:41:@13666.4]
  assign _T_1094 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 123:41:@13667.4]
  assign _T_1096 = {_T_1089,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13669.4]
  assign _T_1098 = {_T_1090,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13671.4]
  assign _T_1100 = {_T_1091,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13673.4]
  assign _T_1102 = {_T_1092,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13675.4]
  assign _T_1104 = {_T_1093,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13677.4]
  assign _T_1106 = {_T_1094,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13679.4]
  assign _T_1107 = _T_1093 ? _T_1104 : _T_1106; // @[Mux.scala 31:69:@13680.4]
  assign _T_1108 = _T_1092 ? _T_1102 : _T_1107; // @[Mux.scala 31:69:@13681.4]
  assign _T_1109 = _T_1091 ? _T_1100 : _T_1108; // @[Mux.scala 31:69:@13682.4]
  assign _T_1110 = _T_1090 ? _T_1098 : _T_1109; // @[Mux.scala 31:69:@13683.4]
  assign _T_1111 = _T_1089 ? _T_1096 : _T_1110; // @[Mux.scala 31:69:@13684.4]
  assign _T_1116 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13691.4]
  assign _T_1119 = _T_1116 & _T_622; // @[MemPrimitives.scala 110:228:@13693.4]
  assign _T_1122 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13695.4]
  assign _T_1125 = _T_1122 & _T_628; // @[MemPrimitives.scala 110:228:@13697.4]
  assign _T_1128 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13699.4]
  assign _T_1131 = _T_1128 & _T_634; // @[MemPrimitives.scala 110:228:@13701.4]
  assign _T_1134 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13703.4]
  assign _T_1137 = _T_1134 & _T_640; // @[MemPrimitives.scala 110:228:@13705.4]
  assign _T_1140 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13707.4]
  assign _T_1143 = _T_1140 & _T_646; // @[MemPrimitives.scala 110:228:@13709.4]
  assign _T_1146 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13711.4]
  assign _T_1149 = _T_1146 & _T_652; // @[MemPrimitives.scala 110:228:@13713.4]
  assign _T_1151 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@13724.4]
  assign _T_1152 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 123:41:@13725.4]
  assign _T_1153 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 123:41:@13726.4]
  assign _T_1154 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 123:41:@13727.4]
  assign _T_1155 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 123:41:@13728.4]
  assign _T_1156 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 123:41:@13729.4]
  assign _T_1158 = {_T_1151,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13731.4]
  assign _T_1160 = {_T_1152,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13733.4]
  assign _T_1162 = {_T_1153,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13735.4]
  assign _T_1164 = {_T_1154,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13737.4]
  assign _T_1166 = {_T_1155,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13739.4]
  assign _T_1168 = {_T_1156,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13741.4]
  assign _T_1169 = _T_1155 ? _T_1166 : _T_1168; // @[Mux.scala 31:69:@13742.4]
  assign _T_1170 = _T_1154 ? _T_1164 : _T_1169; // @[Mux.scala 31:69:@13743.4]
  assign _T_1171 = _T_1153 ? _T_1162 : _T_1170; // @[Mux.scala 31:69:@13744.4]
  assign _T_1172 = _T_1152 ? _T_1160 : _T_1171; // @[Mux.scala 31:69:@13745.4]
  assign _T_1173 = _T_1151 ? _T_1158 : _T_1172; // @[Mux.scala 31:69:@13746.4]
  assign _T_1178 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13753.4]
  assign _T_1181 = _T_1178 & _T_684; // @[MemPrimitives.scala 110:228:@13755.4]
  assign _T_1184 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13757.4]
  assign _T_1187 = _T_1184 & _T_690; // @[MemPrimitives.scala 110:228:@13759.4]
  assign _T_1190 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13761.4]
  assign _T_1193 = _T_1190 & _T_696; // @[MemPrimitives.scala 110:228:@13763.4]
  assign _T_1196 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13765.4]
  assign _T_1199 = _T_1196 & _T_702; // @[MemPrimitives.scala 110:228:@13767.4]
  assign _T_1202 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13769.4]
  assign _T_1205 = _T_1202 & _T_708; // @[MemPrimitives.scala 110:228:@13771.4]
  assign _T_1208 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13773.4]
  assign _T_1211 = _T_1208 & _T_714; // @[MemPrimitives.scala 110:228:@13775.4]
  assign _T_1213 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@13786.4]
  assign _T_1214 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 123:41:@13787.4]
  assign _T_1215 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 123:41:@13788.4]
  assign _T_1216 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 123:41:@13789.4]
  assign _T_1217 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 123:41:@13790.4]
  assign _T_1218 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 123:41:@13791.4]
  assign _T_1220 = {_T_1213,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13793.4]
  assign _T_1222 = {_T_1214,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13795.4]
  assign _T_1224 = {_T_1215,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13797.4]
  assign _T_1226 = {_T_1216,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13799.4]
  assign _T_1228 = {_T_1217,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13801.4]
  assign _T_1230 = {_T_1218,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13803.4]
  assign _T_1231 = _T_1217 ? _T_1228 : _T_1230; // @[Mux.scala 31:69:@13804.4]
  assign _T_1232 = _T_1216 ? _T_1226 : _T_1231; // @[Mux.scala 31:69:@13805.4]
  assign _T_1233 = _T_1215 ? _T_1224 : _T_1232; // @[Mux.scala 31:69:@13806.4]
  assign _T_1234 = _T_1214 ? _T_1222 : _T_1233; // @[Mux.scala 31:69:@13807.4]
  assign _T_1235 = _T_1213 ? _T_1220 : _T_1234; // @[Mux.scala 31:69:@13808.4]
  assign _T_1243 = _T_1116 & _T_746; // @[MemPrimitives.scala 110:228:@13817.4]
  assign _T_1249 = _T_1122 & _T_752; // @[MemPrimitives.scala 110:228:@13821.4]
  assign _T_1255 = _T_1128 & _T_758; // @[MemPrimitives.scala 110:228:@13825.4]
  assign _T_1261 = _T_1134 & _T_764; // @[MemPrimitives.scala 110:228:@13829.4]
  assign _T_1267 = _T_1140 & _T_770; // @[MemPrimitives.scala 110:228:@13833.4]
  assign _T_1273 = _T_1146 & _T_776; // @[MemPrimitives.scala 110:228:@13837.4]
  assign _T_1275 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@13848.4]
  assign _T_1276 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 123:41:@13849.4]
  assign _T_1277 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 123:41:@13850.4]
  assign _T_1278 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 123:41:@13851.4]
  assign _T_1279 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 123:41:@13852.4]
  assign _T_1280 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 123:41:@13853.4]
  assign _T_1282 = {_T_1275,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13855.4]
  assign _T_1284 = {_T_1276,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13857.4]
  assign _T_1286 = {_T_1277,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13859.4]
  assign _T_1288 = {_T_1278,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13861.4]
  assign _T_1290 = {_T_1279,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13863.4]
  assign _T_1292 = {_T_1280,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13865.4]
  assign _T_1293 = _T_1279 ? _T_1290 : _T_1292; // @[Mux.scala 31:69:@13866.4]
  assign _T_1294 = _T_1278 ? _T_1288 : _T_1293; // @[Mux.scala 31:69:@13867.4]
  assign _T_1295 = _T_1277 ? _T_1286 : _T_1294; // @[Mux.scala 31:69:@13868.4]
  assign _T_1296 = _T_1276 ? _T_1284 : _T_1295; // @[Mux.scala 31:69:@13869.4]
  assign _T_1297 = _T_1275 ? _T_1282 : _T_1296; // @[Mux.scala 31:69:@13870.4]
  assign _T_1305 = _T_1178 & _T_808; // @[MemPrimitives.scala 110:228:@13879.4]
  assign _T_1311 = _T_1184 & _T_814; // @[MemPrimitives.scala 110:228:@13883.4]
  assign _T_1317 = _T_1190 & _T_820; // @[MemPrimitives.scala 110:228:@13887.4]
  assign _T_1323 = _T_1196 & _T_826; // @[MemPrimitives.scala 110:228:@13891.4]
  assign _T_1329 = _T_1202 & _T_832; // @[MemPrimitives.scala 110:228:@13895.4]
  assign _T_1335 = _T_1208 & _T_838; // @[MemPrimitives.scala 110:228:@13899.4]
  assign _T_1337 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@13910.4]
  assign _T_1338 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 123:41:@13911.4]
  assign _T_1339 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 123:41:@13912.4]
  assign _T_1340 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 123:41:@13913.4]
  assign _T_1341 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 123:41:@13914.4]
  assign _T_1342 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 123:41:@13915.4]
  assign _T_1344 = {_T_1337,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13917.4]
  assign _T_1346 = {_T_1338,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13919.4]
  assign _T_1348 = {_T_1339,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13921.4]
  assign _T_1350 = {_T_1340,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13923.4]
  assign _T_1352 = {_T_1341,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13925.4]
  assign _T_1354 = {_T_1342,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13927.4]
  assign _T_1355 = _T_1341 ? _T_1352 : _T_1354; // @[Mux.scala 31:69:@13928.4]
  assign _T_1356 = _T_1340 ? _T_1350 : _T_1355; // @[Mux.scala 31:69:@13929.4]
  assign _T_1357 = _T_1339 ? _T_1348 : _T_1356; // @[Mux.scala 31:69:@13930.4]
  assign _T_1358 = _T_1338 ? _T_1346 : _T_1357; // @[Mux.scala 31:69:@13931.4]
  assign _T_1359 = _T_1337 ? _T_1344 : _T_1358; // @[Mux.scala 31:69:@13932.4]
  assign _T_1364 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13939.4]
  assign _T_1367 = _T_1364 & _T_622; // @[MemPrimitives.scala 110:228:@13941.4]
  assign _T_1370 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13943.4]
  assign _T_1373 = _T_1370 & _T_628; // @[MemPrimitives.scala 110:228:@13945.4]
  assign _T_1376 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13947.4]
  assign _T_1379 = _T_1376 & _T_634; // @[MemPrimitives.scala 110:228:@13949.4]
  assign _T_1382 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13951.4]
  assign _T_1385 = _T_1382 & _T_640; // @[MemPrimitives.scala 110:228:@13953.4]
  assign _T_1388 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13955.4]
  assign _T_1391 = _T_1388 & _T_646; // @[MemPrimitives.scala 110:228:@13957.4]
  assign _T_1394 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13959.4]
  assign _T_1397 = _T_1394 & _T_652; // @[MemPrimitives.scala 110:228:@13961.4]
  assign _T_1399 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 123:41:@13972.4]
  assign _T_1400 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 123:41:@13973.4]
  assign _T_1401 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 123:41:@13974.4]
  assign _T_1402 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 123:41:@13975.4]
  assign _T_1403 = StickySelects_12_io_outs_4; // @[MemPrimitives.scala 123:41:@13976.4]
  assign _T_1404 = StickySelects_12_io_outs_5; // @[MemPrimitives.scala 123:41:@13977.4]
  assign _T_1406 = {_T_1399,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13979.4]
  assign _T_1408 = {_T_1400,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13981.4]
  assign _T_1410 = {_T_1401,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13983.4]
  assign _T_1412 = {_T_1402,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13985.4]
  assign _T_1414 = {_T_1403,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13987.4]
  assign _T_1416 = {_T_1404,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13989.4]
  assign _T_1417 = _T_1403 ? _T_1414 : _T_1416; // @[Mux.scala 31:69:@13990.4]
  assign _T_1418 = _T_1402 ? _T_1412 : _T_1417; // @[Mux.scala 31:69:@13991.4]
  assign _T_1419 = _T_1401 ? _T_1410 : _T_1418; // @[Mux.scala 31:69:@13992.4]
  assign _T_1420 = _T_1400 ? _T_1408 : _T_1419; // @[Mux.scala 31:69:@13993.4]
  assign _T_1421 = _T_1399 ? _T_1406 : _T_1420; // @[Mux.scala 31:69:@13994.4]
  assign _T_1426 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14001.4]
  assign _T_1429 = _T_1426 & _T_684; // @[MemPrimitives.scala 110:228:@14003.4]
  assign _T_1432 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14005.4]
  assign _T_1435 = _T_1432 & _T_690; // @[MemPrimitives.scala 110:228:@14007.4]
  assign _T_1438 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14009.4]
  assign _T_1441 = _T_1438 & _T_696; // @[MemPrimitives.scala 110:228:@14011.4]
  assign _T_1444 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14013.4]
  assign _T_1447 = _T_1444 & _T_702; // @[MemPrimitives.scala 110:228:@14015.4]
  assign _T_1450 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14017.4]
  assign _T_1453 = _T_1450 & _T_708; // @[MemPrimitives.scala 110:228:@14019.4]
  assign _T_1456 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14021.4]
  assign _T_1459 = _T_1456 & _T_714; // @[MemPrimitives.scala 110:228:@14023.4]
  assign _T_1461 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 123:41:@14034.4]
  assign _T_1462 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 123:41:@14035.4]
  assign _T_1463 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 123:41:@14036.4]
  assign _T_1464 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 123:41:@14037.4]
  assign _T_1465 = StickySelects_13_io_outs_4; // @[MemPrimitives.scala 123:41:@14038.4]
  assign _T_1466 = StickySelects_13_io_outs_5; // @[MemPrimitives.scala 123:41:@14039.4]
  assign _T_1468 = {_T_1461,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@14041.4]
  assign _T_1470 = {_T_1462,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@14043.4]
  assign _T_1472 = {_T_1463,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@14045.4]
  assign _T_1474 = {_T_1464,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@14047.4]
  assign _T_1476 = {_T_1465,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@14049.4]
  assign _T_1478 = {_T_1466,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@14051.4]
  assign _T_1479 = _T_1465 ? _T_1476 : _T_1478; // @[Mux.scala 31:69:@14052.4]
  assign _T_1480 = _T_1464 ? _T_1474 : _T_1479; // @[Mux.scala 31:69:@14053.4]
  assign _T_1481 = _T_1463 ? _T_1472 : _T_1480; // @[Mux.scala 31:69:@14054.4]
  assign _T_1482 = _T_1462 ? _T_1470 : _T_1481; // @[Mux.scala 31:69:@14055.4]
  assign _T_1483 = _T_1461 ? _T_1468 : _T_1482; // @[Mux.scala 31:69:@14056.4]
  assign _T_1491 = _T_1364 & _T_746; // @[MemPrimitives.scala 110:228:@14065.4]
  assign _T_1497 = _T_1370 & _T_752; // @[MemPrimitives.scala 110:228:@14069.4]
  assign _T_1503 = _T_1376 & _T_758; // @[MemPrimitives.scala 110:228:@14073.4]
  assign _T_1509 = _T_1382 & _T_764; // @[MemPrimitives.scala 110:228:@14077.4]
  assign _T_1515 = _T_1388 & _T_770; // @[MemPrimitives.scala 110:228:@14081.4]
  assign _T_1521 = _T_1394 & _T_776; // @[MemPrimitives.scala 110:228:@14085.4]
  assign _T_1523 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 123:41:@14096.4]
  assign _T_1524 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 123:41:@14097.4]
  assign _T_1525 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 123:41:@14098.4]
  assign _T_1526 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 123:41:@14099.4]
  assign _T_1527 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 123:41:@14100.4]
  assign _T_1528 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 123:41:@14101.4]
  assign _T_1530 = {_T_1523,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@14103.4]
  assign _T_1532 = {_T_1524,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@14105.4]
  assign _T_1534 = {_T_1525,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@14107.4]
  assign _T_1536 = {_T_1526,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@14109.4]
  assign _T_1538 = {_T_1527,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@14111.4]
  assign _T_1540 = {_T_1528,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@14113.4]
  assign _T_1541 = _T_1527 ? _T_1538 : _T_1540; // @[Mux.scala 31:69:@14114.4]
  assign _T_1542 = _T_1526 ? _T_1536 : _T_1541; // @[Mux.scala 31:69:@14115.4]
  assign _T_1543 = _T_1525 ? _T_1534 : _T_1542; // @[Mux.scala 31:69:@14116.4]
  assign _T_1544 = _T_1524 ? _T_1532 : _T_1543; // @[Mux.scala 31:69:@14117.4]
  assign _T_1545 = _T_1523 ? _T_1530 : _T_1544; // @[Mux.scala 31:69:@14118.4]
  assign _T_1553 = _T_1426 & _T_808; // @[MemPrimitives.scala 110:228:@14127.4]
  assign _T_1559 = _T_1432 & _T_814; // @[MemPrimitives.scala 110:228:@14131.4]
  assign _T_1565 = _T_1438 & _T_820; // @[MemPrimitives.scala 110:228:@14135.4]
  assign _T_1571 = _T_1444 & _T_826; // @[MemPrimitives.scala 110:228:@14139.4]
  assign _T_1577 = _T_1450 & _T_832; // @[MemPrimitives.scala 110:228:@14143.4]
  assign _T_1583 = _T_1456 & _T_838; // @[MemPrimitives.scala 110:228:@14147.4]
  assign _T_1585 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 123:41:@14158.4]
  assign _T_1586 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 123:41:@14159.4]
  assign _T_1587 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 123:41:@14160.4]
  assign _T_1588 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 123:41:@14161.4]
  assign _T_1589 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 123:41:@14162.4]
  assign _T_1590 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 123:41:@14163.4]
  assign _T_1592 = {_T_1585,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@14165.4]
  assign _T_1594 = {_T_1586,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@14167.4]
  assign _T_1596 = {_T_1587,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@14169.4]
  assign _T_1598 = {_T_1588,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@14171.4]
  assign _T_1600 = {_T_1589,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@14173.4]
  assign _T_1602 = {_T_1590,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@14175.4]
  assign _T_1603 = _T_1589 ? _T_1600 : _T_1602; // @[Mux.scala 31:69:@14176.4]
  assign _T_1604 = _T_1588 ? _T_1598 : _T_1603; // @[Mux.scala 31:69:@14177.4]
  assign _T_1605 = _T_1587 ? _T_1596 : _T_1604; // @[Mux.scala 31:69:@14178.4]
  assign _T_1606 = _T_1586 ? _T_1594 : _T_1605; // @[Mux.scala 31:69:@14179.4]
  assign _T_1607 = _T_1585 ? _T_1592 : _T_1606; // @[Mux.scala 31:69:@14180.4]
  assign _T_1671 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@14265.4 package.scala 96:25:@14266.4]
  assign _T_1675 = _T_1671 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14275.4]
  assign _T_1668 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@14257.4 package.scala 96:25:@14258.4]
  assign _T_1676 = _T_1668 ? Mem1D_10_io_output : _T_1675; // @[Mux.scala 31:69:@14276.4]
  assign _T_1665 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@14249.4 package.scala 96:25:@14250.4]
  assign _T_1677 = _T_1665 ? Mem1D_8_io_output : _T_1676; // @[Mux.scala 31:69:@14277.4]
  assign _T_1662 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@14241.4 package.scala 96:25:@14242.4]
  assign _T_1678 = _T_1662 ? Mem1D_6_io_output : _T_1677; // @[Mux.scala 31:69:@14278.4]
  assign _T_1659 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@14233.4 package.scala 96:25:@14234.4]
  assign _T_1679 = _T_1659 ? Mem1D_4_io_output : _T_1678; // @[Mux.scala 31:69:@14279.4]
  assign _T_1656 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@14225.4 package.scala 96:25:@14226.4]
  assign _T_1680 = _T_1656 ? Mem1D_2_io_output : _T_1679; // @[Mux.scala 31:69:@14280.4]
  assign _T_1653 = RetimeWrapper_io_out; // @[package.scala 96:25:@14217.4 package.scala 96:25:@14218.4]
  assign _T_1742 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@14361.4 package.scala 96:25:@14362.4]
  assign _T_1746 = _T_1742 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14371.4]
  assign _T_1739 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@14353.4 package.scala 96:25:@14354.4]
  assign _T_1747 = _T_1739 ? Mem1D_11_io_output : _T_1746; // @[Mux.scala 31:69:@14372.4]
  assign _T_1736 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@14345.4 package.scala 96:25:@14346.4]
  assign _T_1748 = _T_1736 ? Mem1D_9_io_output : _T_1747; // @[Mux.scala 31:69:@14373.4]
  assign _T_1733 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@14337.4 package.scala 96:25:@14338.4]
  assign _T_1749 = _T_1733 ? Mem1D_7_io_output : _T_1748; // @[Mux.scala 31:69:@14374.4]
  assign _T_1730 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@14329.4 package.scala 96:25:@14330.4]
  assign _T_1750 = _T_1730 ? Mem1D_5_io_output : _T_1749; // @[Mux.scala 31:69:@14375.4]
  assign _T_1727 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@14321.4 package.scala 96:25:@14322.4]
  assign _T_1751 = _T_1727 ? Mem1D_3_io_output : _T_1750; // @[Mux.scala 31:69:@14376.4]
  assign _T_1724 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@14313.4 package.scala 96:25:@14314.4]
  assign _T_1813 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@14457.4 package.scala 96:25:@14458.4]
  assign _T_1817 = _T_1813 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14467.4]
  assign _T_1810 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@14449.4 package.scala 96:25:@14450.4]
  assign _T_1818 = _T_1810 ? Mem1D_10_io_output : _T_1817; // @[Mux.scala 31:69:@14468.4]
  assign _T_1807 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@14441.4 package.scala 96:25:@14442.4]
  assign _T_1819 = _T_1807 ? Mem1D_8_io_output : _T_1818; // @[Mux.scala 31:69:@14469.4]
  assign _T_1804 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@14433.4 package.scala 96:25:@14434.4]
  assign _T_1820 = _T_1804 ? Mem1D_6_io_output : _T_1819; // @[Mux.scala 31:69:@14470.4]
  assign _T_1801 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@14425.4 package.scala 96:25:@14426.4]
  assign _T_1821 = _T_1801 ? Mem1D_4_io_output : _T_1820; // @[Mux.scala 31:69:@14471.4]
  assign _T_1798 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@14417.4 package.scala 96:25:@14418.4]
  assign _T_1822 = _T_1798 ? Mem1D_2_io_output : _T_1821; // @[Mux.scala 31:69:@14472.4]
  assign _T_1795 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@14409.4 package.scala 96:25:@14410.4]
  assign _T_1884 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@14553.4 package.scala 96:25:@14554.4]
  assign _T_1888 = _T_1884 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14563.4]
  assign _T_1881 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@14545.4 package.scala 96:25:@14546.4]
  assign _T_1889 = _T_1881 ? Mem1D_11_io_output : _T_1888; // @[Mux.scala 31:69:@14564.4]
  assign _T_1878 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@14537.4 package.scala 96:25:@14538.4]
  assign _T_1890 = _T_1878 ? Mem1D_9_io_output : _T_1889; // @[Mux.scala 31:69:@14565.4]
  assign _T_1875 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@14529.4 package.scala 96:25:@14530.4]
  assign _T_1891 = _T_1875 ? Mem1D_7_io_output : _T_1890; // @[Mux.scala 31:69:@14566.4]
  assign _T_1872 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@14521.4 package.scala 96:25:@14522.4]
  assign _T_1892 = _T_1872 ? Mem1D_5_io_output : _T_1891; // @[Mux.scala 31:69:@14567.4]
  assign _T_1869 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@14513.4 package.scala 96:25:@14514.4]
  assign _T_1893 = _T_1869 ? Mem1D_3_io_output : _T_1892; // @[Mux.scala 31:69:@14568.4]
  assign _T_1866 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@14505.4 package.scala 96:25:@14506.4]
  assign _T_1955 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@14649.4 package.scala 96:25:@14650.4]
  assign _T_1959 = _T_1955 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14659.4]
  assign _T_1952 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@14641.4 package.scala 96:25:@14642.4]
  assign _T_1960 = _T_1952 ? Mem1D_10_io_output : _T_1959; // @[Mux.scala 31:69:@14660.4]
  assign _T_1949 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@14633.4 package.scala 96:25:@14634.4]
  assign _T_1961 = _T_1949 ? Mem1D_8_io_output : _T_1960; // @[Mux.scala 31:69:@14661.4]
  assign _T_1946 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@14625.4 package.scala 96:25:@14626.4]
  assign _T_1962 = _T_1946 ? Mem1D_6_io_output : _T_1961; // @[Mux.scala 31:69:@14662.4]
  assign _T_1943 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@14617.4 package.scala 96:25:@14618.4]
  assign _T_1963 = _T_1943 ? Mem1D_4_io_output : _T_1962; // @[Mux.scala 31:69:@14663.4]
  assign _T_1940 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@14609.4 package.scala 96:25:@14610.4]
  assign _T_1964 = _T_1940 ? Mem1D_2_io_output : _T_1963; // @[Mux.scala 31:69:@14664.4]
  assign _T_1937 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@14601.4 package.scala 96:25:@14602.4]
  assign _T_2026 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@14745.4 package.scala 96:25:@14746.4]
  assign _T_2030 = _T_2026 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14755.4]
  assign _T_2023 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@14737.4 package.scala 96:25:@14738.4]
  assign _T_2031 = _T_2023 ? Mem1D_10_io_output : _T_2030; // @[Mux.scala 31:69:@14756.4]
  assign _T_2020 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@14729.4 package.scala 96:25:@14730.4]
  assign _T_2032 = _T_2020 ? Mem1D_8_io_output : _T_2031; // @[Mux.scala 31:69:@14757.4]
  assign _T_2017 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@14721.4 package.scala 96:25:@14722.4]
  assign _T_2033 = _T_2017 ? Mem1D_6_io_output : _T_2032; // @[Mux.scala 31:69:@14758.4]
  assign _T_2014 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@14713.4 package.scala 96:25:@14714.4]
  assign _T_2034 = _T_2014 ? Mem1D_4_io_output : _T_2033; // @[Mux.scala 31:69:@14759.4]
  assign _T_2011 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@14705.4 package.scala 96:25:@14706.4]
  assign _T_2035 = _T_2011 ? Mem1D_2_io_output : _T_2034; // @[Mux.scala 31:69:@14760.4]
  assign _T_2008 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@14697.4 package.scala 96:25:@14698.4]
  assign _T_2097 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@14841.4 package.scala 96:25:@14842.4]
  assign _T_2101 = _T_2097 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14851.4]
  assign _T_2094 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@14833.4 package.scala 96:25:@14834.4]
  assign _T_2102 = _T_2094 ? Mem1D_11_io_output : _T_2101; // @[Mux.scala 31:69:@14852.4]
  assign _T_2091 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@14825.4 package.scala 96:25:@14826.4]
  assign _T_2103 = _T_2091 ? Mem1D_9_io_output : _T_2102; // @[Mux.scala 31:69:@14853.4]
  assign _T_2088 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@14817.4 package.scala 96:25:@14818.4]
  assign _T_2104 = _T_2088 ? Mem1D_7_io_output : _T_2103; // @[Mux.scala 31:69:@14854.4]
  assign _T_2085 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@14809.4 package.scala 96:25:@14810.4]
  assign _T_2105 = _T_2085 ? Mem1D_5_io_output : _T_2104; // @[Mux.scala 31:69:@14855.4]
  assign _T_2082 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@14801.4 package.scala 96:25:@14802.4]
  assign _T_2106 = _T_2082 ? Mem1D_3_io_output : _T_2105; // @[Mux.scala 31:69:@14856.4]
  assign _T_2079 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@14793.4 package.scala 96:25:@14794.4]
  assign _T_2168 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@14937.4 package.scala 96:25:@14938.4]
  assign _T_2172 = _T_2168 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14947.4]
  assign _T_2165 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@14929.4 package.scala 96:25:@14930.4]
  assign _T_2173 = _T_2165 ? Mem1D_11_io_output : _T_2172; // @[Mux.scala 31:69:@14948.4]
  assign _T_2162 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@14921.4 package.scala 96:25:@14922.4]
  assign _T_2174 = _T_2162 ? Mem1D_9_io_output : _T_2173; // @[Mux.scala 31:69:@14949.4]
  assign _T_2159 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@14913.4 package.scala 96:25:@14914.4]
  assign _T_2175 = _T_2159 ? Mem1D_7_io_output : _T_2174; // @[Mux.scala 31:69:@14950.4]
  assign _T_2156 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@14905.4 package.scala 96:25:@14906.4]
  assign _T_2176 = _T_2156 ? Mem1D_5_io_output : _T_2175; // @[Mux.scala 31:69:@14951.4]
  assign _T_2153 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@14897.4 package.scala 96:25:@14898.4]
  assign _T_2177 = _T_2153 ? Mem1D_3_io_output : _T_2176; // @[Mux.scala 31:69:@14952.4]
  assign _T_2150 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@14889.4 package.scala 96:25:@14890.4]
  assign _T_2239 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@15033.4 package.scala 96:25:@15034.4]
  assign _T_2243 = _T_2239 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@15043.4]
  assign _T_2236 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@15025.4 package.scala 96:25:@15026.4]
  assign _T_2244 = _T_2236 ? Mem1D_11_io_output : _T_2243; // @[Mux.scala 31:69:@15044.4]
  assign _T_2233 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@15017.4 package.scala 96:25:@15018.4]
  assign _T_2245 = _T_2233 ? Mem1D_9_io_output : _T_2244; // @[Mux.scala 31:69:@15045.4]
  assign _T_2230 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@15009.4 package.scala 96:25:@15010.4]
  assign _T_2246 = _T_2230 ? Mem1D_7_io_output : _T_2245; // @[Mux.scala 31:69:@15046.4]
  assign _T_2227 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@15001.4 package.scala 96:25:@15002.4]
  assign _T_2247 = _T_2227 ? Mem1D_5_io_output : _T_2246; // @[Mux.scala 31:69:@15047.4]
  assign _T_2224 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@14993.4 package.scala 96:25:@14994.4]
  assign _T_2248 = _T_2224 ? Mem1D_3_io_output : _T_2247; // @[Mux.scala 31:69:@15048.4]
  assign _T_2221 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@14985.4 package.scala 96:25:@14986.4]
  assign _T_2310 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@15129.4 package.scala 96:25:@15130.4]
  assign _T_2314 = _T_2310 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@15139.4]
  assign _T_2307 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@15121.4 package.scala 96:25:@15122.4]
  assign _T_2315 = _T_2307 ? Mem1D_11_io_output : _T_2314; // @[Mux.scala 31:69:@15140.4]
  assign _T_2304 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@15113.4 package.scala 96:25:@15114.4]
  assign _T_2316 = _T_2304 ? Mem1D_9_io_output : _T_2315; // @[Mux.scala 31:69:@15141.4]
  assign _T_2301 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@15105.4 package.scala 96:25:@15106.4]
  assign _T_2317 = _T_2301 ? Mem1D_7_io_output : _T_2316; // @[Mux.scala 31:69:@15142.4]
  assign _T_2298 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@15097.4 package.scala 96:25:@15098.4]
  assign _T_2318 = _T_2298 ? Mem1D_5_io_output : _T_2317; // @[Mux.scala 31:69:@15143.4]
  assign _T_2295 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@15089.4 package.scala 96:25:@15090.4]
  assign _T_2319 = _T_2295 ? Mem1D_3_io_output : _T_2318; // @[Mux.scala 31:69:@15144.4]
  assign _T_2292 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@15081.4 package.scala 96:25:@15082.4]
  assign _T_2381 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@15225.4 package.scala 96:25:@15226.4]
  assign _T_2385 = _T_2381 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@15235.4]
  assign _T_2378 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@15217.4 package.scala 96:25:@15218.4]
  assign _T_2386 = _T_2378 ? Mem1D_10_io_output : _T_2385; // @[Mux.scala 31:69:@15236.4]
  assign _T_2375 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@15209.4 package.scala 96:25:@15210.4]
  assign _T_2387 = _T_2375 ? Mem1D_8_io_output : _T_2386; // @[Mux.scala 31:69:@15237.4]
  assign _T_2372 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@15201.4 package.scala 96:25:@15202.4]
  assign _T_2388 = _T_2372 ? Mem1D_6_io_output : _T_2387; // @[Mux.scala 31:69:@15238.4]
  assign _T_2369 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@15193.4 package.scala 96:25:@15194.4]
  assign _T_2389 = _T_2369 ? Mem1D_4_io_output : _T_2388; // @[Mux.scala 31:69:@15239.4]
  assign _T_2366 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@15185.4 package.scala 96:25:@15186.4]
  assign _T_2390 = _T_2366 ? Mem1D_2_io_output : _T_2389; // @[Mux.scala 31:69:@15240.4]
  assign _T_2363 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@15177.4 package.scala 96:25:@15178.4]
  assign _T_2452 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@15321.4 package.scala 96:25:@15322.4]
  assign _T_2456 = _T_2452 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@15331.4]
  assign _T_2449 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@15313.4 package.scala 96:25:@15314.4]
  assign _T_2457 = _T_2449 ? Mem1D_10_io_output : _T_2456; // @[Mux.scala 31:69:@15332.4]
  assign _T_2446 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@15305.4 package.scala 96:25:@15306.4]
  assign _T_2458 = _T_2446 ? Mem1D_8_io_output : _T_2457; // @[Mux.scala 31:69:@15333.4]
  assign _T_2443 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@15297.4 package.scala 96:25:@15298.4]
  assign _T_2459 = _T_2443 ? Mem1D_6_io_output : _T_2458; // @[Mux.scala 31:69:@15334.4]
  assign _T_2440 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@15289.4 package.scala 96:25:@15290.4]
  assign _T_2460 = _T_2440 ? Mem1D_4_io_output : _T_2459; // @[Mux.scala 31:69:@15335.4]
  assign _T_2437 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@15281.4 package.scala 96:25:@15282.4]
  assign _T_2461 = _T_2437 ? Mem1D_2_io_output : _T_2460; // @[Mux.scala 31:69:@15336.4]
  assign _T_2434 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@15273.4 package.scala 96:25:@15274.4]
  assign io_rPort_11_output_0 = _T_2434 ? Mem1D_io_output : _T_2461; // @[MemPrimitives.scala 148:13:@15338.4]
  assign io_rPort_10_output_0 = _T_2363 ? Mem1D_io_output : _T_2390; // @[MemPrimitives.scala 148:13:@15242.4]
  assign io_rPort_9_output_0 = _T_2292 ? Mem1D_1_io_output : _T_2319; // @[MemPrimitives.scala 148:13:@15146.4]
  assign io_rPort_8_output_0 = _T_2221 ? Mem1D_1_io_output : _T_2248; // @[MemPrimitives.scala 148:13:@15050.4]
  assign io_rPort_7_output_0 = _T_2150 ? Mem1D_1_io_output : _T_2177; // @[MemPrimitives.scala 148:13:@14954.4]
  assign io_rPort_6_output_0 = _T_2079 ? Mem1D_1_io_output : _T_2106; // @[MemPrimitives.scala 148:13:@14858.4]
  assign io_rPort_5_output_0 = _T_2008 ? Mem1D_io_output : _T_2035; // @[MemPrimitives.scala 148:13:@14762.4]
  assign io_rPort_4_output_0 = _T_1937 ? Mem1D_io_output : _T_1964; // @[MemPrimitives.scala 148:13:@14666.4]
  assign io_rPort_3_output_0 = _T_1866 ? Mem1D_1_io_output : _T_1893; // @[MemPrimitives.scala 148:13:@14570.4]
  assign io_rPort_2_output_0 = _T_1795 ? Mem1D_io_output : _T_1822; // @[MemPrimitives.scala 148:13:@14474.4]
  assign io_rPort_1_output_0 = _T_1724 ? Mem1D_1_io_output : _T_1751; // @[MemPrimitives.scala 148:13:@14378.4]
  assign io_rPort_0_output_0 = _T_1653 ? Mem1D_io_output : _T_1680; // @[MemPrimitives.scala 148:13:@14282.4]
  assign Mem1D_clock = clock; // @[:@12748.4]
  assign Mem1D_reset = reset; // @[:@12749.4]
  assign Mem1D_io_r_ofs_0 = _T_677[8:0]; // @[MemPrimitives.scala 127:28:@13254.4]
  assign Mem1D_io_r_backpressure = _T_677[9]; // @[MemPrimitives.scala 128:32:@13255.4]
  assign Mem1D_io_w_ofs_0 = _T_450[8:0]; // @[MemPrimitives.scala 94:28:@13012.4]
  assign Mem1D_io_w_data_0 = _T_450[16:9]; // @[MemPrimitives.scala 95:29:@13013.4]
  assign Mem1D_io_w_en_0 = _T_450[17]; // @[MemPrimitives.scala 96:27:@13014.4]
  assign Mem1D_1_clock = clock; // @[:@12764.4]
  assign Mem1D_1_reset = reset; // @[:@12765.4]
  assign Mem1D_1_io_r_ofs_0 = _T_739[8:0]; // @[MemPrimitives.scala 127:28:@13316.4]
  assign Mem1D_1_io_r_backpressure = _T_739[9]; // @[MemPrimitives.scala 128:32:@13317.4]
  assign Mem1D_1_io_w_ofs_0 = _T_461[8:0]; // @[MemPrimitives.scala 94:28:@13024.4]
  assign Mem1D_1_io_w_data_0 = _T_461[16:9]; // @[MemPrimitives.scala 95:29:@13025.4]
  assign Mem1D_1_io_w_en_0 = _T_461[17]; // @[MemPrimitives.scala 96:27:@13026.4]
  assign Mem1D_2_clock = clock; // @[:@12780.4]
  assign Mem1D_2_reset = reset; // @[:@12781.4]
  assign Mem1D_2_io_r_ofs_0 = _T_801[8:0]; // @[MemPrimitives.scala 127:28:@13378.4]
  assign Mem1D_2_io_r_backpressure = _T_801[9]; // @[MemPrimitives.scala 128:32:@13379.4]
  assign Mem1D_2_io_w_ofs_0 = _T_472[8:0]; // @[MemPrimitives.scala 94:28:@13036.4]
  assign Mem1D_2_io_w_data_0 = _T_472[16:9]; // @[MemPrimitives.scala 95:29:@13037.4]
  assign Mem1D_2_io_w_en_0 = _T_472[17]; // @[MemPrimitives.scala 96:27:@13038.4]
  assign Mem1D_3_clock = clock; // @[:@12796.4]
  assign Mem1D_3_reset = reset; // @[:@12797.4]
  assign Mem1D_3_io_r_ofs_0 = _T_863[8:0]; // @[MemPrimitives.scala 127:28:@13440.4]
  assign Mem1D_3_io_r_backpressure = _T_863[9]; // @[MemPrimitives.scala 128:32:@13441.4]
  assign Mem1D_3_io_w_ofs_0 = _T_483[8:0]; // @[MemPrimitives.scala 94:28:@13048.4]
  assign Mem1D_3_io_w_data_0 = _T_483[16:9]; // @[MemPrimitives.scala 95:29:@13049.4]
  assign Mem1D_3_io_w_en_0 = _T_483[17]; // @[MemPrimitives.scala 96:27:@13050.4]
  assign Mem1D_4_clock = clock; // @[:@12812.4]
  assign Mem1D_4_reset = reset; // @[:@12813.4]
  assign Mem1D_4_io_r_ofs_0 = _T_925[8:0]; // @[MemPrimitives.scala 127:28:@13502.4]
  assign Mem1D_4_io_r_backpressure = _T_925[9]; // @[MemPrimitives.scala 128:32:@13503.4]
  assign Mem1D_4_io_w_ofs_0 = _T_494[8:0]; // @[MemPrimitives.scala 94:28:@13060.4]
  assign Mem1D_4_io_w_data_0 = _T_494[16:9]; // @[MemPrimitives.scala 95:29:@13061.4]
  assign Mem1D_4_io_w_en_0 = _T_494[17]; // @[MemPrimitives.scala 96:27:@13062.4]
  assign Mem1D_5_clock = clock; // @[:@12828.4]
  assign Mem1D_5_reset = reset; // @[:@12829.4]
  assign Mem1D_5_io_r_ofs_0 = _T_987[8:0]; // @[MemPrimitives.scala 127:28:@13564.4]
  assign Mem1D_5_io_r_backpressure = _T_987[9]; // @[MemPrimitives.scala 128:32:@13565.4]
  assign Mem1D_5_io_w_ofs_0 = _T_505[8:0]; // @[MemPrimitives.scala 94:28:@13072.4]
  assign Mem1D_5_io_w_data_0 = _T_505[16:9]; // @[MemPrimitives.scala 95:29:@13073.4]
  assign Mem1D_5_io_w_en_0 = _T_505[17]; // @[MemPrimitives.scala 96:27:@13074.4]
  assign Mem1D_6_clock = clock; // @[:@12844.4]
  assign Mem1D_6_reset = reset; // @[:@12845.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1049[8:0]; // @[MemPrimitives.scala 127:28:@13626.4]
  assign Mem1D_6_io_r_backpressure = _T_1049[9]; // @[MemPrimitives.scala 128:32:@13627.4]
  assign Mem1D_6_io_w_ofs_0 = _T_516[8:0]; // @[MemPrimitives.scala 94:28:@13084.4]
  assign Mem1D_6_io_w_data_0 = _T_516[16:9]; // @[MemPrimitives.scala 95:29:@13085.4]
  assign Mem1D_6_io_w_en_0 = _T_516[17]; // @[MemPrimitives.scala 96:27:@13086.4]
  assign Mem1D_7_clock = clock; // @[:@12860.4]
  assign Mem1D_7_reset = reset; // @[:@12861.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1111[8:0]; // @[MemPrimitives.scala 127:28:@13688.4]
  assign Mem1D_7_io_r_backpressure = _T_1111[9]; // @[MemPrimitives.scala 128:32:@13689.4]
  assign Mem1D_7_io_w_ofs_0 = _T_527[8:0]; // @[MemPrimitives.scala 94:28:@13096.4]
  assign Mem1D_7_io_w_data_0 = _T_527[16:9]; // @[MemPrimitives.scala 95:29:@13097.4]
  assign Mem1D_7_io_w_en_0 = _T_527[17]; // @[MemPrimitives.scala 96:27:@13098.4]
  assign Mem1D_8_clock = clock; // @[:@12876.4]
  assign Mem1D_8_reset = reset; // @[:@12877.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1173[8:0]; // @[MemPrimitives.scala 127:28:@13750.4]
  assign Mem1D_8_io_r_backpressure = _T_1173[9]; // @[MemPrimitives.scala 128:32:@13751.4]
  assign Mem1D_8_io_w_ofs_0 = _T_538[8:0]; // @[MemPrimitives.scala 94:28:@13108.4]
  assign Mem1D_8_io_w_data_0 = _T_538[16:9]; // @[MemPrimitives.scala 95:29:@13109.4]
  assign Mem1D_8_io_w_en_0 = _T_538[17]; // @[MemPrimitives.scala 96:27:@13110.4]
  assign Mem1D_9_clock = clock; // @[:@12892.4]
  assign Mem1D_9_reset = reset; // @[:@12893.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1235[8:0]; // @[MemPrimitives.scala 127:28:@13812.4]
  assign Mem1D_9_io_r_backpressure = _T_1235[9]; // @[MemPrimitives.scala 128:32:@13813.4]
  assign Mem1D_9_io_w_ofs_0 = _T_549[8:0]; // @[MemPrimitives.scala 94:28:@13120.4]
  assign Mem1D_9_io_w_data_0 = _T_549[16:9]; // @[MemPrimitives.scala 95:29:@13121.4]
  assign Mem1D_9_io_w_en_0 = _T_549[17]; // @[MemPrimitives.scala 96:27:@13122.4]
  assign Mem1D_10_clock = clock; // @[:@12908.4]
  assign Mem1D_10_reset = reset; // @[:@12909.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1297[8:0]; // @[MemPrimitives.scala 127:28:@13874.4]
  assign Mem1D_10_io_r_backpressure = _T_1297[9]; // @[MemPrimitives.scala 128:32:@13875.4]
  assign Mem1D_10_io_w_ofs_0 = _T_560[8:0]; // @[MemPrimitives.scala 94:28:@13132.4]
  assign Mem1D_10_io_w_data_0 = _T_560[16:9]; // @[MemPrimitives.scala 95:29:@13133.4]
  assign Mem1D_10_io_w_en_0 = _T_560[17]; // @[MemPrimitives.scala 96:27:@13134.4]
  assign Mem1D_11_clock = clock; // @[:@12924.4]
  assign Mem1D_11_reset = reset; // @[:@12925.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1359[8:0]; // @[MemPrimitives.scala 127:28:@13936.4]
  assign Mem1D_11_io_r_backpressure = _T_1359[9]; // @[MemPrimitives.scala 128:32:@13937.4]
  assign Mem1D_11_io_w_ofs_0 = _T_571[8:0]; // @[MemPrimitives.scala 94:28:@13144.4]
  assign Mem1D_11_io_w_data_0 = _T_571[16:9]; // @[MemPrimitives.scala 95:29:@13145.4]
  assign Mem1D_11_io_w_en_0 = _T_571[17]; // @[MemPrimitives.scala 96:27:@13146.4]
  assign Mem1D_12_clock = clock; // @[:@12940.4]
  assign Mem1D_12_reset = reset; // @[:@12941.4]
  assign Mem1D_12_io_r_ofs_0 = _T_1421[8:0]; // @[MemPrimitives.scala 127:28:@13998.4]
  assign Mem1D_12_io_r_backpressure = _T_1421[9]; // @[MemPrimitives.scala 128:32:@13999.4]
  assign Mem1D_12_io_w_ofs_0 = _T_582[8:0]; // @[MemPrimitives.scala 94:28:@13156.4]
  assign Mem1D_12_io_w_data_0 = _T_582[16:9]; // @[MemPrimitives.scala 95:29:@13157.4]
  assign Mem1D_12_io_w_en_0 = _T_582[17]; // @[MemPrimitives.scala 96:27:@13158.4]
  assign Mem1D_13_clock = clock; // @[:@12956.4]
  assign Mem1D_13_reset = reset; // @[:@12957.4]
  assign Mem1D_13_io_r_ofs_0 = _T_1483[8:0]; // @[MemPrimitives.scala 127:28:@14060.4]
  assign Mem1D_13_io_r_backpressure = _T_1483[9]; // @[MemPrimitives.scala 128:32:@14061.4]
  assign Mem1D_13_io_w_ofs_0 = _T_593[8:0]; // @[MemPrimitives.scala 94:28:@13168.4]
  assign Mem1D_13_io_w_data_0 = _T_593[16:9]; // @[MemPrimitives.scala 95:29:@13169.4]
  assign Mem1D_13_io_w_en_0 = _T_593[17]; // @[MemPrimitives.scala 96:27:@13170.4]
  assign Mem1D_14_clock = clock; // @[:@12972.4]
  assign Mem1D_14_reset = reset; // @[:@12973.4]
  assign Mem1D_14_io_r_ofs_0 = _T_1545[8:0]; // @[MemPrimitives.scala 127:28:@14122.4]
  assign Mem1D_14_io_r_backpressure = _T_1545[9]; // @[MemPrimitives.scala 128:32:@14123.4]
  assign Mem1D_14_io_w_ofs_0 = _T_604[8:0]; // @[MemPrimitives.scala 94:28:@13180.4]
  assign Mem1D_14_io_w_data_0 = _T_604[16:9]; // @[MemPrimitives.scala 95:29:@13181.4]
  assign Mem1D_14_io_w_en_0 = _T_604[17]; // @[MemPrimitives.scala 96:27:@13182.4]
  assign Mem1D_15_clock = clock; // @[:@12988.4]
  assign Mem1D_15_reset = reset; // @[:@12989.4]
  assign Mem1D_15_io_r_ofs_0 = _T_1607[8:0]; // @[MemPrimitives.scala 127:28:@14184.4]
  assign Mem1D_15_io_r_backpressure = _T_1607[9]; // @[MemPrimitives.scala 128:32:@14185.4]
  assign Mem1D_15_io_w_ofs_0 = _T_615[8:0]; // @[MemPrimitives.scala 94:28:@13192.4]
  assign Mem1D_15_io_w_data_0 = _T_615[16:9]; // @[MemPrimitives.scala 95:29:@13193.4]
  assign Mem1D_15_io_w_en_0 = _T_615[17]; // @[MemPrimitives.scala 96:27:@13194.4]
  assign StickySelects_clock = clock; // @[:@13220.4]
  assign StickySelects_reset = reset; // @[:@13221.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_623; // @[MemPrimitives.scala 122:60:@13222.4]
  assign StickySelects_io_ins_1 = io_rPort_2_en_0 & _T_629; // @[MemPrimitives.scala 122:60:@13223.4]
  assign StickySelects_io_ins_2 = io_rPort_4_en_0 & _T_635; // @[MemPrimitives.scala 122:60:@13224.4]
  assign StickySelects_io_ins_3 = io_rPort_5_en_0 & _T_641; // @[MemPrimitives.scala 122:60:@13225.4]
  assign StickySelects_io_ins_4 = io_rPort_10_en_0 & _T_647; // @[MemPrimitives.scala 122:60:@13226.4]
  assign StickySelects_io_ins_5 = io_rPort_11_en_0 & _T_653; // @[MemPrimitives.scala 122:60:@13227.4]
  assign StickySelects_1_clock = clock; // @[:@13282.4]
  assign StickySelects_1_reset = reset; // @[:@13283.4]
  assign StickySelects_1_io_ins_0 = io_rPort_1_en_0 & _T_685; // @[MemPrimitives.scala 122:60:@13284.4]
  assign StickySelects_1_io_ins_1 = io_rPort_3_en_0 & _T_691; // @[MemPrimitives.scala 122:60:@13285.4]
  assign StickySelects_1_io_ins_2 = io_rPort_6_en_0 & _T_697; // @[MemPrimitives.scala 122:60:@13286.4]
  assign StickySelects_1_io_ins_3 = io_rPort_7_en_0 & _T_703; // @[MemPrimitives.scala 122:60:@13287.4]
  assign StickySelects_1_io_ins_4 = io_rPort_8_en_0 & _T_709; // @[MemPrimitives.scala 122:60:@13288.4]
  assign StickySelects_1_io_ins_5 = io_rPort_9_en_0 & _T_715; // @[MemPrimitives.scala 122:60:@13289.4]
  assign StickySelects_2_clock = clock; // @[:@13344.4]
  assign StickySelects_2_reset = reset; // @[:@13345.4]
  assign StickySelects_2_io_ins_0 = io_rPort_0_en_0 & _T_747; // @[MemPrimitives.scala 122:60:@13346.4]
  assign StickySelects_2_io_ins_1 = io_rPort_2_en_0 & _T_753; // @[MemPrimitives.scala 122:60:@13347.4]
  assign StickySelects_2_io_ins_2 = io_rPort_4_en_0 & _T_759; // @[MemPrimitives.scala 122:60:@13348.4]
  assign StickySelects_2_io_ins_3 = io_rPort_5_en_0 & _T_765; // @[MemPrimitives.scala 122:60:@13349.4]
  assign StickySelects_2_io_ins_4 = io_rPort_10_en_0 & _T_771; // @[MemPrimitives.scala 122:60:@13350.4]
  assign StickySelects_2_io_ins_5 = io_rPort_11_en_0 & _T_777; // @[MemPrimitives.scala 122:60:@13351.4]
  assign StickySelects_3_clock = clock; // @[:@13406.4]
  assign StickySelects_3_reset = reset; // @[:@13407.4]
  assign StickySelects_3_io_ins_0 = io_rPort_1_en_0 & _T_809; // @[MemPrimitives.scala 122:60:@13408.4]
  assign StickySelects_3_io_ins_1 = io_rPort_3_en_0 & _T_815; // @[MemPrimitives.scala 122:60:@13409.4]
  assign StickySelects_3_io_ins_2 = io_rPort_6_en_0 & _T_821; // @[MemPrimitives.scala 122:60:@13410.4]
  assign StickySelects_3_io_ins_3 = io_rPort_7_en_0 & _T_827; // @[MemPrimitives.scala 122:60:@13411.4]
  assign StickySelects_3_io_ins_4 = io_rPort_8_en_0 & _T_833; // @[MemPrimitives.scala 122:60:@13412.4]
  assign StickySelects_3_io_ins_5 = io_rPort_9_en_0 & _T_839; // @[MemPrimitives.scala 122:60:@13413.4]
  assign StickySelects_4_clock = clock; // @[:@13468.4]
  assign StickySelects_4_reset = reset; // @[:@13469.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_871; // @[MemPrimitives.scala 122:60:@13470.4]
  assign StickySelects_4_io_ins_1 = io_rPort_2_en_0 & _T_877; // @[MemPrimitives.scala 122:60:@13471.4]
  assign StickySelects_4_io_ins_2 = io_rPort_4_en_0 & _T_883; // @[MemPrimitives.scala 122:60:@13472.4]
  assign StickySelects_4_io_ins_3 = io_rPort_5_en_0 & _T_889; // @[MemPrimitives.scala 122:60:@13473.4]
  assign StickySelects_4_io_ins_4 = io_rPort_10_en_0 & _T_895; // @[MemPrimitives.scala 122:60:@13474.4]
  assign StickySelects_4_io_ins_5 = io_rPort_11_en_0 & _T_901; // @[MemPrimitives.scala 122:60:@13475.4]
  assign StickySelects_5_clock = clock; // @[:@13530.4]
  assign StickySelects_5_reset = reset; // @[:@13531.4]
  assign StickySelects_5_io_ins_0 = io_rPort_1_en_0 & _T_933; // @[MemPrimitives.scala 122:60:@13532.4]
  assign StickySelects_5_io_ins_1 = io_rPort_3_en_0 & _T_939; // @[MemPrimitives.scala 122:60:@13533.4]
  assign StickySelects_5_io_ins_2 = io_rPort_6_en_0 & _T_945; // @[MemPrimitives.scala 122:60:@13534.4]
  assign StickySelects_5_io_ins_3 = io_rPort_7_en_0 & _T_951; // @[MemPrimitives.scala 122:60:@13535.4]
  assign StickySelects_5_io_ins_4 = io_rPort_8_en_0 & _T_957; // @[MemPrimitives.scala 122:60:@13536.4]
  assign StickySelects_5_io_ins_5 = io_rPort_9_en_0 & _T_963; // @[MemPrimitives.scala 122:60:@13537.4]
  assign StickySelects_6_clock = clock; // @[:@13592.4]
  assign StickySelects_6_reset = reset; // @[:@13593.4]
  assign StickySelects_6_io_ins_0 = io_rPort_0_en_0 & _T_995; // @[MemPrimitives.scala 122:60:@13594.4]
  assign StickySelects_6_io_ins_1 = io_rPort_2_en_0 & _T_1001; // @[MemPrimitives.scala 122:60:@13595.4]
  assign StickySelects_6_io_ins_2 = io_rPort_4_en_0 & _T_1007; // @[MemPrimitives.scala 122:60:@13596.4]
  assign StickySelects_6_io_ins_3 = io_rPort_5_en_0 & _T_1013; // @[MemPrimitives.scala 122:60:@13597.4]
  assign StickySelects_6_io_ins_4 = io_rPort_10_en_0 & _T_1019; // @[MemPrimitives.scala 122:60:@13598.4]
  assign StickySelects_6_io_ins_5 = io_rPort_11_en_0 & _T_1025; // @[MemPrimitives.scala 122:60:@13599.4]
  assign StickySelects_7_clock = clock; // @[:@13654.4]
  assign StickySelects_7_reset = reset; // @[:@13655.4]
  assign StickySelects_7_io_ins_0 = io_rPort_1_en_0 & _T_1057; // @[MemPrimitives.scala 122:60:@13656.4]
  assign StickySelects_7_io_ins_1 = io_rPort_3_en_0 & _T_1063; // @[MemPrimitives.scala 122:60:@13657.4]
  assign StickySelects_7_io_ins_2 = io_rPort_6_en_0 & _T_1069; // @[MemPrimitives.scala 122:60:@13658.4]
  assign StickySelects_7_io_ins_3 = io_rPort_7_en_0 & _T_1075; // @[MemPrimitives.scala 122:60:@13659.4]
  assign StickySelects_7_io_ins_4 = io_rPort_8_en_0 & _T_1081; // @[MemPrimitives.scala 122:60:@13660.4]
  assign StickySelects_7_io_ins_5 = io_rPort_9_en_0 & _T_1087; // @[MemPrimitives.scala 122:60:@13661.4]
  assign StickySelects_8_clock = clock; // @[:@13716.4]
  assign StickySelects_8_reset = reset; // @[:@13717.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_1119; // @[MemPrimitives.scala 122:60:@13718.4]
  assign StickySelects_8_io_ins_1 = io_rPort_2_en_0 & _T_1125; // @[MemPrimitives.scala 122:60:@13719.4]
  assign StickySelects_8_io_ins_2 = io_rPort_4_en_0 & _T_1131; // @[MemPrimitives.scala 122:60:@13720.4]
  assign StickySelects_8_io_ins_3 = io_rPort_5_en_0 & _T_1137; // @[MemPrimitives.scala 122:60:@13721.4]
  assign StickySelects_8_io_ins_4 = io_rPort_10_en_0 & _T_1143; // @[MemPrimitives.scala 122:60:@13722.4]
  assign StickySelects_8_io_ins_5 = io_rPort_11_en_0 & _T_1149; // @[MemPrimitives.scala 122:60:@13723.4]
  assign StickySelects_9_clock = clock; // @[:@13778.4]
  assign StickySelects_9_reset = reset; // @[:@13779.4]
  assign StickySelects_9_io_ins_0 = io_rPort_1_en_0 & _T_1181; // @[MemPrimitives.scala 122:60:@13780.4]
  assign StickySelects_9_io_ins_1 = io_rPort_3_en_0 & _T_1187; // @[MemPrimitives.scala 122:60:@13781.4]
  assign StickySelects_9_io_ins_2 = io_rPort_6_en_0 & _T_1193; // @[MemPrimitives.scala 122:60:@13782.4]
  assign StickySelects_9_io_ins_3 = io_rPort_7_en_0 & _T_1199; // @[MemPrimitives.scala 122:60:@13783.4]
  assign StickySelects_9_io_ins_4 = io_rPort_8_en_0 & _T_1205; // @[MemPrimitives.scala 122:60:@13784.4]
  assign StickySelects_9_io_ins_5 = io_rPort_9_en_0 & _T_1211; // @[MemPrimitives.scala 122:60:@13785.4]
  assign StickySelects_10_clock = clock; // @[:@13840.4]
  assign StickySelects_10_reset = reset; // @[:@13841.4]
  assign StickySelects_10_io_ins_0 = io_rPort_0_en_0 & _T_1243; // @[MemPrimitives.scala 122:60:@13842.4]
  assign StickySelects_10_io_ins_1 = io_rPort_2_en_0 & _T_1249; // @[MemPrimitives.scala 122:60:@13843.4]
  assign StickySelects_10_io_ins_2 = io_rPort_4_en_0 & _T_1255; // @[MemPrimitives.scala 122:60:@13844.4]
  assign StickySelects_10_io_ins_3 = io_rPort_5_en_0 & _T_1261; // @[MemPrimitives.scala 122:60:@13845.4]
  assign StickySelects_10_io_ins_4 = io_rPort_10_en_0 & _T_1267; // @[MemPrimitives.scala 122:60:@13846.4]
  assign StickySelects_10_io_ins_5 = io_rPort_11_en_0 & _T_1273; // @[MemPrimitives.scala 122:60:@13847.4]
  assign StickySelects_11_clock = clock; // @[:@13902.4]
  assign StickySelects_11_reset = reset; // @[:@13903.4]
  assign StickySelects_11_io_ins_0 = io_rPort_1_en_0 & _T_1305; // @[MemPrimitives.scala 122:60:@13904.4]
  assign StickySelects_11_io_ins_1 = io_rPort_3_en_0 & _T_1311; // @[MemPrimitives.scala 122:60:@13905.4]
  assign StickySelects_11_io_ins_2 = io_rPort_6_en_0 & _T_1317; // @[MemPrimitives.scala 122:60:@13906.4]
  assign StickySelects_11_io_ins_3 = io_rPort_7_en_0 & _T_1323; // @[MemPrimitives.scala 122:60:@13907.4]
  assign StickySelects_11_io_ins_4 = io_rPort_8_en_0 & _T_1329; // @[MemPrimitives.scala 122:60:@13908.4]
  assign StickySelects_11_io_ins_5 = io_rPort_9_en_0 & _T_1335; // @[MemPrimitives.scala 122:60:@13909.4]
  assign StickySelects_12_clock = clock; // @[:@13964.4]
  assign StickySelects_12_reset = reset; // @[:@13965.4]
  assign StickySelects_12_io_ins_0 = io_rPort_0_en_0 & _T_1367; // @[MemPrimitives.scala 122:60:@13966.4]
  assign StickySelects_12_io_ins_1 = io_rPort_2_en_0 & _T_1373; // @[MemPrimitives.scala 122:60:@13967.4]
  assign StickySelects_12_io_ins_2 = io_rPort_4_en_0 & _T_1379; // @[MemPrimitives.scala 122:60:@13968.4]
  assign StickySelects_12_io_ins_3 = io_rPort_5_en_0 & _T_1385; // @[MemPrimitives.scala 122:60:@13969.4]
  assign StickySelects_12_io_ins_4 = io_rPort_10_en_0 & _T_1391; // @[MemPrimitives.scala 122:60:@13970.4]
  assign StickySelects_12_io_ins_5 = io_rPort_11_en_0 & _T_1397; // @[MemPrimitives.scala 122:60:@13971.4]
  assign StickySelects_13_clock = clock; // @[:@14026.4]
  assign StickySelects_13_reset = reset; // @[:@14027.4]
  assign StickySelects_13_io_ins_0 = io_rPort_1_en_0 & _T_1429; // @[MemPrimitives.scala 122:60:@14028.4]
  assign StickySelects_13_io_ins_1 = io_rPort_3_en_0 & _T_1435; // @[MemPrimitives.scala 122:60:@14029.4]
  assign StickySelects_13_io_ins_2 = io_rPort_6_en_0 & _T_1441; // @[MemPrimitives.scala 122:60:@14030.4]
  assign StickySelects_13_io_ins_3 = io_rPort_7_en_0 & _T_1447; // @[MemPrimitives.scala 122:60:@14031.4]
  assign StickySelects_13_io_ins_4 = io_rPort_8_en_0 & _T_1453; // @[MemPrimitives.scala 122:60:@14032.4]
  assign StickySelects_13_io_ins_5 = io_rPort_9_en_0 & _T_1459; // @[MemPrimitives.scala 122:60:@14033.4]
  assign StickySelects_14_clock = clock; // @[:@14088.4]
  assign StickySelects_14_reset = reset; // @[:@14089.4]
  assign StickySelects_14_io_ins_0 = io_rPort_0_en_0 & _T_1491; // @[MemPrimitives.scala 122:60:@14090.4]
  assign StickySelects_14_io_ins_1 = io_rPort_2_en_0 & _T_1497; // @[MemPrimitives.scala 122:60:@14091.4]
  assign StickySelects_14_io_ins_2 = io_rPort_4_en_0 & _T_1503; // @[MemPrimitives.scala 122:60:@14092.4]
  assign StickySelects_14_io_ins_3 = io_rPort_5_en_0 & _T_1509; // @[MemPrimitives.scala 122:60:@14093.4]
  assign StickySelects_14_io_ins_4 = io_rPort_10_en_0 & _T_1515; // @[MemPrimitives.scala 122:60:@14094.4]
  assign StickySelects_14_io_ins_5 = io_rPort_11_en_0 & _T_1521; // @[MemPrimitives.scala 122:60:@14095.4]
  assign StickySelects_15_clock = clock; // @[:@14150.4]
  assign StickySelects_15_reset = reset; // @[:@14151.4]
  assign StickySelects_15_io_ins_0 = io_rPort_1_en_0 & _T_1553; // @[MemPrimitives.scala 122:60:@14152.4]
  assign StickySelects_15_io_ins_1 = io_rPort_3_en_0 & _T_1559; // @[MemPrimitives.scala 122:60:@14153.4]
  assign StickySelects_15_io_ins_2 = io_rPort_6_en_0 & _T_1565; // @[MemPrimitives.scala 122:60:@14154.4]
  assign StickySelects_15_io_ins_3 = io_rPort_7_en_0 & _T_1571; // @[MemPrimitives.scala 122:60:@14155.4]
  assign StickySelects_15_io_ins_4 = io_rPort_8_en_0 & _T_1577; // @[MemPrimitives.scala 122:60:@14156.4]
  assign StickySelects_15_io_ins_5 = io_rPort_9_en_0 & _T_1583; // @[MemPrimitives.scala 122:60:@14157.4]
  assign RetimeWrapper_clock = clock; // @[:@14213.4]
  assign RetimeWrapper_reset = reset; // @[:@14214.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14216.4]
  assign RetimeWrapper_io_in = _T_623 & io_rPort_0_en_0; // @[package.scala 94:16:@14215.4]
  assign RetimeWrapper_1_clock = clock; // @[:@14221.4]
  assign RetimeWrapper_1_reset = reset; // @[:@14222.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14224.4]
  assign RetimeWrapper_1_io_in = _T_747 & io_rPort_0_en_0; // @[package.scala 94:16:@14223.4]
  assign RetimeWrapper_2_clock = clock; // @[:@14229.4]
  assign RetimeWrapper_2_reset = reset; // @[:@14230.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14232.4]
  assign RetimeWrapper_2_io_in = _T_871 & io_rPort_0_en_0; // @[package.scala 94:16:@14231.4]
  assign RetimeWrapper_3_clock = clock; // @[:@14237.4]
  assign RetimeWrapper_3_reset = reset; // @[:@14238.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14240.4]
  assign RetimeWrapper_3_io_in = _T_995 & io_rPort_0_en_0; // @[package.scala 94:16:@14239.4]
  assign RetimeWrapper_4_clock = clock; // @[:@14245.4]
  assign RetimeWrapper_4_reset = reset; // @[:@14246.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14248.4]
  assign RetimeWrapper_4_io_in = _T_1119 & io_rPort_0_en_0; // @[package.scala 94:16:@14247.4]
  assign RetimeWrapper_5_clock = clock; // @[:@14253.4]
  assign RetimeWrapper_5_reset = reset; // @[:@14254.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14256.4]
  assign RetimeWrapper_5_io_in = _T_1243 & io_rPort_0_en_0; // @[package.scala 94:16:@14255.4]
  assign RetimeWrapper_6_clock = clock; // @[:@14261.4]
  assign RetimeWrapper_6_reset = reset; // @[:@14262.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14264.4]
  assign RetimeWrapper_6_io_in = _T_1367 & io_rPort_0_en_0; // @[package.scala 94:16:@14263.4]
  assign RetimeWrapper_7_clock = clock; // @[:@14269.4]
  assign RetimeWrapper_7_reset = reset; // @[:@14270.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14272.4]
  assign RetimeWrapper_7_io_in = _T_1491 & io_rPort_0_en_0; // @[package.scala 94:16:@14271.4]
  assign RetimeWrapper_8_clock = clock; // @[:@14309.4]
  assign RetimeWrapper_8_reset = reset; // @[:@14310.4]
  assign RetimeWrapper_8_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14312.4]
  assign RetimeWrapper_8_io_in = _T_685 & io_rPort_1_en_0; // @[package.scala 94:16:@14311.4]
  assign RetimeWrapper_9_clock = clock; // @[:@14317.4]
  assign RetimeWrapper_9_reset = reset; // @[:@14318.4]
  assign RetimeWrapper_9_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14320.4]
  assign RetimeWrapper_9_io_in = _T_809 & io_rPort_1_en_0; // @[package.scala 94:16:@14319.4]
  assign RetimeWrapper_10_clock = clock; // @[:@14325.4]
  assign RetimeWrapper_10_reset = reset; // @[:@14326.4]
  assign RetimeWrapper_10_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14328.4]
  assign RetimeWrapper_10_io_in = _T_933 & io_rPort_1_en_0; // @[package.scala 94:16:@14327.4]
  assign RetimeWrapper_11_clock = clock; // @[:@14333.4]
  assign RetimeWrapper_11_reset = reset; // @[:@14334.4]
  assign RetimeWrapper_11_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14336.4]
  assign RetimeWrapper_11_io_in = _T_1057 & io_rPort_1_en_0; // @[package.scala 94:16:@14335.4]
  assign RetimeWrapper_12_clock = clock; // @[:@14341.4]
  assign RetimeWrapper_12_reset = reset; // @[:@14342.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14344.4]
  assign RetimeWrapper_12_io_in = _T_1181 & io_rPort_1_en_0; // @[package.scala 94:16:@14343.4]
  assign RetimeWrapper_13_clock = clock; // @[:@14349.4]
  assign RetimeWrapper_13_reset = reset; // @[:@14350.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14352.4]
  assign RetimeWrapper_13_io_in = _T_1305 & io_rPort_1_en_0; // @[package.scala 94:16:@14351.4]
  assign RetimeWrapper_14_clock = clock; // @[:@14357.4]
  assign RetimeWrapper_14_reset = reset; // @[:@14358.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14360.4]
  assign RetimeWrapper_14_io_in = _T_1429 & io_rPort_1_en_0; // @[package.scala 94:16:@14359.4]
  assign RetimeWrapper_15_clock = clock; // @[:@14365.4]
  assign RetimeWrapper_15_reset = reset; // @[:@14366.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14368.4]
  assign RetimeWrapper_15_io_in = _T_1553 & io_rPort_1_en_0; // @[package.scala 94:16:@14367.4]
  assign RetimeWrapper_16_clock = clock; // @[:@14405.4]
  assign RetimeWrapper_16_reset = reset; // @[:@14406.4]
  assign RetimeWrapper_16_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14408.4]
  assign RetimeWrapper_16_io_in = _T_629 & io_rPort_2_en_0; // @[package.scala 94:16:@14407.4]
  assign RetimeWrapper_17_clock = clock; // @[:@14413.4]
  assign RetimeWrapper_17_reset = reset; // @[:@14414.4]
  assign RetimeWrapper_17_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14416.4]
  assign RetimeWrapper_17_io_in = _T_753 & io_rPort_2_en_0; // @[package.scala 94:16:@14415.4]
  assign RetimeWrapper_18_clock = clock; // @[:@14421.4]
  assign RetimeWrapper_18_reset = reset; // @[:@14422.4]
  assign RetimeWrapper_18_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14424.4]
  assign RetimeWrapper_18_io_in = _T_877 & io_rPort_2_en_0; // @[package.scala 94:16:@14423.4]
  assign RetimeWrapper_19_clock = clock; // @[:@14429.4]
  assign RetimeWrapper_19_reset = reset; // @[:@14430.4]
  assign RetimeWrapper_19_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14432.4]
  assign RetimeWrapper_19_io_in = _T_1001 & io_rPort_2_en_0; // @[package.scala 94:16:@14431.4]
  assign RetimeWrapper_20_clock = clock; // @[:@14437.4]
  assign RetimeWrapper_20_reset = reset; // @[:@14438.4]
  assign RetimeWrapper_20_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14440.4]
  assign RetimeWrapper_20_io_in = _T_1125 & io_rPort_2_en_0; // @[package.scala 94:16:@14439.4]
  assign RetimeWrapper_21_clock = clock; // @[:@14445.4]
  assign RetimeWrapper_21_reset = reset; // @[:@14446.4]
  assign RetimeWrapper_21_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14448.4]
  assign RetimeWrapper_21_io_in = _T_1249 & io_rPort_2_en_0; // @[package.scala 94:16:@14447.4]
  assign RetimeWrapper_22_clock = clock; // @[:@14453.4]
  assign RetimeWrapper_22_reset = reset; // @[:@14454.4]
  assign RetimeWrapper_22_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14456.4]
  assign RetimeWrapper_22_io_in = _T_1373 & io_rPort_2_en_0; // @[package.scala 94:16:@14455.4]
  assign RetimeWrapper_23_clock = clock; // @[:@14461.4]
  assign RetimeWrapper_23_reset = reset; // @[:@14462.4]
  assign RetimeWrapper_23_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14464.4]
  assign RetimeWrapper_23_io_in = _T_1497 & io_rPort_2_en_0; // @[package.scala 94:16:@14463.4]
  assign RetimeWrapper_24_clock = clock; // @[:@14501.4]
  assign RetimeWrapper_24_reset = reset; // @[:@14502.4]
  assign RetimeWrapper_24_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14504.4]
  assign RetimeWrapper_24_io_in = _T_691 & io_rPort_3_en_0; // @[package.scala 94:16:@14503.4]
  assign RetimeWrapper_25_clock = clock; // @[:@14509.4]
  assign RetimeWrapper_25_reset = reset; // @[:@14510.4]
  assign RetimeWrapper_25_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14512.4]
  assign RetimeWrapper_25_io_in = _T_815 & io_rPort_3_en_0; // @[package.scala 94:16:@14511.4]
  assign RetimeWrapper_26_clock = clock; // @[:@14517.4]
  assign RetimeWrapper_26_reset = reset; // @[:@14518.4]
  assign RetimeWrapper_26_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14520.4]
  assign RetimeWrapper_26_io_in = _T_939 & io_rPort_3_en_0; // @[package.scala 94:16:@14519.4]
  assign RetimeWrapper_27_clock = clock; // @[:@14525.4]
  assign RetimeWrapper_27_reset = reset; // @[:@14526.4]
  assign RetimeWrapper_27_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14528.4]
  assign RetimeWrapper_27_io_in = _T_1063 & io_rPort_3_en_0; // @[package.scala 94:16:@14527.4]
  assign RetimeWrapper_28_clock = clock; // @[:@14533.4]
  assign RetimeWrapper_28_reset = reset; // @[:@14534.4]
  assign RetimeWrapper_28_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14536.4]
  assign RetimeWrapper_28_io_in = _T_1187 & io_rPort_3_en_0; // @[package.scala 94:16:@14535.4]
  assign RetimeWrapper_29_clock = clock; // @[:@14541.4]
  assign RetimeWrapper_29_reset = reset; // @[:@14542.4]
  assign RetimeWrapper_29_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14544.4]
  assign RetimeWrapper_29_io_in = _T_1311 & io_rPort_3_en_0; // @[package.scala 94:16:@14543.4]
  assign RetimeWrapper_30_clock = clock; // @[:@14549.4]
  assign RetimeWrapper_30_reset = reset; // @[:@14550.4]
  assign RetimeWrapper_30_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14552.4]
  assign RetimeWrapper_30_io_in = _T_1435 & io_rPort_3_en_0; // @[package.scala 94:16:@14551.4]
  assign RetimeWrapper_31_clock = clock; // @[:@14557.4]
  assign RetimeWrapper_31_reset = reset; // @[:@14558.4]
  assign RetimeWrapper_31_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14560.4]
  assign RetimeWrapper_31_io_in = _T_1559 & io_rPort_3_en_0; // @[package.scala 94:16:@14559.4]
  assign RetimeWrapper_32_clock = clock; // @[:@14597.4]
  assign RetimeWrapper_32_reset = reset; // @[:@14598.4]
  assign RetimeWrapper_32_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14600.4]
  assign RetimeWrapper_32_io_in = _T_635 & io_rPort_4_en_0; // @[package.scala 94:16:@14599.4]
  assign RetimeWrapper_33_clock = clock; // @[:@14605.4]
  assign RetimeWrapper_33_reset = reset; // @[:@14606.4]
  assign RetimeWrapper_33_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14608.4]
  assign RetimeWrapper_33_io_in = _T_759 & io_rPort_4_en_0; // @[package.scala 94:16:@14607.4]
  assign RetimeWrapper_34_clock = clock; // @[:@14613.4]
  assign RetimeWrapper_34_reset = reset; // @[:@14614.4]
  assign RetimeWrapper_34_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14616.4]
  assign RetimeWrapper_34_io_in = _T_883 & io_rPort_4_en_0; // @[package.scala 94:16:@14615.4]
  assign RetimeWrapper_35_clock = clock; // @[:@14621.4]
  assign RetimeWrapper_35_reset = reset; // @[:@14622.4]
  assign RetimeWrapper_35_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14624.4]
  assign RetimeWrapper_35_io_in = _T_1007 & io_rPort_4_en_0; // @[package.scala 94:16:@14623.4]
  assign RetimeWrapper_36_clock = clock; // @[:@14629.4]
  assign RetimeWrapper_36_reset = reset; // @[:@14630.4]
  assign RetimeWrapper_36_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14632.4]
  assign RetimeWrapper_36_io_in = _T_1131 & io_rPort_4_en_0; // @[package.scala 94:16:@14631.4]
  assign RetimeWrapper_37_clock = clock; // @[:@14637.4]
  assign RetimeWrapper_37_reset = reset; // @[:@14638.4]
  assign RetimeWrapper_37_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14640.4]
  assign RetimeWrapper_37_io_in = _T_1255 & io_rPort_4_en_0; // @[package.scala 94:16:@14639.4]
  assign RetimeWrapper_38_clock = clock; // @[:@14645.4]
  assign RetimeWrapper_38_reset = reset; // @[:@14646.4]
  assign RetimeWrapper_38_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14648.4]
  assign RetimeWrapper_38_io_in = _T_1379 & io_rPort_4_en_0; // @[package.scala 94:16:@14647.4]
  assign RetimeWrapper_39_clock = clock; // @[:@14653.4]
  assign RetimeWrapper_39_reset = reset; // @[:@14654.4]
  assign RetimeWrapper_39_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14656.4]
  assign RetimeWrapper_39_io_in = _T_1503 & io_rPort_4_en_0; // @[package.scala 94:16:@14655.4]
  assign RetimeWrapper_40_clock = clock; // @[:@14693.4]
  assign RetimeWrapper_40_reset = reset; // @[:@14694.4]
  assign RetimeWrapper_40_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14696.4]
  assign RetimeWrapper_40_io_in = _T_641 & io_rPort_5_en_0; // @[package.scala 94:16:@14695.4]
  assign RetimeWrapper_41_clock = clock; // @[:@14701.4]
  assign RetimeWrapper_41_reset = reset; // @[:@14702.4]
  assign RetimeWrapper_41_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14704.4]
  assign RetimeWrapper_41_io_in = _T_765 & io_rPort_5_en_0; // @[package.scala 94:16:@14703.4]
  assign RetimeWrapper_42_clock = clock; // @[:@14709.4]
  assign RetimeWrapper_42_reset = reset; // @[:@14710.4]
  assign RetimeWrapper_42_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14712.4]
  assign RetimeWrapper_42_io_in = _T_889 & io_rPort_5_en_0; // @[package.scala 94:16:@14711.4]
  assign RetimeWrapper_43_clock = clock; // @[:@14717.4]
  assign RetimeWrapper_43_reset = reset; // @[:@14718.4]
  assign RetimeWrapper_43_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14720.4]
  assign RetimeWrapper_43_io_in = _T_1013 & io_rPort_5_en_0; // @[package.scala 94:16:@14719.4]
  assign RetimeWrapper_44_clock = clock; // @[:@14725.4]
  assign RetimeWrapper_44_reset = reset; // @[:@14726.4]
  assign RetimeWrapper_44_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14728.4]
  assign RetimeWrapper_44_io_in = _T_1137 & io_rPort_5_en_0; // @[package.scala 94:16:@14727.4]
  assign RetimeWrapper_45_clock = clock; // @[:@14733.4]
  assign RetimeWrapper_45_reset = reset; // @[:@14734.4]
  assign RetimeWrapper_45_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14736.4]
  assign RetimeWrapper_45_io_in = _T_1261 & io_rPort_5_en_0; // @[package.scala 94:16:@14735.4]
  assign RetimeWrapper_46_clock = clock; // @[:@14741.4]
  assign RetimeWrapper_46_reset = reset; // @[:@14742.4]
  assign RetimeWrapper_46_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14744.4]
  assign RetimeWrapper_46_io_in = _T_1385 & io_rPort_5_en_0; // @[package.scala 94:16:@14743.4]
  assign RetimeWrapper_47_clock = clock; // @[:@14749.4]
  assign RetimeWrapper_47_reset = reset; // @[:@14750.4]
  assign RetimeWrapper_47_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14752.4]
  assign RetimeWrapper_47_io_in = _T_1509 & io_rPort_5_en_0; // @[package.scala 94:16:@14751.4]
  assign RetimeWrapper_48_clock = clock; // @[:@14789.4]
  assign RetimeWrapper_48_reset = reset; // @[:@14790.4]
  assign RetimeWrapper_48_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14792.4]
  assign RetimeWrapper_48_io_in = _T_697 & io_rPort_6_en_0; // @[package.scala 94:16:@14791.4]
  assign RetimeWrapper_49_clock = clock; // @[:@14797.4]
  assign RetimeWrapper_49_reset = reset; // @[:@14798.4]
  assign RetimeWrapper_49_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14800.4]
  assign RetimeWrapper_49_io_in = _T_821 & io_rPort_6_en_0; // @[package.scala 94:16:@14799.4]
  assign RetimeWrapper_50_clock = clock; // @[:@14805.4]
  assign RetimeWrapper_50_reset = reset; // @[:@14806.4]
  assign RetimeWrapper_50_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14808.4]
  assign RetimeWrapper_50_io_in = _T_945 & io_rPort_6_en_0; // @[package.scala 94:16:@14807.4]
  assign RetimeWrapper_51_clock = clock; // @[:@14813.4]
  assign RetimeWrapper_51_reset = reset; // @[:@14814.4]
  assign RetimeWrapper_51_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14816.4]
  assign RetimeWrapper_51_io_in = _T_1069 & io_rPort_6_en_0; // @[package.scala 94:16:@14815.4]
  assign RetimeWrapper_52_clock = clock; // @[:@14821.4]
  assign RetimeWrapper_52_reset = reset; // @[:@14822.4]
  assign RetimeWrapper_52_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14824.4]
  assign RetimeWrapper_52_io_in = _T_1193 & io_rPort_6_en_0; // @[package.scala 94:16:@14823.4]
  assign RetimeWrapper_53_clock = clock; // @[:@14829.4]
  assign RetimeWrapper_53_reset = reset; // @[:@14830.4]
  assign RetimeWrapper_53_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14832.4]
  assign RetimeWrapper_53_io_in = _T_1317 & io_rPort_6_en_0; // @[package.scala 94:16:@14831.4]
  assign RetimeWrapper_54_clock = clock; // @[:@14837.4]
  assign RetimeWrapper_54_reset = reset; // @[:@14838.4]
  assign RetimeWrapper_54_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14840.4]
  assign RetimeWrapper_54_io_in = _T_1441 & io_rPort_6_en_0; // @[package.scala 94:16:@14839.4]
  assign RetimeWrapper_55_clock = clock; // @[:@14845.4]
  assign RetimeWrapper_55_reset = reset; // @[:@14846.4]
  assign RetimeWrapper_55_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14848.4]
  assign RetimeWrapper_55_io_in = _T_1565 & io_rPort_6_en_0; // @[package.scala 94:16:@14847.4]
  assign RetimeWrapper_56_clock = clock; // @[:@14885.4]
  assign RetimeWrapper_56_reset = reset; // @[:@14886.4]
  assign RetimeWrapper_56_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14888.4]
  assign RetimeWrapper_56_io_in = _T_703 & io_rPort_7_en_0; // @[package.scala 94:16:@14887.4]
  assign RetimeWrapper_57_clock = clock; // @[:@14893.4]
  assign RetimeWrapper_57_reset = reset; // @[:@14894.4]
  assign RetimeWrapper_57_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14896.4]
  assign RetimeWrapper_57_io_in = _T_827 & io_rPort_7_en_0; // @[package.scala 94:16:@14895.4]
  assign RetimeWrapper_58_clock = clock; // @[:@14901.4]
  assign RetimeWrapper_58_reset = reset; // @[:@14902.4]
  assign RetimeWrapper_58_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14904.4]
  assign RetimeWrapper_58_io_in = _T_951 & io_rPort_7_en_0; // @[package.scala 94:16:@14903.4]
  assign RetimeWrapper_59_clock = clock; // @[:@14909.4]
  assign RetimeWrapper_59_reset = reset; // @[:@14910.4]
  assign RetimeWrapper_59_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14912.4]
  assign RetimeWrapper_59_io_in = _T_1075 & io_rPort_7_en_0; // @[package.scala 94:16:@14911.4]
  assign RetimeWrapper_60_clock = clock; // @[:@14917.4]
  assign RetimeWrapper_60_reset = reset; // @[:@14918.4]
  assign RetimeWrapper_60_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14920.4]
  assign RetimeWrapper_60_io_in = _T_1199 & io_rPort_7_en_0; // @[package.scala 94:16:@14919.4]
  assign RetimeWrapper_61_clock = clock; // @[:@14925.4]
  assign RetimeWrapper_61_reset = reset; // @[:@14926.4]
  assign RetimeWrapper_61_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14928.4]
  assign RetimeWrapper_61_io_in = _T_1323 & io_rPort_7_en_0; // @[package.scala 94:16:@14927.4]
  assign RetimeWrapper_62_clock = clock; // @[:@14933.4]
  assign RetimeWrapper_62_reset = reset; // @[:@14934.4]
  assign RetimeWrapper_62_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14936.4]
  assign RetimeWrapper_62_io_in = _T_1447 & io_rPort_7_en_0; // @[package.scala 94:16:@14935.4]
  assign RetimeWrapper_63_clock = clock; // @[:@14941.4]
  assign RetimeWrapper_63_reset = reset; // @[:@14942.4]
  assign RetimeWrapper_63_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14944.4]
  assign RetimeWrapper_63_io_in = _T_1571 & io_rPort_7_en_0; // @[package.scala 94:16:@14943.4]
  assign RetimeWrapper_64_clock = clock; // @[:@14981.4]
  assign RetimeWrapper_64_reset = reset; // @[:@14982.4]
  assign RetimeWrapper_64_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14984.4]
  assign RetimeWrapper_64_io_in = _T_709 & io_rPort_8_en_0; // @[package.scala 94:16:@14983.4]
  assign RetimeWrapper_65_clock = clock; // @[:@14989.4]
  assign RetimeWrapper_65_reset = reset; // @[:@14990.4]
  assign RetimeWrapper_65_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14992.4]
  assign RetimeWrapper_65_io_in = _T_833 & io_rPort_8_en_0; // @[package.scala 94:16:@14991.4]
  assign RetimeWrapper_66_clock = clock; // @[:@14997.4]
  assign RetimeWrapper_66_reset = reset; // @[:@14998.4]
  assign RetimeWrapper_66_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15000.4]
  assign RetimeWrapper_66_io_in = _T_957 & io_rPort_8_en_0; // @[package.scala 94:16:@14999.4]
  assign RetimeWrapper_67_clock = clock; // @[:@15005.4]
  assign RetimeWrapper_67_reset = reset; // @[:@15006.4]
  assign RetimeWrapper_67_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15008.4]
  assign RetimeWrapper_67_io_in = _T_1081 & io_rPort_8_en_0; // @[package.scala 94:16:@15007.4]
  assign RetimeWrapper_68_clock = clock; // @[:@15013.4]
  assign RetimeWrapper_68_reset = reset; // @[:@15014.4]
  assign RetimeWrapper_68_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15016.4]
  assign RetimeWrapper_68_io_in = _T_1205 & io_rPort_8_en_0; // @[package.scala 94:16:@15015.4]
  assign RetimeWrapper_69_clock = clock; // @[:@15021.4]
  assign RetimeWrapper_69_reset = reset; // @[:@15022.4]
  assign RetimeWrapper_69_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15024.4]
  assign RetimeWrapper_69_io_in = _T_1329 & io_rPort_8_en_0; // @[package.scala 94:16:@15023.4]
  assign RetimeWrapper_70_clock = clock; // @[:@15029.4]
  assign RetimeWrapper_70_reset = reset; // @[:@15030.4]
  assign RetimeWrapper_70_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15032.4]
  assign RetimeWrapper_70_io_in = _T_1453 & io_rPort_8_en_0; // @[package.scala 94:16:@15031.4]
  assign RetimeWrapper_71_clock = clock; // @[:@15037.4]
  assign RetimeWrapper_71_reset = reset; // @[:@15038.4]
  assign RetimeWrapper_71_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15040.4]
  assign RetimeWrapper_71_io_in = _T_1577 & io_rPort_8_en_0; // @[package.scala 94:16:@15039.4]
  assign RetimeWrapper_72_clock = clock; // @[:@15077.4]
  assign RetimeWrapper_72_reset = reset; // @[:@15078.4]
  assign RetimeWrapper_72_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15080.4]
  assign RetimeWrapper_72_io_in = _T_715 & io_rPort_9_en_0; // @[package.scala 94:16:@15079.4]
  assign RetimeWrapper_73_clock = clock; // @[:@15085.4]
  assign RetimeWrapper_73_reset = reset; // @[:@15086.4]
  assign RetimeWrapper_73_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15088.4]
  assign RetimeWrapper_73_io_in = _T_839 & io_rPort_9_en_0; // @[package.scala 94:16:@15087.4]
  assign RetimeWrapper_74_clock = clock; // @[:@15093.4]
  assign RetimeWrapper_74_reset = reset; // @[:@15094.4]
  assign RetimeWrapper_74_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15096.4]
  assign RetimeWrapper_74_io_in = _T_963 & io_rPort_9_en_0; // @[package.scala 94:16:@15095.4]
  assign RetimeWrapper_75_clock = clock; // @[:@15101.4]
  assign RetimeWrapper_75_reset = reset; // @[:@15102.4]
  assign RetimeWrapper_75_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15104.4]
  assign RetimeWrapper_75_io_in = _T_1087 & io_rPort_9_en_0; // @[package.scala 94:16:@15103.4]
  assign RetimeWrapper_76_clock = clock; // @[:@15109.4]
  assign RetimeWrapper_76_reset = reset; // @[:@15110.4]
  assign RetimeWrapper_76_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15112.4]
  assign RetimeWrapper_76_io_in = _T_1211 & io_rPort_9_en_0; // @[package.scala 94:16:@15111.4]
  assign RetimeWrapper_77_clock = clock; // @[:@15117.4]
  assign RetimeWrapper_77_reset = reset; // @[:@15118.4]
  assign RetimeWrapper_77_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15120.4]
  assign RetimeWrapper_77_io_in = _T_1335 & io_rPort_9_en_0; // @[package.scala 94:16:@15119.4]
  assign RetimeWrapper_78_clock = clock; // @[:@15125.4]
  assign RetimeWrapper_78_reset = reset; // @[:@15126.4]
  assign RetimeWrapper_78_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15128.4]
  assign RetimeWrapper_78_io_in = _T_1459 & io_rPort_9_en_0; // @[package.scala 94:16:@15127.4]
  assign RetimeWrapper_79_clock = clock; // @[:@15133.4]
  assign RetimeWrapper_79_reset = reset; // @[:@15134.4]
  assign RetimeWrapper_79_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15136.4]
  assign RetimeWrapper_79_io_in = _T_1583 & io_rPort_9_en_0; // @[package.scala 94:16:@15135.4]
  assign RetimeWrapper_80_clock = clock; // @[:@15173.4]
  assign RetimeWrapper_80_reset = reset; // @[:@15174.4]
  assign RetimeWrapper_80_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15176.4]
  assign RetimeWrapper_80_io_in = _T_647 & io_rPort_10_en_0; // @[package.scala 94:16:@15175.4]
  assign RetimeWrapper_81_clock = clock; // @[:@15181.4]
  assign RetimeWrapper_81_reset = reset; // @[:@15182.4]
  assign RetimeWrapper_81_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15184.4]
  assign RetimeWrapper_81_io_in = _T_771 & io_rPort_10_en_0; // @[package.scala 94:16:@15183.4]
  assign RetimeWrapper_82_clock = clock; // @[:@15189.4]
  assign RetimeWrapper_82_reset = reset; // @[:@15190.4]
  assign RetimeWrapper_82_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15192.4]
  assign RetimeWrapper_82_io_in = _T_895 & io_rPort_10_en_0; // @[package.scala 94:16:@15191.4]
  assign RetimeWrapper_83_clock = clock; // @[:@15197.4]
  assign RetimeWrapper_83_reset = reset; // @[:@15198.4]
  assign RetimeWrapper_83_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15200.4]
  assign RetimeWrapper_83_io_in = _T_1019 & io_rPort_10_en_0; // @[package.scala 94:16:@15199.4]
  assign RetimeWrapper_84_clock = clock; // @[:@15205.4]
  assign RetimeWrapper_84_reset = reset; // @[:@15206.4]
  assign RetimeWrapper_84_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15208.4]
  assign RetimeWrapper_84_io_in = _T_1143 & io_rPort_10_en_0; // @[package.scala 94:16:@15207.4]
  assign RetimeWrapper_85_clock = clock; // @[:@15213.4]
  assign RetimeWrapper_85_reset = reset; // @[:@15214.4]
  assign RetimeWrapper_85_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15216.4]
  assign RetimeWrapper_85_io_in = _T_1267 & io_rPort_10_en_0; // @[package.scala 94:16:@15215.4]
  assign RetimeWrapper_86_clock = clock; // @[:@15221.4]
  assign RetimeWrapper_86_reset = reset; // @[:@15222.4]
  assign RetimeWrapper_86_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15224.4]
  assign RetimeWrapper_86_io_in = _T_1391 & io_rPort_10_en_0; // @[package.scala 94:16:@15223.4]
  assign RetimeWrapper_87_clock = clock; // @[:@15229.4]
  assign RetimeWrapper_87_reset = reset; // @[:@15230.4]
  assign RetimeWrapper_87_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15232.4]
  assign RetimeWrapper_87_io_in = _T_1515 & io_rPort_10_en_0; // @[package.scala 94:16:@15231.4]
  assign RetimeWrapper_88_clock = clock; // @[:@15269.4]
  assign RetimeWrapper_88_reset = reset; // @[:@15270.4]
  assign RetimeWrapper_88_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15272.4]
  assign RetimeWrapper_88_io_in = _T_653 & io_rPort_11_en_0; // @[package.scala 94:16:@15271.4]
  assign RetimeWrapper_89_clock = clock; // @[:@15277.4]
  assign RetimeWrapper_89_reset = reset; // @[:@15278.4]
  assign RetimeWrapper_89_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15280.4]
  assign RetimeWrapper_89_io_in = _T_777 & io_rPort_11_en_0; // @[package.scala 94:16:@15279.4]
  assign RetimeWrapper_90_clock = clock; // @[:@15285.4]
  assign RetimeWrapper_90_reset = reset; // @[:@15286.4]
  assign RetimeWrapper_90_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15288.4]
  assign RetimeWrapper_90_io_in = _T_901 & io_rPort_11_en_0; // @[package.scala 94:16:@15287.4]
  assign RetimeWrapper_91_clock = clock; // @[:@15293.4]
  assign RetimeWrapper_91_reset = reset; // @[:@15294.4]
  assign RetimeWrapper_91_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15296.4]
  assign RetimeWrapper_91_io_in = _T_1025 & io_rPort_11_en_0; // @[package.scala 94:16:@15295.4]
  assign RetimeWrapper_92_clock = clock; // @[:@15301.4]
  assign RetimeWrapper_92_reset = reset; // @[:@15302.4]
  assign RetimeWrapper_92_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15304.4]
  assign RetimeWrapper_92_io_in = _T_1149 & io_rPort_11_en_0; // @[package.scala 94:16:@15303.4]
  assign RetimeWrapper_93_clock = clock; // @[:@15309.4]
  assign RetimeWrapper_93_reset = reset; // @[:@15310.4]
  assign RetimeWrapper_93_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15312.4]
  assign RetimeWrapper_93_io_in = _T_1273 & io_rPort_11_en_0; // @[package.scala 94:16:@15311.4]
  assign RetimeWrapper_94_clock = clock; // @[:@15317.4]
  assign RetimeWrapper_94_reset = reset; // @[:@15318.4]
  assign RetimeWrapper_94_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15320.4]
  assign RetimeWrapper_94_io_in = _T_1397 & io_rPort_11_en_0; // @[package.scala 94:16:@15319.4]
  assign RetimeWrapper_95_clock = clock; // @[:@15325.4]
  assign RetimeWrapper_95_reset = reset; // @[:@15326.4]
  assign RetimeWrapper_95_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15328.4]
  assign RetimeWrapper_95_io_in = _T_1521 & io_rPort_11_en_0; // @[package.scala 94:16:@15327.4]
endmodule
module RetimeWrapper_165( // @[:@15352.2]
  input         clock, // @[:@15353.4]
  input         reset, // @[:@15354.4]
  input         io_flow, // @[:@15355.4]
  input  [31:0] io_in, // @[:@15355.4]
  output [31:0] io_out // @[:@15355.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15357.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15357.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15357.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15357.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15357.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15357.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@15357.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15370.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15369.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15368.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15367.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15366.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15364.4]
endmodule
module RetimeWrapper_167( // @[:@15574.2]
  input         clock, // @[:@15575.4]
  input         reset, // @[:@15576.4]
  input         io_flow, // @[:@15577.4]
  input  [31:0] io_in, // @[:@15577.4]
  output [31:0] io_out // @[:@15577.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15579.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15579.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15579.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15579.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15579.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15579.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@15579.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15592.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15591.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15590.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15589.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15588.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15586.4]
endmodule
module RetimeWrapper_170( // @[:@15827.2]
  input        clock, // @[:@15828.4]
  input        reset, // @[:@15829.4]
  input        io_flow, // @[:@15830.4]
  input  [7:0] io_in, // @[:@15830.4]
  output [7:0] io_out // @[:@15830.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15832.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15832.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15832.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15832.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15832.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15832.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@15832.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15845.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15844.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@15843.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15842.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15841.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15839.4]
endmodule
module RetimeWrapper_174( // @[:@15955.2]
  input         clock, // @[:@15956.4]
  input         reset, // @[:@15957.4]
  input         io_flow, // @[:@15958.4]
  input  [31:0] io_in, // @[:@15958.4]
  output [31:0] io_out // @[:@15958.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15960.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15960.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15960.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15960.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15960.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15960.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@15960.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15973.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15972.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15971.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15970.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15969.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15967.4]
endmodule
module RetimeWrapper_180( // @[:@16461.2]
  input         clock, // @[:@16462.4]
  input         reset, // @[:@16463.4]
  input         io_flow, // @[:@16464.4]
  input  [31:0] io_in, // @[:@16464.4]
  output [31:0] io_out // @[:@16464.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16466.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16466.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16466.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16466.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16466.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16466.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@16466.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16479.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16478.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16477.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16476.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16475.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16473.4]
endmodule
module RetimeWrapper_183( // @[:@16557.2]
  input         clock, // @[:@16558.4]
  input         reset, // @[:@16559.4]
  input         io_flow, // @[:@16560.4]
  input  [31:0] io_in, // @[:@16560.4]
  output [31:0] io_out // @[:@16560.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16562.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16562.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16562.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16562.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16562.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16562.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@16562.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16575.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16574.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16573.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16572.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16571.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16569.4]
endmodule
module RetimeWrapper_187( // @[:@16685.2]
  input         clock, // @[:@16686.4]
  input         reset, // @[:@16687.4]
  input         io_flow, // @[:@16688.4]
  input  [40:0] io_in, // @[:@16688.4]
  output [40:0] io_out // @[:@16688.4]
);
  wire [40:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16690.4]
  wire [40:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16690.4]
  wire [40:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16690.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16690.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16690.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16690.4]
  RetimeShiftRegister #(.WIDTH(41), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@16690.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16703.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16702.4]
  assign sr_init = 41'h0; // @[RetimeShiftRegister.scala 19:16:@16701.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16700.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16699.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16697.4]
endmodule
module RetimeWrapper_188( // @[:@16717.2]
  input         clock, // @[:@16718.4]
  input         reset, // @[:@16719.4]
  input         io_flow, // @[:@16720.4]
  input  [36:0] io_in, // @[:@16720.4]
  output [36:0] io_out // @[:@16720.4]
);
  wire [36:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16722.4]
  wire [36:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16722.4]
  wire [36:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16722.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16722.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16722.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16722.4]
  RetimeShiftRegister #(.WIDTH(37), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@16722.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16735.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16734.4]
  assign sr_init = 37'h0; // @[RetimeShiftRegister.scala 19:16:@16733.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16732.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16731.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16729.4]
endmodule
module RetimeWrapper_190( // @[:@16939.2]
  input         clock, // @[:@16940.4]
  input         reset, // @[:@16941.4]
  input         io_flow, // @[:@16942.4]
  input  [31:0] io_in, // @[:@16942.4]
  output [31:0] io_out // @[:@16942.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16944.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16944.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16944.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16944.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16944.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16944.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(9)) sr ( // @[RetimeShiftRegister.scala 15:20:@16944.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16957.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16956.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16955.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16954.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16953.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16951.4]
endmodule
module RetimeWrapper_192( // @[:@17160.2]
  input         clock, // @[:@17161.4]
  input         reset, // @[:@17162.4]
  input         io_flow, // @[:@17163.4]
  input  [31:0] io_in, // @[:@17163.4]
  output [31:0] io_out // @[:@17163.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17165.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17165.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17165.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17165.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17165.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17165.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@17165.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17178.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17177.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17176.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17175.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17174.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17172.4]
endmodule
module RetimeWrapper_194( // @[:@17224.2]
  input   clock, // @[:@17225.4]
  input   reset, // @[:@17226.4]
  input   io_flow, // @[:@17227.4]
  input   io_in, // @[:@17227.4]
  output  io_out // @[:@17227.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@17229.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@17229.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@17229.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17229.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17229.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17229.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(14)) sr ( // @[RetimeShiftRegister.scala 15:20:@17229.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17242.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17241.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@17240.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17239.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17238.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17236.4]
endmodule
module RetimeWrapper_196( // @[:@17288.2]
  input         clock, // @[:@17289.4]
  input         reset, // @[:@17290.4]
  input         io_flow, // @[:@17291.4]
  input  [31:0] io_in, // @[:@17291.4]
  output [31:0] io_out // @[:@17291.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17293.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17293.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17293.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17293.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17293.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17293.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(13)) sr ( // @[RetimeShiftRegister.scala 15:20:@17293.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17306.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17305.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17304.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17303.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17302.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17300.4]
endmodule
module RetimeWrapper_201( // @[:@17448.2]
  input         clock, // @[:@17449.4]
  input         reset, // @[:@17450.4]
  input         io_flow, // @[:@17451.4]
  input  [31:0] io_in, // @[:@17451.4]
  output [31:0] io_out // @[:@17451.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17453.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17453.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17453.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17453.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17453.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17453.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(10)) sr ( // @[RetimeShiftRegister.scala 15:20:@17453.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17466.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17465.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17464.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17463.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17462.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17460.4]
endmodule
module RetimeWrapper_205( // @[:@17733.2]
  input         clock, // @[:@17734.4]
  input         reset, // @[:@17735.4]
  input         io_flow, // @[:@17736.4]
  input  [31:0] io_in, // @[:@17736.4]
  output [31:0] io_out // @[:@17736.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17738.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17738.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17738.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17738.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17738.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17738.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(14)) sr ( // @[RetimeShiftRegister.scala 15:20:@17738.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17751.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17750.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17749.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17748.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17747.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17745.4]
endmodule
module RetimeWrapper_236( // @[:@19826.2]
  input         clock, // @[:@19827.4]
  input         reset, // @[:@19828.4]
  input         io_flow, // @[:@19829.4]
  input  [31:0] io_in, // @[:@19829.4]
  output [31:0] io_out // @[:@19829.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@19831.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@19831.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@19831.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@19831.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@19831.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@19831.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(11)) sr ( // @[RetimeShiftRegister.scala 15:20:@19831.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@19844.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@19843.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@19842.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@19841.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@19840.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@19838.4]
endmodule
module SimBlackBoxesfix2fixBox_64( // @[:@22573.2]
  input  [7:0] io_a, // @[:@22576.4]
  output [8:0] io_b // @[:@22576.4]
);
  assign io_b = {1'h0,io_a}; // @[SimBlackBoxes.scala 99:40:@22590.4]
endmodule
module __62( // @[:@22592.2]
  input  [7:0] io_b, // @[:@22595.4]
  output [8:0] io_result // @[:@22595.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@22600.4]
  wire [8:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@22600.4]
  SimBlackBoxesfix2fixBox_64 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@22600.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@22613.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@22608.4]
endmodule
module fix2fixBox_29( // @[:@22657.2]
  input  [8:0] io_a, // @[:@22660.4]
  output [7:0] io_b // @[:@22660.4]
);
  assign io_b = io_a[7:0]; // @[Converter.scala 95:38:@22673.4]
endmodule
module x499_x15( // @[:@22675.2]
  input  [7:0] io_a, // @[:@22678.4]
  input  [7:0] io_b, // @[:@22678.4]
  output [7:0] io_result // @[:@22678.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@22686.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@22686.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@22693.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@22693.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@22703.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@22703.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@22691.4 Math.scala 713:14:@22692.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@22698.4 Math.scala 713:14:@22699.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@22700.4]
  __62 _ ( // @[Math.scala 709:24:@22686.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __62 __1 ( // @[Math.scala 709:24:@22693.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_29 fix2fixBox ( // @[Math.scala 141:30:@22703.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@22691.4 Math.scala 713:14:@22692.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@22698.4 Math.scala 713:14:@22699.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@22700.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@22711.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@22689.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@22696.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@22706.4]
endmodule
module RetimeWrapper_278( // @[:@23649.2]
  input        clock, // @[:@23650.4]
  input        reset, // @[:@23651.4]
  input        io_flow, // @[:@23652.4]
  input  [7:0] io_in, // @[:@23652.4]
  output [7:0] io_out // @[:@23652.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@23654.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@23654.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@23654.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@23654.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@23654.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@23654.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@23654.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@23667.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@23666.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@23665.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@23664.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@23663.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@23661.4]
endmodule
module fix2fixBox_36( // @[:@23669.2]
  input        clock, // @[:@23670.4]
  input        reset, // @[:@23671.4]
  input  [8:0] io_a, // @[:@23672.4]
  input        io_flow, // @[:@23672.4]
  output [7:0] io_b // @[:@23672.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@23685.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@23685.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@23685.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@23685.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@23685.4]
  RetimeWrapper_278 RetimeWrapper ( // @[package.scala 93:22:@23685.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@23692.4]
  assign RetimeWrapper_clock = clock; // @[:@23686.4]
  assign RetimeWrapper_reset = reset; // @[:@23687.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@23689.4]
  assign RetimeWrapper_io_in = io_a[7:0]; // @[package.scala 94:16:@23688.4]
endmodule
module x506_sum( // @[:@23694.2]
  input        clock, // @[:@23695.4]
  input        reset, // @[:@23696.4]
  input  [7:0] io_a, // @[:@23697.4]
  input  [7:0] io_b, // @[:@23697.4]
  input        io_flow, // @[:@23697.4]
  output [7:0] io_result // @[:@23697.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@23705.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@23705.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@23712.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@23712.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@23722.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@23722.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@23722.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@23722.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@23722.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@23710.4 Math.scala 713:14:@23711.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@23717.4 Math.scala 713:14:@23718.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@23719.4]
  __62 _ ( // @[Math.scala 709:24:@23705.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __62 __1 ( // @[Math.scala 709:24:@23712.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_36 fix2fixBox ( // @[Math.scala 141:30:@23722.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@23710.4 Math.scala 713:14:@23711.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@23717.4 Math.scala 713:14:@23718.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@23719.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@23730.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@23708.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@23715.4]
  assign fix2fixBox_clock = clock; // @[:@23723.4]
  assign fix2fixBox_reset = reset; // @[:@23724.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@23725.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@23728.4]
endmodule
module RetimeWrapper_280( // @[:@24903.2]
  input         clock, // @[:@24904.4]
  input         reset, // @[:@24905.4]
  input         io_flow, // @[:@24906.4]
  input  [15:0] io_in, // @[:@24906.4]
  output [15:0] io_out // @[:@24906.4]
);
  wire [15:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@24908.4]
  wire [15:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@24908.4]
  wire [15:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@24908.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@24908.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@24908.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@24908.4]
  RetimeShiftRegister #(.WIDTH(16), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@24908.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@24921.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@24920.4]
  assign sr_init = 16'h0; // @[RetimeShiftRegister.scala 19:16:@24919.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@24918.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@24917.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@24915.4]
endmodule
module x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@25019.2]
  input          clock, // @[:@25020.4]
  input          reset, // @[:@25021.4]
  output         io_in_x348_TREADY, // @[:@25022.4]
  input  [255:0] io_in_x348_TDATA, // @[:@25022.4]
  input  [7:0]   io_in_x348_TID, // @[:@25022.4]
  input  [7:0]   io_in_x348_TDEST, // @[:@25022.4]
  output         io_in_x349_TVALID, // @[:@25022.4]
  input          io_in_x349_TREADY, // @[:@25022.4]
  output [255:0] io_in_x349_TDATA, // @[:@25022.4]
  input          io_sigsIn_backpressure, // @[:@25022.4]
  input          io_sigsIn_datapathEn, // @[:@25022.4]
  input          io_sigsIn_break, // @[:@25022.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@25022.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@25022.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@25022.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@25022.4]
  input          io_rr // @[:@25022.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@25036.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@25036.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@25048.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@25048.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@25071.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@25071.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@25071.4]
  wire [15:0] RetimeWrapper_io_in; // @[package.scala 93:22:@25071.4]
  wire [15:0] RetimeWrapper_io_out; // @[package.scala 93:22:@25071.4]
  wire  x385_lb_0_clock; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_reset; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_11_banks_1; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_11_banks_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [8:0] x385_lb_0_io_rPort_11_ofs_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_11_en_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_11_backpressure; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [7:0] x385_lb_0_io_rPort_11_output_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_10_banks_1; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_10_banks_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [8:0] x385_lb_0_io_rPort_10_ofs_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_10_en_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_10_backpressure; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [7:0] x385_lb_0_io_rPort_10_output_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_9_banks_1; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_9_banks_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [8:0] x385_lb_0_io_rPort_9_ofs_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_9_en_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_9_backpressure; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [7:0] x385_lb_0_io_rPort_9_output_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_8_banks_1; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_8_banks_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [8:0] x385_lb_0_io_rPort_8_ofs_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_8_en_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_8_backpressure; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [7:0] x385_lb_0_io_rPort_8_output_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_7_banks_1; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_7_banks_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [8:0] x385_lb_0_io_rPort_7_ofs_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_7_en_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_7_backpressure; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [7:0] x385_lb_0_io_rPort_7_output_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_6_banks_1; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_6_banks_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [8:0] x385_lb_0_io_rPort_6_ofs_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_6_en_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_6_backpressure; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [7:0] x385_lb_0_io_rPort_6_output_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_5_banks_1; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_5_banks_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [8:0] x385_lb_0_io_rPort_5_ofs_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_5_en_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_5_backpressure; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [7:0] x385_lb_0_io_rPort_5_output_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_4_banks_1; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_4_banks_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [8:0] x385_lb_0_io_rPort_4_ofs_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_4_en_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_4_backpressure; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [7:0] x385_lb_0_io_rPort_4_output_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_3_banks_1; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_3_banks_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [8:0] x385_lb_0_io_rPort_3_ofs_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_3_en_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_3_backpressure; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [7:0] x385_lb_0_io_rPort_3_output_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_2_banks_1; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_2_banks_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [8:0] x385_lb_0_io_rPort_2_ofs_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_2_en_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_2_backpressure; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [7:0] x385_lb_0_io_rPort_2_output_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_1_banks_1; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_1_banks_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [8:0] x385_lb_0_io_rPort_1_ofs_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_1_en_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_1_backpressure; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [7:0] x385_lb_0_io_rPort_1_output_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_0_banks_1; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_rPort_0_banks_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [8:0] x385_lb_0_io_rPort_0_ofs_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_0_en_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_rPort_0_backpressure; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [7:0] x385_lb_0_io_rPort_0_output_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_wPort_1_banks_1; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_wPort_1_banks_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [8:0] x385_lb_0_io_wPort_1_ofs_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [7:0] x385_lb_0_io_wPort_1_data_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_wPort_1_en_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_wPort_0_banks_1; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [2:0] x385_lb_0_io_wPort_0_banks_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [8:0] x385_lb_0_io_wPort_0_ofs_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire [7:0] x385_lb_0_io_wPort_0_data_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  x385_lb_0_io_wPort_0_en_0; // @[m_x385_lb_0.scala 39:17:@25081.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@25231.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@25231.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@25231.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@25231.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@25231.4]
  wire  x588_sub_1_clock; // @[Math.scala 191:24:@25281.4]
  wire  x588_sub_1_reset; // @[Math.scala 191:24:@25281.4]
  wire [31:0] x588_sub_1_io_a; // @[Math.scala 191:24:@25281.4]
  wire [31:0] x588_sub_1_io_b; // @[Math.scala 191:24:@25281.4]
  wire  x588_sub_1_io_flow; // @[Math.scala 191:24:@25281.4]
  wire [31:0] x588_sub_1_io_result; // @[Math.scala 191:24:@25281.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@25300.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@25300.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@25300.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@25300.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@25300.4]
  wire  x398_sum_1_clock; // @[Math.scala 150:24:@25309.4]
  wire  x398_sum_1_reset; // @[Math.scala 150:24:@25309.4]
  wire [31:0] x398_sum_1_io_a; // @[Math.scala 150:24:@25309.4]
  wire [31:0] x398_sum_1_io_b; // @[Math.scala 150:24:@25309.4]
  wire  x398_sum_1_io_flow; // @[Math.scala 150:24:@25309.4]
  wire [31:0] x398_sum_1_io_result; // @[Math.scala 150:24:@25309.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@25319.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@25319.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@25319.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@25319.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@25319.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@25328.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@25328.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@25328.4]
  wire [7:0] RetimeWrapper_4_io_in; // @[package.scala 93:22:@25328.4]
  wire [7:0] RetimeWrapper_4_io_out; // @[package.scala 93:22:@25328.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@25337.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@25337.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@25337.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@25337.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@25337.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@25346.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@25346.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@25346.4]
  wire [31:0] RetimeWrapper_6_io_in; // @[package.scala 93:22:@25346.4]
  wire [31:0] RetimeWrapper_6_io_out; // @[package.scala 93:22:@25346.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@25355.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@25355.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@25355.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@25355.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@25355.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@25364.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@25364.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@25364.4]
  wire [31:0] RetimeWrapper_8_io_in; // @[package.scala 93:22:@25364.4]
  wire [31:0] RetimeWrapper_8_io_out; // @[package.scala 93:22:@25364.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@25375.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@25375.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@25375.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@25375.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@25375.4]
  wire  x400_rdcol_1_clock; // @[Math.scala 150:24:@25398.4]
  wire  x400_rdcol_1_reset; // @[Math.scala 150:24:@25398.4]
  wire [31:0] x400_rdcol_1_io_a; // @[Math.scala 150:24:@25398.4]
  wire [31:0] x400_rdcol_1_io_b; // @[Math.scala 150:24:@25398.4]
  wire  x400_rdcol_1_io_flow; // @[Math.scala 150:24:@25398.4]
  wire [31:0] x400_rdcol_1_io_result; // @[Math.scala 150:24:@25398.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@25430.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@25430.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@25430.4]
  wire [31:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@25430.4]
  wire [31:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@25430.4]
  wire  x404_sum_1_clock; // @[Math.scala 150:24:@25439.4]
  wire  x404_sum_1_reset; // @[Math.scala 150:24:@25439.4]
  wire [31:0] x404_sum_1_io_a; // @[Math.scala 150:24:@25439.4]
  wire [31:0] x404_sum_1_io_b; // @[Math.scala 150:24:@25439.4]
  wire  x404_sum_1_io_flow; // @[Math.scala 150:24:@25439.4]
  wire [31:0] x404_sum_1_io_result; // @[Math.scala 150:24:@25439.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@25449.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@25449.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@25449.4]
  wire [31:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@25449.4]
  wire [31:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@25449.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@25458.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@25458.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@25458.4]
  wire [31:0] RetimeWrapper_12_io_in; // @[package.scala 93:22:@25458.4]
  wire [31:0] RetimeWrapper_12_io_out; // @[package.scala 93:22:@25458.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@25467.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@25467.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@25467.4]
  wire [7:0] RetimeWrapper_13_io_in; // @[package.scala 93:22:@25467.4]
  wire [7:0] RetimeWrapper_13_io_out; // @[package.scala 93:22:@25467.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@25478.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@25478.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@25478.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@25478.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@25478.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@25499.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@25499.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@25499.4]
  wire [31:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@25499.4]
  wire [31:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@25499.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@25526.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@25526.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@25526.4]
  wire [31:0] RetimeWrapper_16_io_in; // @[package.scala 93:22:@25526.4]
  wire [31:0] RetimeWrapper_16_io_out; // @[package.scala 93:22:@25526.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@25542.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@25542.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@25542.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@25542.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@25542.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@25554.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@25554.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@25554.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@25554.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@25554.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@25590.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@25590.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@25590.4]
  wire [40:0] RetimeWrapper_19_io_in; // @[package.scala 93:22:@25590.4]
  wire [40:0] RetimeWrapper_19_io_out; // @[package.scala 93:22:@25590.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@25602.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@25602.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@25602.4]
  wire [36:0] RetimeWrapper_20_io_in; // @[package.scala 93:22:@25602.4]
  wire [36:0] RetimeWrapper_20_io_out; // @[package.scala 93:22:@25602.4]
  wire  x594_sub_1_clock; // @[Math.scala 191:24:@25612.4]
  wire  x594_sub_1_reset; // @[Math.scala 191:24:@25612.4]
  wire [31:0] x594_sub_1_io_a; // @[Math.scala 191:24:@25612.4]
  wire [31:0] x594_sub_1_io_b; // @[Math.scala 191:24:@25612.4]
  wire  x594_sub_1_io_flow; // @[Math.scala 191:24:@25612.4]
  wire [31:0] x594_sub_1_io_result; // @[Math.scala 191:24:@25612.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@25622.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@25622.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@25622.4]
  wire [31:0] RetimeWrapper_21_io_in; // @[package.scala 93:22:@25622.4]
  wire [31:0] RetimeWrapper_21_io_out; // @[package.scala 93:22:@25622.4]
  wire  x415_sum_1_clock; // @[Math.scala 150:24:@25631.4]
  wire  x415_sum_1_reset; // @[Math.scala 150:24:@25631.4]
  wire [31:0] x415_sum_1_io_a; // @[Math.scala 150:24:@25631.4]
  wire [31:0] x415_sum_1_io_b; // @[Math.scala 150:24:@25631.4]
  wire  x415_sum_1_io_flow; // @[Math.scala 150:24:@25631.4]
  wire [31:0] x415_sum_1_io_result; // @[Math.scala 150:24:@25631.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@25641.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@25641.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@25641.4]
  wire [31:0] RetimeWrapper_22_io_in; // @[package.scala 93:22:@25641.4]
  wire [31:0] RetimeWrapper_22_io_out; // @[package.scala 93:22:@25641.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@25650.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@25650.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@25650.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@25650.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@25650.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@25659.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@25659.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@25659.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@25659.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@25659.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@25668.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@25668.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@25668.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@25668.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@25668.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@25677.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@25677.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@25677.4]
  wire [31:0] RetimeWrapper_26_io_in; // @[package.scala 93:22:@25677.4]
  wire [31:0] RetimeWrapper_26_io_out; // @[package.scala 93:22:@25677.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@25686.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@25686.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@25686.4]
  wire [31:0] RetimeWrapper_27_io_in; // @[package.scala 93:22:@25686.4]
  wire [31:0] RetimeWrapper_27_io_out; // @[package.scala 93:22:@25686.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@25698.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@25698.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@25698.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@25698.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@25698.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@25719.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@25719.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@25719.4]
  wire [31:0] RetimeWrapper_29_io_in; // @[package.scala 93:22:@25719.4]
  wire [31:0] RetimeWrapper_29_io_out; // @[package.scala 93:22:@25719.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@25738.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@25738.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@25738.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@25738.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@25738.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@25750.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@25750.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@25750.4]
  wire [31:0] RetimeWrapper_31_io_in; // @[package.scala 93:22:@25750.4]
  wire [31:0] RetimeWrapper_31_io_out; // @[package.scala 93:22:@25750.4]
  wire  x421_sum_1_clock; // @[Math.scala 150:24:@25759.4]
  wire  x421_sum_1_reset; // @[Math.scala 150:24:@25759.4]
  wire [31:0] x421_sum_1_io_a; // @[Math.scala 150:24:@25759.4]
  wire [31:0] x421_sum_1_io_b; // @[Math.scala 150:24:@25759.4]
  wire  x421_sum_1_io_flow; // @[Math.scala 150:24:@25759.4]
  wire [31:0] x421_sum_1_io_result; // @[Math.scala 150:24:@25759.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@25769.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@25769.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@25769.4]
  wire [31:0] RetimeWrapper_32_io_in; // @[package.scala 93:22:@25769.4]
  wire [31:0] RetimeWrapper_32_io_out; // @[package.scala 93:22:@25769.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@25778.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@25778.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@25778.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@25778.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@25778.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@25787.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@25787.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@25787.4]
  wire [31:0] RetimeWrapper_34_io_in; // @[package.scala 93:22:@25787.4]
  wire [31:0] RetimeWrapper_34_io_out; // @[package.scala 93:22:@25787.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@25799.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@25799.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@25799.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@25799.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@25799.4]
  wire  x424_rdcol_1_clock; // @[Math.scala 150:24:@25822.4]
  wire  x424_rdcol_1_reset; // @[Math.scala 150:24:@25822.4]
  wire [31:0] x424_rdcol_1_io_a; // @[Math.scala 150:24:@25822.4]
  wire [31:0] x424_rdcol_1_io_b; // @[Math.scala 150:24:@25822.4]
  wire  x424_rdcol_1_io_flow; // @[Math.scala 150:24:@25822.4]
  wire [31:0] x424_rdcol_1_io_result; // @[Math.scala 150:24:@25822.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@25842.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@25842.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@25842.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@25842.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@25842.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@25874.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@25874.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@25874.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@25874.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@25874.4]
  wire  x430_sum_1_clock; // @[Math.scala 150:24:@25883.4]
  wire  x430_sum_1_reset; // @[Math.scala 150:24:@25883.4]
  wire [31:0] x430_sum_1_io_a; // @[Math.scala 150:24:@25883.4]
  wire [31:0] x430_sum_1_io_b; // @[Math.scala 150:24:@25883.4]
  wire  x430_sum_1_io_flow; // @[Math.scala 150:24:@25883.4]
  wire [31:0] x430_sum_1_io_result; // @[Math.scala 150:24:@25883.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@25893.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@25893.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@25893.4]
  wire [31:0] RetimeWrapper_38_io_in; // @[package.scala 93:22:@25893.4]
  wire [31:0] RetimeWrapper_38_io_out; // @[package.scala 93:22:@25893.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@25902.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@25902.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@25902.4]
  wire [31:0] RetimeWrapper_39_io_in; // @[package.scala 93:22:@25902.4]
  wire [31:0] RetimeWrapper_39_io_out; // @[package.scala 93:22:@25902.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@25911.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@25911.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@25911.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@25911.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@25911.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@25923.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@25923.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@25923.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@25923.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@25923.4]
  wire  x433_rdcol_1_clock; // @[Math.scala 150:24:@25946.4]
  wire  x433_rdcol_1_reset; // @[Math.scala 150:24:@25946.4]
  wire [31:0] x433_rdcol_1_io_a; // @[Math.scala 150:24:@25946.4]
  wire [31:0] x433_rdcol_1_io_b; // @[Math.scala 150:24:@25946.4]
  wire  x433_rdcol_1_io_flow; // @[Math.scala 150:24:@25946.4]
  wire [31:0] x433_rdcol_1_io_result; // @[Math.scala 150:24:@25946.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@25966.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@25966.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@25966.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@25966.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@25966.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@25998.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@25998.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@25998.4]
  wire [31:0] RetimeWrapper_43_io_in; // @[package.scala 93:22:@25998.4]
  wire [31:0] RetimeWrapper_43_io_out; // @[package.scala 93:22:@25998.4]
  wire  x439_sum_1_clock; // @[Math.scala 150:24:@26007.4]
  wire  x439_sum_1_reset; // @[Math.scala 150:24:@26007.4]
  wire [31:0] x439_sum_1_io_a; // @[Math.scala 150:24:@26007.4]
  wire [31:0] x439_sum_1_io_b; // @[Math.scala 150:24:@26007.4]
  wire  x439_sum_1_io_flow; // @[Math.scala 150:24:@26007.4]
  wire [31:0] x439_sum_1_io_result; // @[Math.scala 150:24:@26007.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@26017.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@26017.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@26017.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@26017.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@26017.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@26026.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@26026.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@26026.4]
  wire [31:0] RetimeWrapper_45_io_in; // @[package.scala 93:22:@26026.4]
  wire [31:0] RetimeWrapper_45_io_out; // @[package.scala 93:22:@26026.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@26035.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@26035.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@26035.4]
  wire [31:0] RetimeWrapper_46_io_in; // @[package.scala 93:22:@26035.4]
  wire [31:0] RetimeWrapper_46_io_out; // @[package.scala 93:22:@26035.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@26047.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@26047.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@26047.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@26047.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@26047.4]
  wire  x442_rdrow_1_clock; // @[Math.scala 191:24:@26072.4]
  wire  x442_rdrow_1_reset; // @[Math.scala 191:24:@26072.4]
  wire [31:0] x442_rdrow_1_io_a; // @[Math.scala 191:24:@26072.4]
  wire [31:0] x442_rdrow_1_io_b; // @[Math.scala 191:24:@26072.4]
  wire  x442_rdrow_1_io_flow; // @[Math.scala 191:24:@26072.4]
  wire [31:0] x442_rdrow_1_io_result; // @[Math.scala 191:24:@26072.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@26103.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@26103.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@26103.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@26103.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@26103.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@26137.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@26137.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@26137.4]
  wire [40:0] RetimeWrapper_49_io_in; // @[package.scala 93:22:@26137.4]
  wire [40:0] RetimeWrapper_49_io_out; // @[package.scala 93:22:@26137.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@26149.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@26149.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@26149.4]
  wire [36:0] RetimeWrapper_50_io_in; // @[package.scala 93:22:@26149.4]
  wire [36:0] RetimeWrapper_50_io_out; // @[package.scala 93:22:@26149.4]
  wire  x601_sub_1_clock; // @[Math.scala 191:24:@26159.4]
  wire  x601_sub_1_reset; // @[Math.scala 191:24:@26159.4]
  wire [31:0] x601_sub_1_io_a; // @[Math.scala 191:24:@26159.4]
  wire [31:0] x601_sub_1_io_b; // @[Math.scala 191:24:@26159.4]
  wire  x601_sub_1_io_flow; // @[Math.scala 191:24:@26159.4]
  wire [31:0] x601_sub_1_io_result; // @[Math.scala 191:24:@26159.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@26169.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@26169.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@26169.4]
  wire [31:0] RetimeWrapper_51_io_in; // @[package.scala 93:22:@26169.4]
  wire [31:0] RetimeWrapper_51_io_out; // @[package.scala 93:22:@26169.4]
  wire  x450_sum_1_clock; // @[Math.scala 150:24:@26178.4]
  wire  x450_sum_1_reset; // @[Math.scala 150:24:@26178.4]
  wire [31:0] x450_sum_1_io_a; // @[Math.scala 150:24:@26178.4]
  wire [31:0] x450_sum_1_io_b; // @[Math.scala 150:24:@26178.4]
  wire  x450_sum_1_io_flow; // @[Math.scala 150:24:@26178.4]
  wire [31:0] x450_sum_1_io_result; // @[Math.scala 150:24:@26178.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@26188.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@26188.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@26188.4]
  wire [31:0] RetimeWrapper_52_io_in; // @[package.scala 93:22:@26188.4]
  wire [31:0] RetimeWrapper_52_io_out; // @[package.scala 93:22:@26188.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@26197.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@26197.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@26197.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@26197.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@26197.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@26206.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@26206.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@26206.4]
  wire [31:0] RetimeWrapper_54_io_in; // @[package.scala 93:22:@26206.4]
  wire [31:0] RetimeWrapper_54_io_out; // @[package.scala 93:22:@26206.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@26218.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@26218.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@26218.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@26218.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@26218.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@26239.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@26239.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@26239.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@26239.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@26239.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@26251.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@26251.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@26251.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@26251.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@26251.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@26263.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@26263.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@26263.4]
  wire [31:0] RetimeWrapper_58_io_in; // @[package.scala 93:22:@26263.4]
  wire [31:0] RetimeWrapper_58_io_out; // @[package.scala 93:22:@26263.4]
  wire  x455_sum_1_clock; // @[Math.scala 150:24:@26272.4]
  wire  x455_sum_1_reset; // @[Math.scala 150:24:@26272.4]
  wire [31:0] x455_sum_1_io_a; // @[Math.scala 150:24:@26272.4]
  wire [31:0] x455_sum_1_io_b; // @[Math.scala 150:24:@26272.4]
  wire  x455_sum_1_io_flow; // @[Math.scala 150:24:@26272.4]
  wire [31:0] x455_sum_1_io_result; // @[Math.scala 150:24:@26272.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@26282.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@26282.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@26282.4]
  wire [31:0] RetimeWrapper_59_io_in; // @[package.scala 93:22:@26282.4]
  wire [31:0] RetimeWrapper_59_io_out; // @[package.scala 93:22:@26282.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@26291.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@26291.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@26291.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@26291.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@26291.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@26303.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@26303.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@26303.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@26303.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@26303.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@26327.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@26327.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@26327.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@26327.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@26327.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@26339.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@26339.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@26339.4]
  wire [31:0] RetimeWrapper_63_io_in; // @[package.scala 93:22:@26339.4]
  wire [31:0] RetimeWrapper_63_io_out; // @[package.scala 93:22:@26339.4]
  wire  x460_sum_1_clock; // @[Math.scala 150:24:@26348.4]
  wire  x460_sum_1_reset; // @[Math.scala 150:24:@26348.4]
  wire [31:0] x460_sum_1_io_a; // @[Math.scala 150:24:@26348.4]
  wire [31:0] x460_sum_1_io_b; // @[Math.scala 150:24:@26348.4]
  wire  x460_sum_1_io_flow; // @[Math.scala 150:24:@26348.4]
  wire [31:0] x460_sum_1_io_result; // @[Math.scala 150:24:@26348.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@26358.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@26358.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@26358.4]
  wire [31:0] RetimeWrapper_64_io_in; // @[package.scala 93:22:@26358.4]
  wire [31:0] RetimeWrapper_64_io_out; // @[package.scala 93:22:@26358.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@26367.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@26367.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@26367.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@26367.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@26367.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@26379.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@26379.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@26379.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@26379.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@26379.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@26403.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@26403.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@26403.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@26403.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@26403.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@26415.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@26415.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@26415.4]
  wire [31:0] RetimeWrapper_68_io_in; // @[package.scala 93:22:@26415.4]
  wire [31:0] RetimeWrapper_68_io_out; // @[package.scala 93:22:@26415.4]
  wire  x465_sum_1_clock; // @[Math.scala 150:24:@26424.4]
  wire  x465_sum_1_reset; // @[Math.scala 150:24:@26424.4]
  wire [31:0] x465_sum_1_io_a; // @[Math.scala 150:24:@26424.4]
  wire [31:0] x465_sum_1_io_b; // @[Math.scala 150:24:@26424.4]
  wire  x465_sum_1_io_flow; // @[Math.scala 150:24:@26424.4]
  wire [31:0] x465_sum_1_io_result; // @[Math.scala 150:24:@26424.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@26434.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@26434.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@26434.4]
  wire [31:0] RetimeWrapper_69_io_in; // @[package.scala 93:22:@26434.4]
  wire [31:0] RetimeWrapper_69_io_out; // @[package.scala 93:22:@26434.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@26443.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@26443.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@26443.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@26443.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@26443.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@26455.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@26455.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@26455.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@26455.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@26455.4]
  wire  x468_rdrow_1_clock; // @[Math.scala 191:24:@26480.4]
  wire  x468_rdrow_1_reset; // @[Math.scala 191:24:@26480.4]
  wire [31:0] x468_rdrow_1_io_a; // @[Math.scala 191:24:@26480.4]
  wire [31:0] x468_rdrow_1_io_b; // @[Math.scala 191:24:@26480.4]
  wire  x468_rdrow_1_io_flow; // @[Math.scala 191:24:@26480.4]
  wire [31:0] x468_rdrow_1_io_result; // @[Math.scala 191:24:@26480.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@26511.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@26511.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@26511.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@26511.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@26511.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@26545.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@26545.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@26545.4]
  wire [40:0] RetimeWrapper_73_io_in; // @[package.scala 93:22:@26545.4]
  wire [40:0] RetimeWrapper_73_io_out; // @[package.scala 93:22:@26545.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@26557.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@26557.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@26557.4]
  wire [36:0] RetimeWrapper_74_io_in; // @[package.scala 93:22:@26557.4]
  wire [36:0] RetimeWrapper_74_io_out; // @[package.scala 93:22:@26557.4]
  wire  x606_sub_1_clock; // @[Math.scala 191:24:@26567.4]
  wire  x606_sub_1_reset; // @[Math.scala 191:24:@26567.4]
  wire [31:0] x606_sub_1_io_a; // @[Math.scala 191:24:@26567.4]
  wire [31:0] x606_sub_1_io_b; // @[Math.scala 191:24:@26567.4]
  wire  x606_sub_1_io_flow; // @[Math.scala 191:24:@26567.4]
  wire [31:0] x606_sub_1_io_result; // @[Math.scala 191:24:@26567.4]
  wire  x476_sum_1_clock; // @[Math.scala 150:24:@26577.4]
  wire  x476_sum_1_reset; // @[Math.scala 150:24:@26577.4]
  wire [31:0] x476_sum_1_io_a; // @[Math.scala 150:24:@26577.4]
  wire [31:0] x476_sum_1_io_b; // @[Math.scala 150:24:@26577.4]
  wire  x476_sum_1_io_flow; // @[Math.scala 150:24:@26577.4]
  wire [31:0] x476_sum_1_io_result; // @[Math.scala 150:24:@26577.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@26587.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@26587.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@26587.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@26587.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@26587.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@26596.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@26596.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@26596.4]
  wire [31:0] RetimeWrapper_76_io_in; // @[package.scala 93:22:@26596.4]
  wire [31:0] RetimeWrapper_76_io_out; // @[package.scala 93:22:@26596.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@26605.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@26605.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@26605.4]
  wire [31:0] RetimeWrapper_77_io_in; // @[package.scala 93:22:@26605.4]
  wire [31:0] RetimeWrapper_77_io_out; // @[package.scala 93:22:@26605.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@26617.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@26617.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@26617.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@26617.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@26617.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@26641.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@26641.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@26641.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@26641.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@26641.4]
  wire  x481_sum_1_clock; // @[Math.scala 150:24:@26653.4]
  wire  x481_sum_1_reset; // @[Math.scala 150:24:@26653.4]
  wire [31:0] x481_sum_1_io_a; // @[Math.scala 150:24:@26653.4]
  wire [31:0] x481_sum_1_io_b; // @[Math.scala 150:24:@26653.4]
  wire  x481_sum_1_io_flow; // @[Math.scala 150:24:@26653.4]
  wire [31:0] x481_sum_1_io_result; // @[Math.scala 150:24:@26653.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@26663.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@26663.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@26663.4]
  wire [31:0] RetimeWrapper_80_io_in; // @[package.scala 93:22:@26663.4]
  wire [31:0] RetimeWrapper_80_io_out; // @[package.scala 93:22:@26663.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@26672.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@26672.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@26672.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@26672.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@26672.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@26684.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@26684.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@26684.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@26684.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@26684.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@26708.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@26708.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@26708.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@26708.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@26708.4]
  wire  x486_sum_1_clock; // @[Math.scala 150:24:@26720.4]
  wire  x486_sum_1_reset; // @[Math.scala 150:24:@26720.4]
  wire [31:0] x486_sum_1_io_a; // @[Math.scala 150:24:@26720.4]
  wire [31:0] x486_sum_1_io_b; // @[Math.scala 150:24:@26720.4]
  wire  x486_sum_1_io_flow; // @[Math.scala 150:24:@26720.4]
  wire [31:0] x486_sum_1_io_result; // @[Math.scala 150:24:@26720.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@26730.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@26730.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@26730.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@26730.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@26730.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@26739.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@26739.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@26739.4]
  wire [31:0] RetimeWrapper_85_io_in; // @[package.scala 93:22:@26739.4]
  wire [31:0] RetimeWrapper_85_io_out; // @[package.scala 93:22:@26739.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@26751.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@26751.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@26751.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@26751.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@26751.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@26775.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@26775.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@26775.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@26775.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@26775.4]
  wire  x491_sum_1_clock; // @[Math.scala 150:24:@26787.4]
  wire  x491_sum_1_reset; // @[Math.scala 150:24:@26787.4]
  wire [31:0] x491_sum_1_io_a; // @[Math.scala 150:24:@26787.4]
  wire [31:0] x491_sum_1_io_b; // @[Math.scala 150:24:@26787.4]
  wire  x491_sum_1_io_flow; // @[Math.scala 150:24:@26787.4]
  wire [31:0] x491_sum_1_io_result; // @[Math.scala 150:24:@26787.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@26797.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@26797.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@26797.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@26797.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@26797.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@26806.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@26806.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@26806.4]
  wire [31:0] RetimeWrapper_89_io_in; // @[package.scala 93:22:@26806.4]
  wire [31:0] RetimeWrapper_89_io_out; // @[package.scala 93:22:@26806.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@26818.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@26818.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@26818.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@26818.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@26818.4]
  wire [7:0] x499_x15_1_io_a; // @[Math.scala 150:24:@26864.4]
  wire [7:0] x499_x15_1_io_b; // @[Math.scala 150:24:@26864.4]
  wire [7:0] x499_x15_1_io_result; // @[Math.scala 150:24:@26864.4]
  wire [7:0] x500_x16_1_io_a; // @[Math.scala 150:24:@26876.4]
  wire [7:0] x500_x16_1_io_b; // @[Math.scala 150:24:@26876.4]
  wire [7:0] x500_x16_1_io_result; // @[Math.scala 150:24:@26876.4]
  wire [7:0] x501_x15_1_io_a; // @[Math.scala 150:24:@26886.4]
  wire [7:0] x501_x15_1_io_b; // @[Math.scala 150:24:@26886.4]
  wire [7:0] x501_x15_1_io_result; // @[Math.scala 150:24:@26886.4]
  wire [7:0] x502_x16_1_io_a; // @[Math.scala 150:24:@26896.4]
  wire [7:0] x502_x16_1_io_b; // @[Math.scala 150:24:@26896.4]
  wire [7:0] x502_x16_1_io_result; // @[Math.scala 150:24:@26896.4]
  wire [7:0] x503_x15_1_io_a; // @[Math.scala 150:24:@26906.4]
  wire [7:0] x503_x15_1_io_b; // @[Math.scala 150:24:@26906.4]
  wire [7:0] x503_x15_1_io_result; // @[Math.scala 150:24:@26906.4]
  wire [7:0] x504_x16_1_io_a; // @[Math.scala 150:24:@26916.4]
  wire [7:0] x504_x16_1_io_b; // @[Math.scala 150:24:@26916.4]
  wire [7:0] x504_x16_1_io_result; // @[Math.scala 150:24:@26916.4]
  wire [7:0] x505_x15_1_io_a; // @[Math.scala 150:24:@26926.4]
  wire [7:0] x505_x15_1_io_b; // @[Math.scala 150:24:@26926.4]
  wire [7:0] x505_x15_1_io_result; // @[Math.scala 150:24:@26926.4]
  wire  x506_sum_1_clock; // @[Math.scala 150:24:@26936.4]
  wire  x506_sum_1_reset; // @[Math.scala 150:24:@26936.4]
  wire [7:0] x506_sum_1_io_a; // @[Math.scala 150:24:@26936.4]
  wire [7:0] x506_sum_1_io_b; // @[Math.scala 150:24:@26936.4]
  wire  x506_sum_1_io_flow; // @[Math.scala 150:24:@26936.4]
  wire [7:0] x506_sum_1_io_result; // @[Math.scala 150:24:@26936.4]
  wire [7:0] x513_x15_1_io_a; // @[Math.scala 150:24:@26978.4]
  wire [7:0] x513_x15_1_io_b; // @[Math.scala 150:24:@26978.4]
  wire [7:0] x513_x15_1_io_result; // @[Math.scala 150:24:@26978.4]
  wire [7:0] x514_x16_1_io_a; // @[Math.scala 150:24:@26988.4]
  wire [7:0] x514_x16_1_io_b; // @[Math.scala 150:24:@26988.4]
  wire [7:0] x514_x16_1_io_result; // @[Math.scala 150:24:@26988.4]
  wire [7:0] x515_x15_1_io_a; // @[Math.scala 150:24:@26998.4]
  wire [7:0] x515_x15_1_io_b; // @[Math.scala 150:24:@26998.4]
  wire [7:0] x515_x15_1_io_result; // @[Math.scala 150:24:@26998.4]
  wire [7:0] x516_x16_1_io_a; // @[Math.scala 150:24:@27008.4]
  wire [7:0] x516_x16_1_io_b; // @[Math.scala 150:24:@27008.4]
  wire [7:0] x516_x16_1_io_result; // @[Math.scala 150:24:@27008.4]
  wire [7:0] x517_x15_1_io_a; // @[Math.scala 150:24:@27018.4]
  wire [7:0] x517_x15_1_io_b; // @[Math.scala 150:24:@27018.4]
  wire [7:0] x517_x15_1_io_result; // @[Math.scala 150:24:@27018.4]
  wire [7:0] x518_x16_1_io_a; // @[Math.scala 150:24:@27028.4]
  wire [7:0] x518_x16_1_io_b; // @[Math.scala 150:24:@27028.4]
  wire [7:0] x518_x16_1_io_result; // @[Math.scala 150:24:@27028.4]
  wire [7:0] x519_x15_1_io_a; // @[Math.scala 150:24:@27038.4]
  wire [7:0] x519_x15_1_io_b; // @[Math.scala 150:24:@27038.4]
  wire [7:0] x519_x15_1_io_result; // @[Math.scala 150:24:@27038.4]
  wire  x520_sum_1_clock; // @[Math.scala 150:24:@27048.4]
  wire  x520_sum_1_reset; // @[Math.scala 150:24:@27048.4]
  wire [7:0] x520_sum_1_io_a; // @[Math.scala 150:24:@27048.4]
  wire [7:0] x520_sum_1_io_b; // @[Math.scala 150:24:@27048.4]
  wire  x520_sum_1_io_flow; // @[Math.scala 150:24:@27048.4]
  wire [7:0] x520_sum_1_io_result; // @[Math.scala 150:24:@27048.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@27071.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@27071.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@27071.4]
  wire [15:0] RetimeWrapper_91_io_in; // @[package.scala 93:22:@27071.4]
  wire [15:0] RetimeWrapper_91_io_out; // @[package.scala 93:22:@27071.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@27080.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@27080.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@27080.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@27080.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@27080.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@27089.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@27089.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@27089.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@27089.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@27089.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@27098.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@27098.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@27098.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@27098.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@27098.4]
  wire  b381; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 62:18:@25056.4]
  wire  b382; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 63:18:@25057.4]
  wire  _T_205; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 67:30:@25059.4]
  wire  _T_206; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 67:37:@25060.4]
  wire  _T_210; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 69:76:@25065.4]
  wire  _T_211; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 69:62:@25066.4]
  wire  _T_213; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 69:101:@25067.4]
  wire [15:0] x612_x383_D1_0_number; // @[package.scala 96:25:@25076.4 package.scala 96:25:@25077.4]
  wire [31:0] b379_number; // @[Math.scala 712:22:@25041.4 Math.scala 713:14:@25042.4]
  wire [31:0] _T_242; // @[Math.scala 499:52:@25185.4]
  wire  x388; // @[Math.scala 499:44:@25193.4]
  wire  x389; // @[Math.scala 499:44:@25200.4]
  wire  x390; // @[Math.scala 499:44:@25207.4]
  wire [31:0] _T_289; // @[Mux.scala 19:72:@25219.4]
  wire [31:0] _T_291; // @[Mux.scala 19:72:@25220.4]
  wire [31:0] _T_293; // @[Mux.scala 19:72:@25221.4]
  wire [31:0] _T_295; // @[Mux.scala 19:72:@25223.4]
  wire [31:0] x613_x391_D2_number; // @[package.scala 96:25:@25236.4 package.scala 96:25:@25237.4]
  wire [31:0] _T_310; // @[Math.scala 406:49:@25243.4]
  wire [31:0] _T_312; // @[Math.scala 406:56:@25245.4]
  wire [31:0] _T_313; // @[Math.scala 406:56:@25246.4]
  wire [31:0] b380_number; // @[Math.scala 712:22:@25053.4 Math.scala 713:14:@25054.4]
  wire [31:0] _T_322; // @[Math.scala 406:49:@25254.4]
  wire [31:0] _T_324; // @[Math.scala 406:56:@25256.4]
  wire [31:0] _T_325; // @[Math.scala 406:56:@25257.4]
  wire  _T_330; // @[FixedPoint.scala 50:25:@25263.4]
  wire [1:0] _T_334; // @[Bitwise.scala 72:12:@25265.4]
  wire [29:0] _T_335; // @[FixedPoint.scala 18:52:@25266.4]
  wire [31:0] x395_number; // @[Cat.scala 30:58:@25267.4]
  wire [40:0] _GEN_0; // @[Math.scala 450:32:@25272.4]
  wire [40:0] _T_340; // @[Math.scala 450:32:@25272.4]
  wire [36:0] _GEN_1; // @[Math.scala 450:32:@25277.4]
  wire [36:0] _T_344; // @[Math.scala 450:32:@25277.4]
  wire  _T_351; // @[FixedPoint.scala 50:25:@25292.4]
  wire [1:0] _T_355; // @[Bitwise.scala 72:12:@25294.4]
  wire [29:0] _T_356; // @[FixedPoint.scala 18:52:@25295.4]
  wire  _T_383; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 127:101:@25372.4]
  wire  _T_387; // @[package.scala 96:25:@25380.4 package.scala 96:25:@25381.4]
  wire  _T_389; // @[implicits.scala 55:10:@25382.4]
  wire  _T_390; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 127:118:@25383.4]
  wire  _T_392; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 127:206:@25385.4]
  wire  _T_393; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 127:225:@25386.4]
  wire  x615_b381_D5; // @[package.scala 96:25:@25324.4 package.scala 96:25:@25325.4]
  wire  _T_394; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 127:251:@25387.4]
  wire  x619_b382_D5; // @[package.scala 96:25:@25360.4 package.scala 96:25:@25361.4]
  wire [31:0] x400_rdcol_number; // @[Math.scala 154:22:@25404.4 Math.scala 155:14:@25405.4]
  wire [31:0] _T_411; // @[Math.scala 406:49:@25413.4]
  wire [31:0] _T_413; // @[Math.scala 406:56:@25415.4]
  wire [31:0] _T_414; // @[Math.scala 406:56:@25416.4]
  wire  _T_419; // @[FixedPoint.scala 50:25:@25422.4]
  wire [1:0] _T_423; // @[Bitwise.scala 72:12:@25424.4]
  wire [29:0] _T_424; // @[FixedPoint.scala 18:52:@25425.4]
  wire  _T_446; // @[package.scala 96:25:@25483.4 package.scala 96:25:@25484.4]
  wire  _T_448; // @[implicits.scala 55:10:@25485.4]
  wire  _T_449; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 150:118:@25486.4]
  wire  _T_451; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 150:206:@25488.4]
  wire  _T_452; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 150:225:@25489.4]
  wire  _T_453; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 150:251:@25490.4]
  wire [31:0] x625_b379_D8_number; // @[package.scala 96:25:@25504.4 package.scala 96:25:@25505.4]
  wire [31:0] _T_465; // @[Math.scala 406:49:@25511.4]
  wire [31:0] _T_467; // @[Math.scala 406:56:@25513.4]
  wire [31:0] _T_468; // @[Math.scala 406:56:@25514.4]
  wire [31:0] x590_number; // @[implicits.scala 133:21:@25515.4]
  wire  x408; // @[Math.scala 465:44:@25523.4]
  wire [31:0] x626_x400_rdcol_D8_number; // @[package.scala 96:25:@25531.4 package.scala 96:25:@25532.4]
  wire [31:0] _T_486; // @[Math.scala 465:37:@25537.4]
  wire  x409; // @[Math.scala 465:44:@25539.4]
  wire  x627_x408_D1; // @[package.scala 96:25:@25547.4 package.scala 96:25:@25548.4]
  wire  x628_x410_D1; // @[package.scala 96:25:@25559.4 package.scala 96:25:@25560.4]
  wire [31:0] _T_506; // @[Math.scala 406:49:@25569.4]
  wire [31:0] _T_508; // @[Math.scala 406:56:@25571.4]
  wire [31:0] _T_509; // @[Math.scala 406:56:@25572.4]
  wire  _T_516; // @[FixedPoint.scala 50:25:@25580.4]
  wire [1:0] _T_520; // @[Bitwise.scala 72:12:@25582.4]
  wire [29:0] _T_521; // @[FixedPoint.scala 18:52:@25583.4]
  wire [31:0] x413_number; // @[Cat.scala 30:58:@25584.4]
  wire [40:0] _GEN_2; // @[Math.scala 450:32:@25589.4]
  wire [36:0] _GEN_3; // @[Math.scala 450:32:@25601.4]
  wire  _T_573; // @[package.scala 96:25:@25703.4 package.scala 96:25:@25704.4]
  wire  _T_575; // @[implicits.scala 55:10:@25705.4]
  wire  _T_576; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 208:194:@25706.4]
  wire  x631_x411_D4; // @[package.scala 96:25:@25655.4 package.scala 96:25:@25656.4]
  wire  _T_577; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 208:283:@25707.4]
  wire  x632_b381_D14; // @[package.scala 96:25:@25664.4 package.scala 96:25:@25665.4]
  wire  _T_578; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 208:291:@25708.4]
  wire  x633_b382_D14; // @[package.scala 96:25:@25673.4 package.scala 96:25:@25674.4]
  wire [31:0] x636_b380_D8_number; // @[package.scala 96:25:@25724.4 package.scala 96:25:@25725.4]
  wire [31:0] _T_589; // @[Math.scala 465:37:@25730.4]
  wire  x418; // @[Math.scala 465:44:@25732.4]
  wire  x637_x419_D1; // @[package.scala 96:25:@25743.4 package.scala 96:25:@25744.4]
  wire  _T_625; // @[package.scala 96:25:@25804.4 package.scala 96:25:@25805.4]
  wire  _T_627; // @[implicits.scala 55:10:@25806.4]
  wire  _T_628; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 235:194:@25807.4]
  wire  x640_x420_D5; // @[package.scala 96:25:@25783.4 package.scala 96:25:@25784.4]
  wire  _T_629; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 235:283:@25808.4]
  wire  _T_630; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 235:291:@25809.4]
  wire [31:0] x424_rdcol_number; // @[Math.scala 154:22:@25828.4 Math.scala 155:14:@25829.4]
  wire [31:0] _T_645; // @[Math.scala 465:37:@25834.4]
  wire  x425; // @[Math.scala 465:44:@25836.4]
  wire  x642_x426_D1; // @[package.scala 96:25:@25847.4 package.scala 96:25:@25848.4]
  wire [31:0] _T_664; // @[Math.scala 406:56:@25859.4]
  wire [31:0] _T_665; // @[Math.scala 406:56:@25860.4]
  wire  _T_670; // @[FixedPoint.scala 50:25:@25866.4]
  wire [1:0] _T_674; // @[Bitwise.scala 72:12:@25868.4]
  wire [29:0] _T_675; // @[FixedPoint.scala 18:52:@25869.4]
  wire  _T_703; // @[package.scala 96:25:@25928.4 package.scala 96:25:@25929.4]
  wire  _T_705; // @[implicits.scala 55:10:@25930.4]
  wire  _T_706; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 266:194:@25931.4]
  wire  x646_x427_D4; // @[package.scala 96:25:@25916.4 package.scala 96:25:@25917.4]
  wire  _T_707; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 266:283:@25932.4]
  wire  _T_708; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 266:291:@25933.4]
  wire [31:0] x433_rdcol_number; // @[Math.scala 154:22:@25952.4 Math.scala 155:14:@25953.4]
  wire [31:0] _T_723; // @[Math.scala 465:37:@25958.4]
  wire  x434; // @[Math.scala 465:44:@25960.4]
  wire  x647_x435_D1; // @[package.scala 96:25:@25971.4 package.scala 96:25:@25972.4]
  wire [31:0] _T_742; // @[Math.scala 406:56:@25983.4]
  wire [31:0] _T_743; // @[Math.scala 406:56:@25984.4]
  wire  _T_748; // @[FixedPoint.scala 50:25:@25990.4]
  wire [1:0] _T_752; // @[Bitwise.scala 72:12:@25992.4]
  wire [29:0] _T_753; // @[FixedPoint.scala 18:52:@25993.4]
  wire  _T_781; // @[package.scala 96:25:@26052.4 package.scala 96:25:@26053.4]
  wire  _T_783; // @[implicits.scala 55:10:@26054.4]
  wire  _T_784; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 303:194:@26055.4]
  wire  x649_x436_D4; // @[package.scala 96:25:@26022.4 package.scala 96:25:@26023.4]
  wire  _T_785; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 303:283:@26056.4]
  wire  _T_786; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 303:291:@26057.4]
  wire [31:0] x442_rdrow_number; // @[Math.scala 195:22:@26078.4 Math.scala 196:14:@26079.4]
  wire [31:0] _T_805; // @[Math.scala 406:49:@26085.4]
  wire [31:0] _T_807; // @[Math.scala 406:56:@26087.4]
  wire [31:0] _T_808; // @[Math.scala 406:56:@26088.4]
  wire [31:0] x597_number; // @[implicits.scala 133:21:@26089.4]
  wire  x444; // @[Math.scala 465:44:@26097.4]
  wire  x652_x445_D1; // @[package.scala 96:25:@26108.4 package.scala 96:25:@26109.4]
  wire [31:0] _T_832; // @[Math.scala 406:49:@26118.4]
  wire [31:0] _T_834; // @[Math.scala 406:56:@26120.4]
  wire [31:0] _T_835; // @[Math.scala 406:56:@26121.4]
  wire  _T_840; // @[FixedPoint.scala 50:25:@26127.4]
  wire [1:0] _T_844; // @[Bitwise.scala 72:12:@26129.4]
  wire [29:0] _T_845; // @[FixedPoint.scala 18:52:@26130.4]
  wire [31:0] x448_number; // @[Cat.scala 30:58:@26131.4]
  wire [40:0] _GEN_4; // @[Math.scala 450:32:@26136.4]
  wire [36:0] _GEN_5; // @[Math.scala 450:32:@26148.4]
  wire  _T_888; // @[package.scala 96:25:@26223.4 package.scala 96:25:@26224.4]
  wire  _T_890; // @[implicits.scala 55:10:@26225.4]
  wire  _T_891; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 344:194:@26226.4]
  wire  x655_x446_D4; // @[package.scala 96:25:@26202.4 package.scala 96:25:@26203.4]
  wire  _T_892; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 344:283:@26227.4]
  wire  _T_893; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 344:291:@26228.4]
  wire  x657_x418_D1; // @[package.scala 96:25:@26244.4 package.scala 96:25:@26245.4]
  wire  x658_x453_D1; // @[package.scala 96:25:@26256.4 package.scala 96:25:@26257.4]
  wire  _T_929; // @[package.scala 96:25:@26308.4 package.scala 96:25:@26309.4]
  wire  _T_931; // @[implicits.scala 55:10:@26310.4]
  wire  _T_932; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 367:194:@26311.4]
  wire  x661_x454_D4; // @[package.scala 96:25:@26296.4 package.scala 96:25:@26297.4]
  wire  _T_933; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 367:283:@26312.4]
  wire  _T_934; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 367:291:@26313.4]
  wire  x662_x458_D1; // @[package.scala 96:25:@26332.4 package.scala 96:25:@26333.4]
  wire  _T_967; // @[package.scala 96:25:@26384.4 package.scala 96:25:@26385.4]
  wire  _T_969; // @[implicits.scala 55:10:@26386.4]
  wire  _T_970; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 388:194:@26387.4]
  wire  x665_x459_D4; // @[package.scala 96:25:@26372.4 package.scala 96:25:@26373.4]
  wire  _T_971; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 388:283:@26388.4]
  wire  _T_972; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 388:291:@26389.4]
  wire  x666_x463_D1; // @[package.scala 96:25:@26408.4 package.scala 96:25:@26409.4]
  wire  _T_1005; // @[package.scala 96:25:@26460.4 package.scala 96:25:@26461.4]
  wire  _T_1007; // @[implicits.scala 55:10:@26462.4]
  wire  _T_1008; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 415:194:@26463.4]
  wire  x669_x464_D4; // @[package.scala 96:25:@26448.4 package.scala 96:25:@26449.4]
  wire  _T_1009; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 415:283:@26464.4]
  wire  _T_1010; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 415:326:@26465.4]
  wire [31:0] x468_rdrow_number; // @[Math.scala 195:22:@26486.4 Math.scala 196:14:@26487.4]
  wire [31:0] _T_1029; // @[Math.scala 406:49:@26493.4]
  wire [31:0] _T_1031; // @[Math.scala 406:56:@26495.4]
  wire [31:0] _T_1032; // @[Math.scala 406:56:@26496.4]
  wire [31:0] x602_number; // @[implicits.scala 133:21:@26497.4]
  wire  x470; // @[Math.scala 465:44:@26505.4]
  wire  x670_x471_D1; // @[package.scala 96:25:@26516.4 package.scala 96:25:@26517.4]
  wire [31:0] _T_1056; // @[Math.scala 406:49:@26526.4]
  wire [31:0] _T_1058; // @[Math.scala 406:56:@26528.4]
  wire [31:0] _T_1059; // @[Math.scala 406:56:@26529.4]
  wire  _T_1064; // @[FixedPoint.scala 50:25:@26535.4]
  wire [1:0] _T_1068; // @[Bitwise.scala 72:12:@26537.4]
  wire [29:0] _T_1069; // @[FixedPoint.scala 18:52:@26538.4]
  wire [31:0] x474_number; // @[Cat.scala 30:58:@26539.4]
  wire [40:0] _GEN_6; // @[Math.scala 450:32:@26544.4]
  wire [36:0] _GEN_7; // @[Math.scala 450:32:@26556.4]
  wire  _T_1109; // @[package.scala 96:25:@26622.4 package.scala 96:25:@26623.4]
  wire  _T_1111; // @[implicits.scala 55:10:@26624.4]
  wire  _T_1112; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 454:194:@26625.4]
  wire  x671_x472_D4; // @[package.scala 96:25:@26592.4 package.scala 96:25:@26593.4]
  wire  _T_1113; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 454:283:@26626.4]
  wire  _T_1114; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 454:291:@26627.4]
  wire  x674_x479_D1; // @[package.scala 96:25:@26646.4 package.scala 96:25:@26647.4]
  wire  _T_1144; // @[package.scala 96:25:@26689.4 package.scala 96:25:@26690.4]
  wire  _T_1146; // @[implicits.scala 55:10:@26691.4]
  wire  _T_1147; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 473:194:@26692.4]
  wire  x676_x480_D4; // @[package.scala 96:25:@26677.4 package.scala 96:25:@26678.4]
  wire  _T_1148; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 473:283:@26693.4]
  wire  _T_1149; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 473:291:@26694.4]
  wire  x677_x484_D1; // @[package.scala 96:25:@26713.4 package.scala 96:25:@26714.4]
  wire  _T_1179; // @[package.scala 96:25:@26756.4 package.scala 96:25:@26757.4]
  wire  _T_1181; // @[implicits.scala 55:10:@26758.4]
  wire  _T_1182; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 492:194:@26759.4]
  wire  x678_x485_D4; // @[package.scala 96:25:@26735.4 package.scala 96:25:@26736.4]
  wire  _T_1183; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 492:283:@26760.4]
  wire  _T_1184; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 492:291:@26761.4]
  wire  x680_x489_D1; // @[package.scala 96:25:@26780.4 package.scala 96:25:@26781.4]
  wire  _T_1214; // @[package.scala 96:25:@26823.4 package.scala 96:25:@26824.4]
  wire  _T_1216; // @[implicits.scala 55:10:@26825.4]
  wire  _T_1217; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 511:194:@26826.4]
  wire  x681_x490_D4; // @[package.scala 96:25:@26802.4 package.scala 96:25:@26803.4]
  wire  _T_1218; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 511:283:@26827.4]
  wire  _T_1219; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 511:291:@26828.4]
  wire [7:0] x422_rd_0_number; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 231:29:@25795.4 sm_x526_inr_Foreach_SAMPLER_BOX.scala 235:338:@25816.4]
  wire [8:0] _GEN_8; // @[Math.scala 450:32:@26840.4]
  wire [8:0] _T_1225; // @[Math.scala 450:32:@26840.4]
  wire [7:0] x451_rd_0_number; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 340:29:@26214.4 sm_x526_inr_Foreach_SAMPLER_BOX.scala 344:408:@26235.4]
  wire [8:0] _GEN_9; // @[Math.scala 450:32:@26845.4]
  wire [8:0] _T_1229; // @[Math.scala 450:32:@26845.4]
  wire [7:0] x456_rd_0_number; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 363:29:@26299.4 sm_x526_inr_Foreach_SAMPLER_BOX.scala 367:408:@26320.4]
  wire [9:0] _GEN_10; // @[Math.scala 450:32:@26850.4]
  wire [9:0] _T_1233; // @[Math.scala 450:32:@26850.4]
  wire [7:0] x461_rd_0_number; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 384:29:@26375.4 sm_x526_inr_Foreach_SAMPLER_BOX.scala 388:408:@26396.4]
  wire [8:0] _GEN_11; // @[Math.scala 450:32:@26855.4]
  wire [8:0] _T_1237; // @[Math.scala 450:32:@26855.4]
  wire [7:0] x482_rd_0_number; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 469:29:@26680.4 sm_x526_inr_Foreach_SAMPLER_BOX.scala 473:408:@26701.4]
  wire [8:0] _GEN_12; // @[Math.scala 450:32:@26860.4]
  wire [8:0] _T_1241; // @[Math.scala 450:32:@26860.4]
  wire [7:0] x506_sum_number; // @[Math.scala 154:22:@26942.4 Math.scala 155:14:@26943.4]
  wire [3:0] _T_1276; // @[FixedPoint.scala 18:52:@26948.4]
  wire [7:0] x507_number; // @[Cat.scala 30:58:@26949.4]
  wire [7:0] x431_rd_0_number; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 262:29:@25919.4 sm_x526_inr_Foreach_SAMPLER_BOX.scala 266:338:@25940.4]
  wire [8:0] _GEN_13; // @[Math.scala 450:32:@26954.4]
  wire [8:0] _T_1281; // @[Math.scala 450:32:@26954.4]
  wire [8:0] _GEN_14; // @[Math.scala 450:32:@26959.4]
  wire [8:0] _T_1285; // @[Math.scala 450:32:@26959.4]
  wire [9:0] _GEN_15; // @[Math.scala 450:32:@26964.4]
  wire [9:0] _T_1289; // @[Math.scala 450:32:@26964.4]
  wire [7:0] x466_rd_0_number; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 411:29:@26451.4 sm_x526_inr_Foreach_SAMPLER_BOX.scala 415:443:@26472.4]
  wire [8:0] _GEN_16; // @[Math.scala 450:32:@26969.4]
  wire [8:0] _T_1293; // @[Math.scala 450:32:@26969.4]
  wire [7:0] x487_rd_0_number; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 488:29:@26747.4 sm_x526_inr_Foreach_SAMPLER_BOX.scala 492:408:@26768.4]
  wire [8:0] _GEN_17; // @[Math.scala 450:32:@26974.4]
  wire [8:0] _T_1297; // @[Math.scala 450:32:@26974.4]
  wire [7:0] x520_sum_number; // @[Math.scala 154:22:@27054.4 Math.scala 155:14:@27055.4]
  wire [3:0] _T_1330; // @[FixedPoint.scala 18:52:@27060.4]
  wire [7:0] x521_number; // @[Cat.scala 30:58:@27061.4]
  wire  _T_1353; // @[package.scala 96:25:@27103.4 package.scala 96:25:@27104.4]
  wire  _T_1355; // @[implicits.scala 55:10:@27105.4]
  wire  x684_b381_D20; // @[package.scala 96:25:@27094.4 package.scala 96:25:@27095.4]
  wire  _T_1356; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 587:117:@27106.4]
  wire  x683_b382_D20; // @[package.scala 96:25:@27085.4 package.scala 96:25:@27086.4]
  wire  _T_1357; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 587:123:@27107.4]
  wire [31:0] x617_x398_sum_D1_number; // @[package.scala 96:25:@25342.4 package.scala 96:25:@25343.4]
  wire [31:0] x618_x584_D3_number; // @[package.scala 96:25:@25351.4 package.scala 96:25:@25352.4]
  wire [31:0] x620_x585_D5_number; // @[package.scala 96:25:@25369.4 package.scala 96:25:@25370.4]
  wire [31:0] x622_x404_sum_D1_number; // @[package.scala 96:25:@25454.4 package.scala 96:25:@25455.4]
  wire [31:0] x623_x589_D4_number; // @[package.scala 96:25:@25463.4 package.scala 96:25:@25464.4]
  wire [40:0] _T_528; // @[package.scala 96:25:@25595.4 package.scala 96:25:@25596.4]
  wire [36:0] _T_534; // @[package.scala 96:25:@25607.4 package.scala 96:25:@25608.4]
  wire [31:0] x630_x591_D6_number; // @[package.scala 96:25:@25646.4 package.scala 96:25:@25647.4]
  wire [31:0] x634_x589_D13_number; // @[package.scala 96:25:@25682.4 package.scala 96:25:@25683.4]
  wire [31:0] x635_x415_sum_D3_number; // @[package.scala 96:25:@25691.4 package.scala 96:25:@25692.4]
  wire [31:0] x639_x421_sum_D3_number; // @[package.scala 96:25:@25774.4 package.scala 96:25:@25775.4]
  wire [31:0] x641_x585_D14_number; // @[package.scala 96:25:@25792.4 package.scala 96:25:@25793.4]
  wire [31:0] x644_x430_sum_D3_number; // @[package.scala 96:25:@25898.4 package.scala 96:25:@25899.4]
  wire [31:0] x645_x595_D5_number; // @[package.scala 96:25:@25907.4 package.scala 96:25:@25908.4]
  wire [31:0] x650_x439_sum_D3_number; // @[package.scala 96:25:@26031.4 package.scala 96:25:@26032.4]
  wire [31:0] x651_x596_D5_number; // @[package.scala 96:25:@26040.4 package.scala 96:25:@26041.4]
  wire [40:0] _T_852; // @[package.scala 96:25:@26142.4 package.scala 96:25:@26143.4]
  wire [36:0] _T_858; // @[package.scala 96:25:@26154.4 package.scala 96:25:@26155.4]
  wire [31:0] x654_x598_D5_number; // @[package.scala 96:25:@26193.4 package.scala 96:25:@26194.4]
  wire [31:0] x656_x450_sum_D2_number; // @[package.scala 96:25:@26211.4 package.scala 96:25:@26212.4]
  wire [31:0] x660_x455_sum_D2_number; // @[package.scala 96:25:@26287.4 package.scala 96:25:@26288.4]
  wire [31:0] x664_x460_sum_D2_number; // @[package.scala 96:25:@26363.4 package.scala 96:25:@26364.4]
  wire [31:0] x668_x465_sum_D2_number; // @[package.scala 96:25:@26439.4 package.scala 96:25:@26440.4]
  wire [40:0] _T_1076; // @[package.scala 96:25:@26550.4 package.scala 96:25:@26551.4]
  wire [36:0] _T_1082; // @[package.scala 96:25:@26562.4 package.scala 96:25:@26563.4]
  wire [31:0] x672_x476_sum_D2_number; // @[package.scala 96:25:@26601.4 package.scala 96:25:@26602.4]
  wire [31:0] x673_x603_D5_number; // @[package.scala 96:25:@26610.4 package.scala 96:25:@26611.4]
  wire [31:0] x675_x481_sum_D2_number; // @[package.scala 96:25:@26668.4 package.scala 96:25:@26669.4]
  wire [31:0] x679_x486_sum_D2_number; // @[package.scala 96:25:@26744.4 package.scala 96:25:@26745.4]
  wire [31:0] x682_x491_sum_D2_number; // @[package.scala 96:25:@26811.4 package.scala 96:25:@26812.4]
  _ _ ( // @[Math.scala 709:24:@25036.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@25048.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@25071.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x385_lb_0 x385_lb_0 ( // @[m_x385_lb_0.scala 39:17:@25081.4]
    .clock(x385_lb_0_clock),
    .reset(x385_lb_0_reset),
    .io_rPort_11_banks_1(x385_lb_0_io_rPort_11_banks_1),
    .io_rPort_11_banks_0(x385_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x385_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x385_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x385_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x385_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_1(x385_lb_0_io_rPort_10_banks_1),
    .io_rPort_10_banks_0(x385_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x385_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x385_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x385_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x385_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_1(x385_lb_0_io_rPort_9_banks_1),
    .io_rPort_9_banks_0(x385_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x385_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x385_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x385_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x385_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_1(x385_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x385_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x385_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x385_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x385_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x385_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x385_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x385_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x385_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x385_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x385_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x385_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x385_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x385_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x385_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x385_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x385_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x385_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x385_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x385_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x385_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x385_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x385_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x385_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x385_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x385_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x385_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x385_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x385_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x385_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x385_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x385_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x385_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x385_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x385_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x385_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x385_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x385_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x385_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x385_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x385_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x385_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x385_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x385_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x385_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x385_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x385_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x385_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x385_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x385_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x385_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x385_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x385_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x385_lb_0_io_rPort_0_output_0),
    .io_wPort_1_banks_1(x385_lb_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x385_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x385_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x385_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x385_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x385_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x385_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x385_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x385_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x385_lb_0_io_wPort_0_en_0)
  );
  RetimeWrapper_165 RetimeWrapper_1 ( // @[package.scala 93:22:@25231.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x577_sub x588_sub_1 ( // @[Math.scala 191:24:@25281.4]
    .clock(x588_sub_1_clock),
    .reset(x588_sub_1_reset),
    .io_a(x588_sub_1_io_a),
    .io_b(x588_sub_1_io_b),
    .io_flow(x588_sub_1_io_flow),
    .io_result(x588_sub_1_io_result)
  );
  RetimeWrapper_167 RetimeWrapper_2 ( // @[package.scala 93:22:@25300.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x362_sum x398_sum_1 ( // @[Math.scala 150:24:@25309.4]
    .clock(x398_sum_1_clock),
    .reset(x398_sum_1_reset),
    .io_a(x398_sum_1_io_a),
    .io_b(x398_sum_1_io_b),
    .io_flow(x398_sum_1_io_flow),
    .io_result(x398_sum_1_io_result)
  );
  RetimeWrapper_21 RetimeWrapper_3 ( // @[package.scala 93:22:@25319.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_170 RetimeWrapper_4 ( // @[package.scala 93:22:@25328.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_5 ( // @[package.scala 93:22:@25337.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_167 RetimeWrapper_6 ( // @[package.scala 93:22:@25346.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_7 ( // @[package.scala 93:22:@25355.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_174 RetimeWrapper_8 ( // @[package.scala 93:22:@25364.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_9 ( // @[package.scala 93:22:@25375.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  x362_sum x400_rdcol_1 ( // @[Math.scala 150:24:@25398.4]
    .clock(x400_rdcol_1_clock),
    .reset(x400_rdcol_1_reset),
    .io_a(x400_rdcol_1_io_a),
    .io_b(x400_rdcol_1_io_b),
    .io_flow(x400_rdcol_1_io_flow),
    .io_result(x400_rdcol_1_io_result)
  );
  RetimeWrapper_165 RetimeWrapper_10 ( // @[package.scala 93:22:@25430.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  x362_sum x404_sum_1 ( // @[Math.scala 150:24:@25439.4]
    .clock(x404_sum_1_clock),
    .reset(x404_sum_1_reset),
    .io_a(x404_sum_1_io_a),
    .io_b(x404_sum_1_io_b),
    .io_flow(x404_sum_1_io_flow),
    .io_result(x404_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_11 ( // @[package.scala 93:22:@25449.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_180 RetimeWrapper_12 ( // @[package.scala 93:22:@25458.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_170 RetimeWrapper_13 ( // @[package.scala 93:22:@25467.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_14 ( // @[package.scala 93:22:@25478.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_183 RetimeWrapper_15 ( // @[package.scala 93:22:@25499.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_183 RetimeWrapper_16 ( // @[package.scala 93:22:@25526.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper RetimeWrapper_17 ( // @[package.scala 93:22:@25542.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper RetimeWrapper_18 ( // @[package.scala 93:22:@25554.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_187 RetimeWrapper_19 ( // @[package.scala 93:22:@25590.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_188 RetimeWrapper_20 ( // @[package.scala 93:22:@25602.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  x577_sub x594_sub_1 ( // @[Math.scala 191:24:@25612.4]
    .clock(x594_sub_1_clock),
    .reset(x594_sub_1_reset),
    .io_a(x594_sub_1_io_a),
    .io_b(x594_sub_1_io_b),
    .io_flow(x594_sub_1_io_flow),
    .io_result(x594_sub_1_io_result)
  );
  RetimeWrapper_190 RetimeWrapper_21 ( // @[package.scala 93:22:@25622.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  x362_sum x415_sum_1 ( // @[Math.scala 150:24:@25631.4]
    .clock(x415_sum_1_clock),
    .reset(x415_sum_1_reset),
    .io_a(x415_sum_1_io_a),
    .io_b(x415_sum_1_io_b),
    .io_flow(x415_sum_1_io_flow),
    .io_result(x415_sum_1_io_result)
  );
  RetimeWrapper_192 RetimeWrapper_22 ( // @[package.scala 93:22:@25641.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_23 ( // @[package.scala 93:22:@25650.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_194 RetimeWrapper_24 ( // @[package.scala 93:22:@25659.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_194 RetimeWrapper_25 ( // @[package.scala 93:22:@25668.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_196 RetimeWrapper_26 ( // @[package.scala 93:22:@25677.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_167 RetimeWrapper_27 ( // @[package.scala 93:22:@25686.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_194 RetimeWrapper_28 ( // @[package.scala 93:22:@25698.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_183 RetimeWrapper_29 ( // @[package.scala 93:22:@25719.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper RetimeWrapper_30 ( // @[package.scala 93:22:@25738.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_201 RetimeWrapper_31 ( // @[package.scala 93:22:@25750.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  x362_sum x421_sum_1 ( // @[Math.scala 150:24:@25759.4]
    .clock(x421_sum_1_clock),
    .reset(x421_sum_1_reset),
    .io_a(x421_sum_1_io_a),
    .io_b(x421_sum_1_io_b),
    .io_flow(x421_sum_1_io_flow),
    .io_result(x421_sum_1_io_result)
  );
  RetimeWrapper_167 RetimeWrapper_32 ( // @[package.scala 93:22:@25769.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_33 ( // @[package.scala 93:22:@25778.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_205 RetimeWrapper_34 ( // @[package.scala 93:22:@25787.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_194 RetimeWrapper_35 ( // @[package.scala 93:22:@25799.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  x362_sum x424_rdcol_1 ( // @[Math.scala 150:24:@25822.4]
    .clock(x424_rdcol_1_clock),
    .reset(x424_rdcol_1_reset),
    .io_a(x424_rdcol_1_io_a),
    .io_b(x424_rdcol_1_io_b),
    .io_flow(x424_rdcol_1_io_flow),
    .io_result(x424_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_36 ( // @[package.scala 93:22:@25842.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_37 ( // @[package.scala 93:22:@25874.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  x362_sum x430_sum_1 ( // @[Math.scala 150:24:@25883.4]
    .clock(x430_sum_1_clock),
    .reset(x430_sum_1_reset),
    .io_a(x430_sum_1_io_a),
    .io_b(x430_sum_1_io_b),
    .io_flow(x430_sum_1_io_flow),
    .io_result(x430_sum_1_io_result)
  );
  RetimeWrapper_167 RetimeWrapper_38 ( // @[package.scala 93:22:@25893.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_174 RetimeWrapper_39 ( // @[package.scala 93:22:@25902.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_40 ( // @[package.scala 93:22:@25911.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_194 RetimeWrapper_41 ( // @[package.scala 93:22:@25923.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  x362_sum x433_rdcol_1 ( // @[Math.scala 150:24:@25946.4]
    .clock(x433_rdcol_1_clock),
    .reset(x433_rdcol_1_reset),
    .io_a(x433_rdcol_1_io_a),
    .io_b(x433_rdcol_1_io_b),
    .io_flow(x433_rdcol_1_io_flow),
    .io_result(x433_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_42 ( // @[package.scala 93:22:@25966.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_43 ( // @[package.scala 93:22:@25998.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  x362_sum x439_sum_1 ( // @[Math.scala 150:24:@26007.4]
    .clock(x439_sum_1_clock),
    .reset(x439_sum_1_reset),
    .io_a(x439_sum_1_io_a),
    .io_b(x439_sum_1_io_b),
    .io_flow(x439_sum_1_io_flow),
    .io_result(x439_sum_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_44 ( // @[package.scala 93:22:@26017.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_167 RetimeWrapper_45 ( // @[package.scala 93:22:@26026.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_174 RetimeWrapper_46 ( // @[package.scala 93:22:@26035.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_194 RetimeWrapper_47 ( // @[package.scala 93:22:@26047.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  x577_sub x442_rdrow_1 ( // @[Math.scala 191:24:@26072.4]
    .clock(x442_rdrow_1_clock),
    .reset(x442_rdrow_1_reset),
    .io_a(x442_rdrow_1_io_a),
    .io_b(x442_rdrow_1_io_b),
    .io_flow(x442_rdrow_1_io_flow),
    .io_result(x442_rdrow_1_io_result)
  );
  RetimeWrapper RetimeWrapper_48 ( // @[package.scala 93:22:@26103.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_187 RetimeWrapper_49 ( // @[package.scala 93:22:@26137.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_188 RetimeWrapper_50 ( // @[package.scala 93:22:@26149.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  x577_sub x601_sub_1 ( // @[Math.scala 191:24:@26159.4]
    .clock(x601_sub_1_clock),
    .reset(x601_sub_1_reset),
    .io_a(x601_sub_1_io_a),
    .io_b(x601_sub_1_io_b),
    .io_flow(x601_sub_1_io_flow),
    .io_result(x601_sub_1_io_result)
  );
  RetimeWrapper_201 RetimeWrapper_51 ( // @[package.scala 93:22:@26169.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  x362_sum x450_sum_1 ( // @[Math.scala 150:24:@26178.4]
    .clock(x450_sum_1_clock),
    .reset(x450_sum_1_reset),
    .io_a(x450_sum_1_io_a),
    .io_b(x450_sum_1_io_b),
    .io_flow(x450_sum_1_io_flow),
    .io_result(x450_sum_1_io_result)
  );
  RetimeWrapper_174 RetimeWrapper_52 ( // @[package.scala 93:22:@26188.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_53 ( // @[package.scala 93:22:@26197.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_165 RetimeWrapper_54 ( // @[package.scala 93:22:@26206.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_194 RetimeWrapper_55 ( // @[package.scala 93:22:@26218.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper RetimeWrapper_56 ( // @[package.scala 93:22:@26239.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper RetimeWrapper_57 ( // @[package.scala 93:22:@26251.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_236 RetimeWrapper_58 ( // @[package.scala 93:22:@26263.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  x362_sum x455_sum_1 ( // @[Math.scala 150:24:@26272.4]
    .clock(x455_sum_1_clock),
    .reset(x455_sum_1_reset),
    .io_a(x455_sum_1_io_a),
    .io_b(x455_sum_1_io_b),
    .io_flow(x455_sum_1_io_flow),
    .io_result(x455_sum_1_io_result)
  );
  RetimeWrapper_165 RetimeWrapper_59 ( // @[package.scala 93:22:@26282.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_60 ( // @[package.scala 93:22:@26291.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_194 RetimeWrapper_61 ( // @[package.scala 93:22:@26303.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper RetimeWrapper_62 ( // @[package.scala 93:22:@26327.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_165 RetimeWrapper_63 ( // @[package.scala 93:22:@26339.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  x362_sum x460_sum_1 ( // @[Math.scala 150:24:@26348.4]
    .clock(x460_sum_1_clock),
    .reset(x460_sum_1_reset),
    .io_a(x460_sum_1_io_a),
    .io_b(x460_sum_1_io_b),
    .io_flow(x460_sum_1_io_flow),
    .io_result(x460_sum_1_io_result)
  );
  RetimeWrapper_165 RetimeWrapper_64 ( // @[package.scala 93:22:@26358.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_65 ( // @[package.scala 93:22:@26367.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_194 RetimeWrapper_66 ( // @[package.scala 93:22:@26379.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper RetimeWrapper_67 ( // @[package.scala 93:22:@26403.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_165 RetimeWrapper_68 ( // @[package.scala 93:22:@26415.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  x362_sum x465_sum_1 ( // @[Math.scala 150:24:@26424.4]
    .clock(x465_sum_1_clock),
    .reset(x465_sum_1_reset),
    .io_a(x465_sum_1_io_a),
    .io_b(x465_sum_1_io_b),
    .io_flow(x465_sum_1_io_flow),
    .io_result(x465_sum_1_io_result)
  );
  RetimeWrapper_165 RetimeWrapper_69 ( // @[package.scala 93:22:@26434.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_70 ( // @[package.scala 93:22:@26443.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_194 RetimeWrapper_71 ( // @[package.scala 93:22:@26455.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  x577_sub x468_rdrow_1 ( // @[Math.scala 191:24:@26480.4]
    .clock(x468_rdrow_1_clock),
    .reset(x468_rdrow_1_reset),
    .io_a(x468_rdrow_1_io_a),
    .io_b(x468_rdrow_1_io_b),
    .io_flow(x468_rdrow_1_io_flow),
    .io_result(x468_rdrow_1_io_result)
  );
  RetimeWrapper RetimeWrapper_72 ( // @[package.scala 93:22:@26511.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_187 RetimeWrapper_73 ( // @[package.scala 93:22:@26545.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_188 RetimeWrapper_74 ( // @[package.scala 93:22:@26557.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  x577_sub x606_sub_1 ( // @[Math.scala 191:24:@26567.4]
    .clock(x606_sub_1_clock),
    .reset(x606_sub_1_reset),
    .io_a(x606_sub_1_io_a),
    .io_b(x606_sub_1_io_b),
    .io_flow(x606_sub_1_io_flow),
    .io_result(x606_sub_1_io_result)
  );
  x362_sum x476_sum_1 ( // @[Math.scala 150:24:@26577.4]
    .clock(x476_sum_1_clock),
    .reset(x476_sum_1_reset),
    .io_a(x476_sum_1_io_a),
    .io_b(x476_sum_1_io_b),
    .io_flow(x476_sum_1_io_flow),
    .io_result(x476_sum_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_75 ( // @[package.scala 93:22:@26587.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_165 RetimeWrapper_76 ( // @[package.scala 93:22:@26596.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_174 RetimeWrapper_77 ( // @[package.scala 93:22:@26605.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_194 RetimeWrapper_78 ( // @[package.scala 93:22:@26617.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper RetimeWrapper_79 ( // @[package.scala 93:22:@26641.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  x362_sum x481_sum_1 ( // @[Math.scala 150:24:@26653.4]
    .clock(x481_sum_1_clock),
    .reset(x481_sum_1_reset),
    .io_a(x481_sum_1_io_a),
    .io_b(x481_sum_1_io_b),
    .io_flow(x481_sum_1_io_flow),
    .io_result(x481_sum_1_io_result)
  );
  RetimeWrapper_165 RetimeWrapper_80 ( // @[package.scala 93:22:@26663.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_81 ( // @[package.scala 93:22:@26672.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_194 RetimeWrapper_82 ( // @[package.scala 93:22:@26684.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper RetimeWrapper_83 ( // @[package.scala 93:22:@26708.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  x362_sum x486_sum_1 ( // @[Math.scala 150:24:@26720.4]
    .clock(x486_sum_1_clock),
    .reset(x486_sum_1_reset),
    .io_a(x486_sum_1_io_a),
    .io_b(x486_sum_1_io_b),
    .io_flow(x486_sum_1_io_flow),
    .io_result(x486_sum_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_84 ( // @[package.scala 93:22:@26730.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_165 RetimeWrapper_85 ( // @[package.scala 93:22:@26739.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_194 RetimeWrapper_86 ( // @[package.scala 93:22:@26751.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper RetimeWrapper_87 ( // @[package.scala 93:22:@26775.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  x362_sum x491_sum_1 ( // @[Math.scala 150:24:@26787.4]
    .clock(x491_sum_1_clock),
    .reset(x491_sum_1_reset),
    .io_a(x491_sum_1_io_a),
    .io_b(x491_sum_1_io_b),
    .io_flow(x491_sum_1_io_flow),
    .io_result(x491_sum_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_88 ( // @[package.scala 93:22:@26797.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_165 RetimeWrapper_89 ( // @[package.scala 93:22:@26806.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_194 RetimeWrapper_90 ( // @[package.scala 93:22:@26818.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  x499_x15 x499_x15_1 ( // @[Math.scala 150:24:@26864.4]
    .io_a(x499_x15_1_io_a),
    .io_b(x499_x15_1_io_b),
    .io_result(x499_x15_1_io_result)
  );
  x499_x15 x500_x16_1 ( // @[Math.scala 150:24:@26876.4]
    .io_a(x500_x16_1_io_a),
    .io_b(x500_x16_1_io_b),
    .io_result(x500_x16_1_io_result)
  );
  x499_x15 x501_x15_1 ( // @[Math.scala 150:24:@26886.4]
    .io_a(x501_x15_1_io_a),
    .io_b(x501_x15_1_io_b),
    .io_result(x501_x15_1_io_result)
  );
  x499_x15 x502_x16_1 ( // @[Math.scala 150:24:@26896.4]
    .io_a(x502_x16_1_io_a),
    .io_b(x502_x16_1_io_b),
    .io_result(x502_x16_1_io_result)
  );
  x499_x15 x503_x15_1 ( // @[Math.scala 150:24:@26906.4]
    .io_a(x503_x15_1_io_a),
    .io_b(x503_x15_1_io_b),
    .io_result(x503_x15_1_io_result)
  );
  x499_x15 x504_x16_1 ( // @[Math.scala 150:24:@26916.4]
    .io_a(x504_x16_1_io_a),
    .io_b(x504_x16_1_io_b),
    .io_result(x504_x16_1_io_result)
  );
  x499_x15 x505_x15_1 ( // @[Math.scala 150:24:@26926.4]
    .io_a(x505_x15_1_io_a),
    .io_b(x505_x15_1_io_b),
    .io_result(x505_x15_1_io_result)
  );
  x506_sum x506_sum_1 ( // @[Math.scala 150:24:@26936.4]
    .clock(x506_sum_1_clock),
    .reset(x506_sum_1_reset),
    .io_a(x506_sum_1_io_a),
    .io_b(x506_sum_1_io_b),
    .io_flow(x506_sum_1_io_flow),
    .io_result(x506_sum_1_io_result)
  );
  x499_x15 x513_x15_1 ( // @[Math.scala 150:24:@26978.4]
    .io_a(x513_x15_1_io_a),
    .io_b(x513_x15_1_io_b),
    .io_result(x513_x15_1_io_result)
  );
  x499_x15 x514_x16_1 ( // @[Math.scala 150:24:@26988.4]
    .io_a(x514_x16_1_io_a),
    .io_b(x514_x16_1_io_b),
    .io_result(x514_x16_1_io_result)
  );
  x499_x15 x515_x15_1 ( // @[Math.scala 150:24:@26998.4]
    .io_a(x515_x15_1_io_a),
    .io_b(x515_x15_1_io_b),
    .io_result(x515_x15_1_io_result)
  );
  x499_x15 x516_x16_1 ( // @[Math.scala 150:24:@27008.4]
    .io_a(x516_x16_1_io_a),
    .io_b(x516_x16_1_io_b),
    .io_result(x516_x16_1_io_result)
  );
  x499_x15 x517_x15_1 ( // @[Math.scala 150:24:@27018.4]
    .io_a(x517_x15_1_io_a),
    .io_b(x517_x15_1_io_b),
    .io_result(x517_x15_1_io_result)
  );
  x499_x15 x518_x16_1 ( // @[Math.scala 150:24:@27028.4]
    .io_a(x518_x16_1_io_a),
    .io_b(x518_x16_1_io_b),
    .io_result(x518_x16_1_io_result)
  );
  x499_x15 x519_x15_1 ( // @[Math.scala 150:24:@27038.4]
    .io_a(x519_x15_1_io_a),
    .io_b(x519_x15_1_io_b),
    .io_result(x519_x15_1_io_result)
  );
  x506_sum x520_sum_1 ( // @[Math.scala 150:24:@27048.4]
    .clock(x520_sum_1_clock),
    .reset(x520_sum_1_reset),
    .io_a(x520_sum_1_io_a),
    .io_b(x520_sum_1_io_b),
    .io_flow(x520_sum_1_io_flow),
    .io_result(x520_sum_1_io_result)
  );
  RetimeWrapper_280 RetimeWrapper_91 ( // @[package.scala 93:22:@27071.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_92 ( // @[package.scala 93:22:@27080.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_93 ( // @[package.scala 93:22:@27089.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_94 ( // @[package.scala 93:22:@27098.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  assign b381 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 62:18:@25056.4]
  assign b382 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 63:18:@25057.4]
  assign _T_205 = b381 & b382; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 67:30:@25059.4]
  assign _T_206 = _T_205 & io_sigsIn_datapathEn; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 67:37:@25060.4]
  assign _T_210 = io_in_x348_TID == 8'h0; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 69:76:@25065.4]
  assign _T_211 = _T_206 & _T_210; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 69:62:@25066.4]
  assign _T_213 = io_in_x348_TDEST == 8'h0; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 69:101:@25067.4]
  assign x612_x383_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@25076.4 package.scala 96:25:@25077.4]
  assign b379_number = __io_result; // @[Math.scala 712:22:@25041.4 Math.scala 713:14:@25042.4]
  assign _T_242 = $signed(b379_number); // @[Math.scala 499:52:@25185.4]
  assign x388 = $signed(32'sh1) == $signed(_T_242); // @[Math.scala 499:44:@25193.4]
  assign x389 = $signed(32'sh2) == $signed(_T_242); // @[Math.scala 499:44:@25200.4]
  assign x390 = $signed(32'sh3) == $signed(_T_242); // @[Math.scala 499:44:@25207.4]
  assign _T_289 = x388 ? 32'h1 : 32'h0; // @[Mux.scala 19:72:@25219.4]
  assign _T_291 = x389 ? 32'h2 : 32'h0; // @[Mux.scala 19:72:@25220.4]
  assign _T_293 = x390 ? 32'h3 : 32'h0; // @[Mux.scala 19:72:@25221.4]
  assign _T_295 = _T_289 | _T_291; // @[Mux.scala 19:72:@25223.4]
  assign x613_x391_D2_number = RetimeWrapper_1_io_out; // @[package.scala 96:25:@25236.4 package.scala 96:25:@25237.4]
  assign _T_310 = $signed(x613_x391_D2_number); // @[Math.scala 406:49:@25243.4]
  assign _T_312 = $signed(_T_310) & $signed(32'sh3); // @[Math.scala 406:56:@25245.4]
  assign _T_313 = $signed(_T_312); // @[Math.scala 406:56:@25246.4]
  assign b380_number = __1_io_result; // @[Math.scala 712:22:@25053.4 Math.scala 713:14:@25054.4]
  assign _T_322 = $signed(b380_number); // @[Math.scala 406:49:@25254.4]
  assign _T_324 = $signed(_T_322) & $signed(32'sh3); // @[Math.scala 406:56:@25256.4]
  assign _T_325 = $signed(_T_324); // @[Math.scala 406:56:@25257.4]
  assign _T_330 = x613_x391_D2_number[31]; // @[FixedPoint.scala 50:25:@25263.4]
  assign _T_334 = _T_330 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@25265.4]
  assign _T_335 = x613_x391_D2_number[31:2]; // @[FixedPoint.scala 18:52:@25266.4]
  assign x395_number = {_T_334,_T_335}; // @[Cat.scala 30:58:@25267.4]
  assign _GEN_0 = {{9'd0}, x395_number}; // @[Math.scala 450:32:@25272.4]
  assign _T_340 = _GEN_0 << 9; // @[Math.scala 450:32:@25272.4]
  assign _GEN_1 = {{5'd0}, x395_number}; // @[Math.scala 450:32:@25277.4]
  assign _T_344 = _GEN_1 << 5; // @[Math.scala 450:32:@25277.4]
  assign _T_351 = b380_number[31]; // @[FixedPoint.scala 50:25:@25292.4]
  assign _T_355 = _T_351 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@25294.4]
  assign _T_356 = b380_number[31:2]; // @[FixedPoint.scala 18:52:@25295.4]
  assign _T_383 = ~ io_sigsIn_break; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 127:101:@25372.4]
  assign _T_387 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@25380.4 package.scala 96:25:@25381.4]
  assign _T_389 = io_rr ? _T_387 : 1'h0; // @[implicits.scala 55:10:@25382.4]
  assign _T_390 = _T_383 & _T_389; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 127:118:@25383.4]
  assign _T_392 = _T_390 & _T_383; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 127:206:@25385.4]
  assign _T_393 = _T_392 & io_sigsIn_backpressure; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 127:225:@25386.4]
  assign x615_b381_D5 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@25324.4 package.scala 96:25:@25325.4]
  assign _T_394 = _T_393 & x615_b381_D5; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 127:251:@25387.4]
  assign x619_b382_D5 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@25360.4 package.scala 96:25:@25361.4]
  assign x400_rdcol_number = x400_rdcol_1_io_result; // @[Math.scala 154:22:@25404.4 Math.scala 155:14:@25405.4]
  assign _T_411 = $signed(x400_rdcol_number); // @[Math.scala 406:49:@25413.4]
  assign _T_413 = $signed(_T_411) & $signed(32'sh3); // @[Math.scala 406:56:@25415.4]
  assign _T_414 = $signed(_T_413); // @[Math.scala 406:56:@25416.4]
  assign _T_419 = x400_rdcol_number[31]; // @[FixedPoint.scala 50:25:@25422.4]
  assign _T_423 = _T_419 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@25424.4]
  assign _T_424 = x400_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@25425.4]
  assign _T_446 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@25483.4 package.scala 96:25:@25484.4]
  assign _T_448 = io_rr ? _T_446 : 1'h0; // @[implicits.scala 55:10:@25485.4]
  assign _T_449 = _T_383 & _T_448; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 150:118:@25486.4]
  assign _T_451 = _T_449 & _T_383; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 150:206:@25488.4]
  assign _T_452 = _T_451 & io_sigsIn_backpressure; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 150:225:@25489.4]
  assign _T_453 = _T_452 & x615_b381_D5; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 150:251:@25490.4]
  assign x625_b379_D8_number = RetimeWrapper_15_io_out; // @[package.scala 96:25:@25504.4 package.scala 96:25:@25505.4]
  assign _T_465 = $signed(x625_b379_D8_number); // @[Math.scala 406:49:@25511.4]
  assign _T_467 = $signed(_T_465) & $signed(32'sh3); // @[Math.scala 406:56:@25513.4]
  assign _T_468 = $signed(_T_467); // @[Math.scala 406:56:@25514.4]
  assign x590_number = $unsigned(_T_468); // @[implicits.scala 133:21:@25515.4]
  assign x408 = $signed(_T_465) < $signed(32'sh0); // @[Math.scala 465:44:@25523.4]
  assign x626_x400_rdcol_D8_number = RetimeWrapper_16_io_out; // @[package.scala 96:25:@25531.4 package.scala 96:25:@25532.4]
  assign _T_486 = $signed(x626_x400_rdcol_D8_number); // @[Math.scala 465:37:@25537.4]
  assign x409 = $signed(_T_486) < $signed(32'sh0); // @[Math.scala 465:44:@25539.4]
  assign x627_x408_D1 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@25547.4 package.scala 96:25:@25548.4]
  assign x628_x410_D1 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@25559.4 package.scala 96:25:@25560.4]
  assign _T_506 = $signed(x590_number); // @[Math.scala 406:49:@25569.4]
  assign _T_508 = $signed(_T_506) & $signed(32'sh3); // @[Math.scala 406:56:@25571.4]
  assign _T_509 = $signed(_T_508); // @[Math.scala 406:56:@25572.4]
  assign _T_516 = x590_number[31]; // @[FixedPoint.scala 50:25:@25580.4]
  assign _T_520 = _T_516 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@25582.4]
  assign _T_521 = x590_number[31:2]; // @[FixedPoint.scala 18:52:@25583.4]
  assign x413_number = {_T_520,_T_521}; // @[Cat.scala 30:58:@25584.4]
  assign _GEN_2 = {{9'd0}, x413_number}; // @[Math.scala 450:32:@25589.4]
  assign _GEN_3 = {{5'd0}, x413_number}; // @[Math.scala 450:32:@25601.4]
  assign _T_573 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@25703.4 package.scala 96:25:@25704.4]
  assign _T_575 = io_rr ? _T_573 : 1'h0; // @[implicits.scala 55:10:@25705.4]
  assign _T_576 = _T_383 & _T_575; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 208:194:@25706.4]
  assign x631_x411_D4 = RetimeWrapper_23_io_out; // @[package.scala 96:25:@25655.4 package.scala 96:25:@25656.4]
  assign _T_577 = _T_576 & x631_x411_D4; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 208:283:@25707.4]
  assign x632_b381_D14 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@25664.4 package.scala 96:25:@25665.4]
  assign _T_578 = _T_577 & x632_b381_D14; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 208:291:@25708.4]
  assign x633_b382_D14 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@25673.4 package.scala 96:25:@25674.4]
  assign x636_b380_D8_number = RetimeWrapper_29_io_out; // @[package.scala 96:25:@25724.4 package.scala 96:25:@25725.4]
  assign _T_589 = $signed(x636_b380_D8_number); // @[Math.scala 465:37:@25730.4]
  assign x418 = $signed(_T_589) < $signed(32'sh0); // @[Math.scala 465:44:@25732.4]
  assign x637_x419_D1 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@25743.4 package.scala 96:25:@25744.4]
  assign _T_625 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@25804.4 package.scala 96:25:@25805.4]
  assign _T_627 = io_rr ? _T_625 : 1'h0; // @[implicits.scala 55:10:@25806.4]
  assign _T_628 = _T_383 & _T_627; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 235:194:@25807.4]
  assign x640_x420_D5 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@25783.4 package.scala 96:25:@25784.4]
  assign _T_629 = _T_628 & x640_x420_D5; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 235:283:@25808.4]
  assign _T_630 = _T_629 & x632_b381_D14; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 235:291:@25809.4]
  assign x424_rdcol_number = x424_rdcol_1_io_result; // @[Math.scala 154:22:@25828.4 Math.scala 155:14:@25829.4]
  assign _T_645 = $signed(x424_rdcol_number); // @[Math.scala 465:37:@25834.4]
  assign x425 = $signed(_T_645) < $signed(32'sh0); // @[Math.scala 465:44:@25836.4]
  assign x642_x426_D1 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@25847.4 package.scala 96:25:@25848.4]
  assign _T_664 = $signed(_T_645) & $signed(32'sh3); // @[Math.scala 406:56:@25859.4]
  assign _T_665 = $signed(_T_664); // @[Math.scala 406:56:@25860.4]
  assign _T_670 = x424_rdcol_number[31]; // @[FixedPoint.scala 50:25:@25866.4]
  assign _T_674 = _T_670 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@25868.4]
  assign _T_675 = x424_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@25869.4]
  assign _T_703 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@25928.4 package.scala 96:25:@25929.4]
  assign _T_705 = io_rr ? _T_703 : 1'h0; // @[implicits.scala 55:10:@25930.4]
  assign _T_706 = _T_383 & _T_705; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 266:194:@25931.4]
  assign x646_x427_D4 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@25916.4 package.scala 96:25:@25917.4]
  assign _T_707 = _T_706 & x646_x427_D4; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 266:283:@25932.4]
  assign _T_708 = _T_707 & x632_b381_D14; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 266:291:@25933.4]
  assign x433_rdcol_number = x433_rdcol_1_io_result; // @[Math.scala 154:22:@25952.4 Math.scala 155:14:@25953.4]
  assign _T_723 = $signed(x433_rdcol_number); // @[Math.scala 465:37:@25958.4]
  assign x434 = $signed(_T_723) < $signed(32'sh0); // @[Math.scala 465:44:@25960.4]
  assign x647_x435_D1 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@25971.4 package.scala 96:25:@25972.4]
  assign _T_742 = $signed(_T_723) & $signed(32'sh3); // @[Math.scala 406:56:@25983.4]
  assign _T_743 = $signed(_T_742); // @[Math.scala 406:56:@25984.4]
  assign _T_748 = x433_rdcol_number[31]; // @[FixedPoint.scala 50:25:@25990.4]
  assign _T_752 = _T_748 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@25992.4]
  assign _T_753 = x433_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@25993.4]
  assign _T_781 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@26052.4 package.scala 96:25:@26053.4]
  assign _T_783 = io_rr ? _T_781 : 1'h0; // @[implicits.scala 55:10:@26054.4]
  assign _T_784 = _T_383 & _T_783; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 303:194:@26055.4]
  assign x649_x436_D4 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@26022.4 package.scala 96:25:@26023.4]
  assign _T_785 = _T_784 & x649_x436_D4; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 303:283:@26056.4]
  assign _T_786 = _T_785 & x632_b381_D14; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 303:291:@26057.4]
  assign x442_rdrow_number = x442_rdrow_1_io_result; // @[Math.scala 195:22:@26078.4 Math.scala 196:14:@26079.4]
  assign _T_805 = $signed(x442_rdrow_number); // @[Math.scala 406:49:@26085.4]
  assign _T_807 = $signed(_T_805) & $signed(32'sh3); // @[Math.scala 406:56:@26087.4]
  assign _T_808 = $signed(_T_807); // @[Math.scala 406:56:@26088.4]
  assign x597_number = $unsigned(_T_808); // @[implicits.scala 133:21:@26089.4]
  assign x444 = $signed(_T_805) < $signed(32'sh0); // @[Math.scala 465:44:@26097.4]
  assign x652_x445_D1 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@26108.4 package.scala 96:25:@26109.4]
  assign _T_832 = $signed(x597_number); // @[Math.scala 406:49:@26118.4]
  assign _T_834 = $signed(_T_832) & $signed(32'sh3); // @[Math.scala 406:56:@26120.4]
  assign _T_835 = $signed(_T_834); // @[Math.scala 406:56:@26121.4]
  assign _T_840 = x597_number[31]; // @[FixedPoint.scala 50:25:@26127.4]
  assign _T_844 = _T_840 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@26129.4]
  assign _T_845 = x597_number[31:2]; // @[FixedPoint.scala 18:52:@26130.4]
  assign x448_number = {_T_844,_T_845}; // @[Cat.scala 30:58:@26131.4]
  assign _GEN_4 = {{9'd0}, x448_number}; // @[Math.scala 450:32:@26136.4]
  assign _GEN_5 = {{5'd0}, x448_number}; // @[Math.scala 450:32:@26148.4]
  assign _T_888 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@26223.4 package.scala 96:25:@26224.4]
  assign _T_890 = io_rr ? _T_888 : 1'h0; // @[implicits.scala 55:10:@26225.4]
  assign _T_891 = _T_383 & _T_890; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 344:194:@26226.4]
  assign x655_x446_D4 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@26202.4 package.scala 96:25:@26203.4]
  assign _T_892 = _T_891 & x655_x446_D4; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 344:283:@26227.4]
  assign _T_893 = _T_892 & x632_b381_D14; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 344:291:@26228.4]
  assign x657_x418_D1 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@26244.4 package.scala 96:25:@26245.4]
  assign x658_x453_D1 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@26256.4 package.scala 96:25:@26257.4]
  assign _T_929 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@26308.4 package.scala 96:25:@26309.4]
  assign _T_931 = io_rr ? _T_929 : 1'h0; // @[implicits.scala 55:10:@26310.4]
  assign _T_932 = _T_383 & _T_931; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 367:194:@26311.4]
  assign x661_x454_D4 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@26296.4 package.scala 96:25:@26297.4]
  assign _T_933 = _T_932 & x661_x454_D4; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 367:283:@26312.4]
  assign _T_934 = _T_933 & x632_b381_D14; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 367:291:@26313.4]
  assign x662_x458_D1 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@26332.4 package.scala 96:25:@26333.4]
  assign _T_967 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@26384.4 package.scala 96:25:@26385.4]
  assign _T_969 = io_rr ? _T_967 : 1'h0; // @[implicits.scala 55:10:@26386.4]
  assign _T_970 = _T_383 & _T_969; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 388:194:@26387.4]
  assign x665_x459_D4 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@26372.4 package.scala 96:25:@26373.4]
  assign _T_971 = _T_970 & x665_x459_D4; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 388:283:@26388.4]
  assign _T_972 = _T_971 & x632_b381_D14; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 388:291:@26389.4]
  assign x666_x463_D1 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@26408.4 package.scala 96:25:@26409.4]
  assign _T_1005 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@26460.4 package.scala 96:25:@26461.4]
  assign _T_1007 = io_rr ? _T_1005 : 1'h0; // @[implicits.scala 55:10:@26462.4]
  assign _T_1008 = _T_383 & _T_1007; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 415:194:@26463.4]
  assign x669_x464_D4 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@26448.4 package.scala 96:25:@26449.4]
  assign _T_1009 = _T_1008 & x669_x464_D4; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 415:283:@26464.4]
  assign _T_1010 = _T_1009 & x632_b381_D14; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 415:326:@26465.4]
  assign x468_rdrow_number = x468_rdrow_1_io_result; // @[Math.scala 195:22:@26486.4 Math.scala 196:14:@26487.4]
  assign _T_1029 = $signed(x468_rdrow_number); // @[Math.scala 406:49:@26493.4]
  assign _T_1031 = $signed(_T_1029) & $signed(32'sh3); // @[Math.scala 406:56:@26495.4]
  assign _T_1032 = $signed(_T_1031); // @[Math.scala 406:56:@26496.4]
  assign x602_number = $unsigned(_T_1032); // @[implicits.scala 133:21:@26497.4]
  assign x470 = $signed(_T_1029) < $signed(32'sh0); // @[Math.scala 465:44:@26505.4]
  assign x670_x471_D1 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@26516.4 package.scala 96:25:@26517.4]
  assign _T_1056 = $signed(x602_number); // @[Math.scala 406:49:@26526.4]
  assign _T_1058 = $signed(_T_1056) & $signed(32'sh3); // @[Math.scala 406:56:@26528.4]
  assign _T_1059 = $signed(_T_1058); // @[Math.scala 406:56:@26529.4]
  assign _T_1064 = x602_number[31]; // @[FixedPoint.scala 50:25:@26535.4]
  assign _T_1068 = _T_1064 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@26537.4]
  assign _T_1069 = x602_number[31:2]; // @[FixedPoint.scala 18:52:@26538.4]
  assign x474_number = {_T_1068,_T_1069}; // @[Cat.scala 30:58:@26539.4]
  assign _GEN_6 = {{9'd0}, x474_number}; // @[Math.scala 450:32:@26544.4]
  assign _GEN_7 = {{5'd0}, x474_number}; // @[Math.scala 450:32:@26556.4]
  assign _T_1109 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@26622.4 package.scala 96:25:@26623.4]
  assign _T_1111 = io_rr ? _T_1109 : 1'h0; // @[implicits.scala 55:10:@26624.4]
  assign _T_1112 = _T_383 & _T_1111; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 454:194:@26625.4]
  assign x671_x472_D4 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@26592.4 package.scala 96:25:@26593.4]
  assign _T_1113 = _T_1112 & x671_x472_D4; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 454:283:@26626.4]
  assign _T_1114 = _T_1113 & x632_b381_D14; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 454:291:@26627.4]
  assign x674_x479_D1 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@26646.4 package.scala 96:25:@26647.4]
  assign _T_1144 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@26689.4 package.scala 96:25:@26690.4]
  assign _T_1146 = io_rr ? _T_1144 : 1'h0; // @[implicits.scala 55:10:@26691.4]
  assign _T_1147 = _T_383 & _T_1146; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 473:194:@26692.4]
  assign x676_x480_D4 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@26677.4 package.scala 96:25:@26678.4]
  assign _T_1148 = _T_1147 & x676_x480_D4; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 473:283:@26693.4]
  assign _T_1149 = _T_1148 & x632_b381_D14; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 473:291:@26694.4]
  assign x677_x484_D1 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@26713.4 package.scala 96:25:@26714.4]
  assign _T_1179 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@26756.4 package.scala 96:25:@26757.4]
  assign _T_1181 = io_rr ? _T_1179 : 1'h0; // @[implicits.scala 55:10:@26758.4]
  assign _T_1182 = _T_383 & _T_1181; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 492:194:@26759.4]
  assign x678_x485_D4 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@26735.4 package.scala 96:25:@26736.4]
  assign _T_1183 = _T_1182 & x678_x485_D4; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 492:283:@26760.4]
  assign _T_1184 = _T_1183 & x632_b381_D14; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 492:291:@26761.4]
  assign x680_x489_D1 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@26780.4 package.scala 96:25:@26781.4]
  assign _T_1214 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@26823.4 package.scala 96:25:@26824.4]
  assign _T_1216 = io_rr ? _T_1214 : 1'h0; // @[implicits.scala 55:10:@26825.4]
  assign _T_1217 = _T_383 & _T_1216; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 511:194:@26826.4]
  assign x681_x490_D4 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@26802.4 package.scala 96:25:@26803.4]
  assign _T_1218 = _T_1217 & x681_x490_D4; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 511:283:@26827.4]
  assign _T_1219 = _T_1218 & x632_b381_D14; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 511:291:@26828.4]
  assign x422_rd_0_number = x385_lb_0_io_rPort_11_output_0; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 231:29:@25795.4 sm_x526_inr_Foreach_SAMPLER_BOX.scala 235:338:@25816.4]
  assign _GEN_8 = {{1'd0}, x422_rd_0_number}; // @[Math.scala 450:32:@26840.4]
  assign _T_1225 = _GEN_8 << 1; // @[Math.scala 450:32:@26840.4]
  assign x451_rd_0_number = x385_lb_0_io_rPort_6_output_0; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 340:29:@26214.4 sm_x526_inr_Foreach_SAMPLER_BOX.scala 344:408:@26235.4]
  assign _GEN_9 = {{1'd0}, x451_rd_0_number}; // @[Math.scala 450:32:@26845.4]
  assign _T_1229 = _GEN_9 << 1; // @[Math.scala 450:32:@26845.4]
  assign x456_rd_0_number = x385_lb_0_io_rPort_4_output_0; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 363:29:@26299.4 sm_x526_inr_Foreach_SAMPLER_BOX.scala 367:408:@26320.4]
  assign _GEN_10 = {{2'd0}, x456_rd_0_number}; // @[Math.scala 450:32:@26850.4]
  assign _T_1233 = _GEN_10 << 2; // @[Math.scala 450:32:@26850.4]
  assign x461_rd_0_number = x385_lb_0_io_rPort_3_output_0; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 384:29:@26375.4 sm_x526_inr_Foreach_SAMPLER_BOX.scala 388:408:@26396.4]
  assign _GEN_11 = {{1'd0}, x461_rd_0_number}; // @[Math.scala 450:32:@26855.4]
  assign _T_1237 = _GEN_11 << 1; // @[Math.scala 450:32:@26855.4]
  assign x482_rd_0_number = x385_lb_0_io_rPort_10_output_0; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 469:29:@26680.4 sm_x526_inr_Foreach_SAMPLER_BOX.scala 473:408:@26701.4]
  assign _GEN_12 = {{1'd0}, x482_rd_0_number}; // @[Math.scala 450:32:@26860.4]
  assign _T_1241 = _GEN_12 << 1; // @[Math.scala 450:32:@26860.4]
  assign x506_sum_number = x506_sum_1_io_result; // @[Math.scala 154:22:@26942.4 Math.scala 155:14:@26943.4]
  assign _T_1276 = x506_sum_number[7:4]; // @[FixedPoint.scala 18:52:@26948.4]
  assign x507_number = {4'h0,_T_1276}; // @[Cat.scala 30:58:@26949.4]
  assign x431_rd_0_number = x385_lb_0_io_rPort_8_output_0; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 262:29:@25919.4 sm_x526_inr_Foreach_SAMPLER_BOX.scala 266:338:@25940.4]
  assign _GEN_13 = {{1'd0}, x431_rd_0_number}; // @[Math.scala 450:32:@26954.4]
  assign _T_1281 = _GEN_13 << 1; // @[Math.scala 450:32:@26954.4]
  assign _GEN_14 = {{1'd0}, x456_rd_0_number}; // @[Math.scala 450:32:@26959.4]
  assign _T_1285 = _GEN_14 << 1; // @[Math.scala 450:32:@26959.4]
  assign _GEN_15 = {{2'd0}, x461_rd_0_number}; // @[Math.scala 450:32:@26964.4]
  assign _T_1289 = _GEN_15 << 2; // @[Math.scala 450:32:@26964.4]
  assign x466_rd_0_number = x385_lb_0_io_rPort_5_output_0; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 411:29:@26451.4 sm_x526_inr_Foreach_SAMPLER_BOX.scala 415:443:@26472.4]
  assign _GEN_16 = {{1'd0}, x466_rd_0_number}; // @[Math.scala 450:32:@26969.4]
  assign _T_1293 = _GEN_16 << 1; // @[Math.scala 450:32:@26969.4]
  assign x487_rd_0_number = x385_lb_0_io_rPort_9_output_0; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 488:29:@26747.4 sm_x526_inr_Foreach_SAMPLER_BOX.scala 492:408:@26768.4]
  assign _GEN_17 = {{1'd0}, x487_rd_0_number}; // @[Math.scala 450:32:@26974.4]
  assign _T_1297 = _GEN_17 << 1; // @[Math.scala 450:32:@26974.4]
  assign x520_sum_number = x520_sum_1_io_result; // @[Math.scala 154:22:@27054.4 Math.scala 155:14:@27055.4]
  assign _T_1330 = x520_sum_number[7:4]; // @[FixedPoint.scala 18:52:@27060.4]
  assign x521_number = {4'h0,_T_1330}; // @[Cat.scala 30:58:@27061.4]
  assign _T_1353 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@27103.4 package.scala 96:25:@27104.4]
  assign _T_1355 = io_rr ? _T_1353 : 1'h0; // @[implicits.scala 55:10:@27105.4]
  assign x684_b381_D20 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@27094.4 package.scala 96:25:@27095.4]
  assign _T_1356 = _T_1355 & x684_b381_D20; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 587:117:@27106.4]
  assign x683_b382_D20 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@27085.4 package.scala 96:25:@27086.4]
  assign _T_1357 = _T_1356 & x683_b382_D20; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 587:123:@27107.4]
  assign x617_x398_sum_D1_number = RetimeWrapper_5_io_out; // @[package.scala 96:25:@25342.4 package.scala 96:25:@25343.4]
  assign x618_x584_D3_number = RetimeWrapper_6_io_out; // @[package.scala 96:25:@25351.4 package.scala 96:25:@25352.4]
  assign x620_x585_D5_number = RetimeWrapper_8_io_out; // @[package.scala 96:25:@25369.4 package.scala 96:25:@25370.4]
  assign x622_x404_sum_D1_number = RetimeWrapper_11_io_out; // @[package.scala 96:25:@25454.4 package.scala 96:25:@25455.4]
  assign x623_x589_D4_number = RetimeWrapper_12_io_out; // @[package.scala 96:25:@25463.4 package.scala 96:25:@25464.4]
  assign _T_528 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@25595.4 package.scala 96:25:@25596.4]
  assign _T_534 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@25607.4 package.scala 96:25:@25608.4]
  assign x630_x591_D6_number = RetimeWrapper_22_io_out; // @[package.scala 96:25:@25646.4 package.scala 96:25:@25647.4]
  assign x634_x589_D13_number = RetimeWrapper_26_io_out; // @[package.scala 96:25:@25682.4 package.scala 96:25:@25683.4]
  assign x635_x415_sum_D3_number = RetimeWrapper_27_io_out; // @[package.scala 96:25:@25691.4 package.scala 96:25:@25692.4]
  assign x639_x421_sum_D3_number = RetimeWrapper_32_io_out; // @[package.scala 96:25:@25774.4 package.scala 96:25:@25775.4]
  assign x641_x585_D14_number = RetimeWrapper_34_io_out; // @[package.scala 96:25:@25792.4 package.scala 96:25:@25793.4]
  assign x644_x430_sum_D3_number = RetimeWrapper_38_io_out; // @[package.scala 96:25:@25898.4 package.scala 96:25:@25899.4]
  assign x645_x595_D5_number = RetimeWrapper_39_io_out; // @[package.scala 96:25:@25907.4 package.scala 96:25:@25908.4]
  assign x650_x439_sum_D3_number = RetimeWrapper_45_io_out; // @[package.scala 96:25:@26031.4 package.scala 96:25:@26032.4]
  assign x651_x596_D5_number = RetimeWrapper_46_io_out; // @[package.scala 96:25:@26040.4 package.scala 96:25:@26041.4]
  assign _T_852 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@26142.4 package.scala 96:25:@26143.4]
  assign _T_858 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@26154.4 package.scala 96:25:@26155.4]
  assign x654_x598_D5_number = RetimeWrapper_52_io_out; // @[package.scala 96:25:@26193.4 package.scala 96:25:@26194.4]
  assign x656_x450_sum_D2_number = RetimeWrapper_54_io_out; // @[package.scala 96:25:@26211.4 package.scala 96:25:@26212.4]
  assign x660_x455_sum_D2_number = RetimeWrapper_59_io_out; // @[package.scala 96:25:@26287.4 package.scala 96:25:@26288.4]
  assign x664_x460_sum_D2_number = RetimeWrapper_64_io_out; // @[package.scala 96:25:@26363.4 package.scala 96:25:@26364.4]
  assign x668_x465_sum_D2_number = RetimeWrapper_69_io_out; // @[package.scala 96:25:@26439.4 package.scala 96:25:@26440.4]
  assign _T_1076 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@26550.4 package.scala 96:25:@26551.4]
  assign _T_1082 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@26562.4 package.scala 96:25:@26563.4]
  assign x672_x476_sum_D2_number = RetimeWrapper_76_io_out; // @[package.scala 96:25:@26601.4 package.scala 96:25:@26602.4]
  assign x673_x603_D5_number = RetimeWrapper_77_io_out; // @[package.scala 96:25:@26610.4 package.scala 96:25:@26611.4]
  assign x675_x481_sum_D2_number = RetimeWrapper_80_io_out; // @[package.scala 96:25:@26668.4 package.scala 96:25:@26669.4]
  assign x679_x486_sum_D2_number = RetimeWrapper_85_io_out; // @[package.scala 96:25:@26744.4 package.scala 96:25:@26745.4]
  assign x682_x491_sum_D2_number = RetimeWrapper_89_io_out; // @[package.scala 96:25:@26811.4 package.scala 96:25:@26812.4]
  assign io_in_x348_TREADY = _T_211 & _T_213; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 67:22:@25061.4 sm_x526_inr_Foreach_SAMPLER_BOX.scala 69:22:@25069.4]
  assign io_in_x349_TVALID = _T_1357 & io_sigsIn_backpressure; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 587:22:@27109.4]
  assign io_in_x349_TDATA = {{240'd0}, RetimeWrapper_91_io_out}; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 588:24:@27110.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@25039.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@25051.4]
  assign RetimeWrapper_clock = clock; // @[:@25072.4]
  assign RetimeWrapper_reset = reset; // @[:@25073.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25075.4]
  assign RetimeWrapper_io_in = io_in_x348_TDATA[15:0]; // @[package.scala 94:16:@25074.4]
  assign x385_lb_0_clock = clock; // @[:@25082.4]
  assign x385_lb_0_reset = reset; // @[:@25083.4]
  assign x385_lb_0_io_rPort_11_banks_1 = x641_x585_D14_number[2:0]; // @[MemInterfaceType.scala 106:58:@25812.4]
  assign x385_lb_0_io_rPort_11_banks_0 = x630_x591_D6_number[2:0]; // @[MemInterfaceType.scala 106:58:@25811.4]
  assign x385_lb_0_io_rPort_11_ofs_0 = x639_x421_sum_D3_number[8:0]; // @[MemInterfaceType.scala 107:54:@25813.4]
  assign x385_lb_0_io_rPort_11_en_0 = _T_630 & x633_b382_D14; // @[MemInterfaceType.scala 110:79:@25815.4]
  assign x385_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@25814.4]
  assign x385_lb_0_io_rPort_10_banks_1 = x641_x585_D14_number[2:0]; // @[MemInterfaceType.scala 106:58:@26697.4]
  assign x385_lb_0_io_rPort_10_banks_0 = x673_x603_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@26696.4]
  assign x385_lb_0_io_rPort_10_ofs_0 = x675_x481_sum_D2_number[8:0]; // @[MemInterfaceType.scala 107:54:@26698.4]
  assign x385_lb_0_io_rPort_10_en_0 = _T_1149 & x633_b382_D14; // @[MemInterfaceType.scala 110:79:@26700.4]
  assign x385_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26699.4]
  assign x385_lb_0_io_rPort_9_banks_1 = x645_x595_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@26764.4]
  assign x385_lb_0_io_rPort_9_banks_0 = x673_x603_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@26763.4]
  assign x385_lb_0_io_rPort_9_ofs_0 = x679_x486_sum_D2_number[8:0]; // @[MemInterfaceType.scala 107:54:@26765.4]
  assign x385_lb_0_io_rPort_9_en_0 = _T_1184 & x633_b382_D14; // @[MemInterfaceType.scala 110:79:@26767.4]
  assign x385_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26766.4]
  assign x385_lb_0_io_rPort_8_banks_1 = x645_x595_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@25936.4]
  assign x385_lb_0_io_rPort_8_banks_0 = x630_x591_D6_number[2:0]; // @[MemInterfaceType.scala 106:58:@25935.4]
  assign x385_lb_0_io_rPort_8_ofs_0 = x644_x430_sum_D3_number[8:0]; // @[MemInterfaceType.scala 107:54:@25937.4]
  assign x385_lb_0_io_rPort_8_en_0 = _T_708 & x633_b382_D14; // @[MemInterfaceType.scala 110:79:@25939.4]
  assign x385_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@25938.4]
  assign x385_lb_0_io_rPort_7_banks_1 = x634_x589_D13_number[2:0]; // @[MemInterfaceType.scala 106:58:@26630.4]
  assign x385_lb_0_io_rPort_7_banks_0 = x673_x603_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@26629.4]
  assign x385_lb_0_io_rPort_7_ofs_0 = x672_x476_sum_D2_number[8:0]; // @[MemInterfaceType.scala 107:54:@26631.4]
  assign x385_lb_0_io_rPort_7_en_0 = _T_1114 & x633_b382_D14; // @[MemInterfaceType.scala 110:79:@26633.4]
  assign x385_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26632.4]
  assign x385_lb_0_io_rPort_6_banks_1 = x634_x589_D13_number[2:0]; // @[MemInterfaceType.scala 106:58:@26231.4]
  assign x385_lb_0_io_rPort_6_banks_0 = x654_x598_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@26230.4]
  assign x385_lb_0_io_rPort_6_ofs_0 = x656_x450_sum_D2_number[8:0]; // @[MemInterfaceType.scala 107:54:@26232.4]
  assign x385_lb_0_io_rPort_6_en_0 = _T_893 & x633_b382_D14; // @[MemInterfaceType.scala 110:79:@26234.4]
  assign x385_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26233.4]
  assign x385_lb_0_io_rPort_5_banks_1 = x651_x596_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@26468.4]
  assign x385_lb_0_io_rPort_5_banks_0 = x654_x598_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@26467.4]
  assign x385_lb_0_io_rPort_5_ofs_0 = x668_x465_sum_D2_number[8:0]; // @[MemInterfaceType.scala 107:54:@26469.4]
  assign x385_lb_0_io_rPort_5_en_0 = _T_1010 & x633_b382_D14; // @[MemInterfaceType.scala 110:79:@26471.4]
  assign x385_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26470.4]
  assign x385_lb_0_io_rPort_4_banks_1 = x641_x585_D14_number[2:0]; // @[MemInterfaceType.scala 106:58:@26316.4]
  assign x385_lb_0_io_rPort_4_banks_0 = x654_x598_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@26315.4]
  assign x385_lb_0_io_rPort_4_ofs_0 = x660_x455_sum_D2_number[8:0]; // @[MemInterfaceType.scala 107:54:@26317.4]
  assign x385_lb_0_io_rPort_4_en_0 = _T_934 & x633_b382_D14; // @[MemInterfaceType.scala 110:79:@26319.4]
  assign x385_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26318.4]
  assign x385_lb_0_io_rPort_3_banks_1 = x645_x595_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@26392.4]
  assign x385_lb_0_io_rPort_3_banks_0 = x654_x598_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@26391.4]
  assign x385_lb_0_io_rPort_3_ofs_0 = x664_x460_sum_D2_number[8:0]; // @[MemInterfaceType.scala 107:54:@26393.4]
  assign x385_lb_0_io_rPort_3_en_0 = _T_972 & x633_b382_D14; // @[MemInterfaceType.scala 110:79:@26395.4]
  assign x385_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26394.4]
  assign x385_lb_0_io_rPort_2_banks_1 = x651_x596_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@26831.4]
  assign x385_lb_0_io_rPort_2_banks_0 = x673_x603_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@26830.4]
  assign x385_lb_0_io_rPort_2_ofs_0 = x682_x491_sum_D2_number[8:0]; // @[MemInterfaceType.scala 107:54:@26832.4]
  assign x385_lb_0_io_rPort_2_en_0 = _T_1219 & x633_b382_D14; // @[MemInterfaceType.scala 110:79:@26834.4]
  assign x385_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26833.4]
  assign x385_lb_0_io_rPort_1_banks_1 = x634_x589_D13_number[2:0]; // @[MemInterfaceType.scala 106:58:@25711.4]
  assign x385_lb_0_io_rPort_1_banks_0 = x630_x591_D6_number[2:0]; // @[MemInterfaceType.scala 106:58:@25710.4]
  assign x385_lb_0_io_rPort_1_ofs_0 = x635_x415_sum_D3_number[8:0]; // @[MemInterfaceType.scala 107:54:@25712.4]
  assign x385_lb_0_io_rPort_1_en_0 = _T_578 & x633_b382_D14; // @[MemInterfaceType.scala 110:79:@25714.4]
  assign x385_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@25713.4]
  assign x385_lb_0_io_rPort_0_banks_1 = x651_x596_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@26060.4]
  assign x385_lb_0_io_rPort_0_banks_0 = x630_x591_D6_number[2:0]; // @[MemInterfaceType.scala 106:58:@26059.4]
  assign x385_lb_0_io_rPort_0_ofs_0 = x650_x439_sum_D3_number[8:0]; // @[MemInterfaceType.scala 107:54:@26061.4]
  assign x385_lb_0_io_rPort_0_en_0 = _T_786 & x633_b382_D14; // @[MemInterfaceType.scala 110:79:@26063.4]
  assign x385_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26062.4]
  assign x385_lb_0_io_wPort_1_banks_1 = x623_x589_D4_number[2:0]; // @[MemInterfaceType.scala 88:58:@25493.4]
  assign x385_lb_0_io_wPort_1_banks_0 = x618_x584_D3_number[2:0]; // @[MemInterfaceType.scala 88:58:@25492.4]
  assign x385_lb_0_io_wPort_1_ofs_0 = x622_x404_sum_D1_number[8:0]; // @[MemInterfaceType.scala 89:54:@25494.4]
  assign x385_lb_0_io_wPort_1_data_0 = RetimeWrapper_13_io_out; // @[MemInterfaceType.scala 90:56:@25495.4]
  assign x385_lb_0_io_wPort_1_en_0 = _T_453 & x619_b382_D5; // @[MemInterfaceType.scala 93:57:@25497.4]
  assign x385_lb_0_io_wPort_0_banks_1 = x620_x585_D5_number[2:0]; // @[MemInterfaceType.scala 88:58:@25390.4]
  assign x385_lb_0_io_wPort_0_banks_0 = x618_x584_D3_number[2:0]; // @[MemInterfaceType.scala 88:58:@25389.4]
  assign x385_lb_0_io_wPort_0_ofs_0 = x617_x398_sum_D1_number[8:0]; // @[MemInterfaceType.scala 89:54:@25391.4]
  assign x385_lb_0_io_wPort_0_data_0 = RetimeWrapper_4_io_out; // @[MemInterfaceType.scala 90:56:@25392.4]
  assign x385_lb_0_io_wPort_0_en_0 = _T_394 & x619_b382_D5; // @[MemInterfaceType.scala 93:57:@25394.4]
  assign RetimeWrapper_1_clock = clock; // @[:@25232.4]
  assign RetimeWrapper_1_reset = reset; // @[:@25233.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25235.4]
  assign RetimeWrapper_1_io_in = _T_295 | _T_293; // @[package.scala 94:16:@25234.4]
  assign x588_sub_1_clock = clock; // @[:@25282.4]
  assign x588_sub_1_reset = reset; // @[:@25283.4]
  assign x588_sub_1_io_a = _T_340[31:0]; // @[Math.scala 192:17:@25284.4]
  assign x588_sub_1_io_b = _T_344[31:0]; // @[Math.scala 193:17:@25285.4]
  assign x588_sub_1_io_flow = io_in_x349_TREADY; // @[Math.scala 194:20:@25286.4]
  assign RetimeWrapper_2_clock = clock; // @[:@25301.4]
  assign RetimeWrapper_2_reset = reset; // @[:@25302.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25304.4]
  assign RetimeWrapper_2_io_in = {_T_355,_T_356}; // @[package.scala 94:16:@25303.4]
  assign x398_sum_1_clock = clock; // @[:@25310.4]
  assign x398_sum_1_reset = reset; // @[:@25311.4]
  assign x398_sum_1_io_a = x588_sub_1_io_result; // @[Math.scala 151:17:@25312.4]
  assign x398_sum_1_io_b = RetimeWrapper_2_io_out; // @[Math.scala 152:17:@25313.4]
  assign x398_sum_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@25314.4]
  assign RetimeWrapper_3_clock = clock; // @[:@25320.4]
  assign RetimeWrapper_3_reset = reset; // @[:@25321.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25323.4]
  assign RetimeWrapper_3_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@25322.4]
  assign RetimeWrapper_4_clock = clock; // @[:@25329.4]
  assign RetimeWrapper_4_reset = reset; // @[:@25330.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25332.4]
  assign RetimeWrapper_4_io_in = x612_x383_D1_0_number[7:0]; // @[package.scala 94:16:@25331.4]
  assign RetimeWrapper_5_clock = clock; // @[:@25338.4]
  assign RetimeWrapper_5_reset = reset; // @[:@25339.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25341.4]
  assign RetimeWrapper_5_io_in = x398_sum_1_io_result; // @[package.scala 94:16:@25340.4]
  assign RetimeWrapper_6_clock = clock; // @[:@25347.4]
  assign RetimeWrapper_6_reset = reset; // @[:@25348.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25350.4]
  assign RetimeWrapper_6_io_in = $unsigned(_T_313); // @[package.scala 94:16:@25349.4]
  assign RetimeWrapper_7_clock = clock; // @[:@25356.4]
  assign RetimeWrapper_7_reset = reset; // @[:@25357.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25359.4]
  assign RetimeWrapper_7_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@25358.4]
  assign RetimeWrapper_8_clock = clock; // @[:@25365.4]
  assign RetimeWrapper_8_reset = reset; // @[:@25366.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25368.4]
  assign RetimeWrapper_8_io_in = $unsigned(_T_325); // @[package.scala 94:16:@25367.4]
  assign RetimeWrapper_9_clock = clock; // @[:@25376.4]
  assign RetimeWrapper_9_reset = reset; // @[:@25377.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25379.4]
  assign RetimeWrapper_9_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@25378.4]
  assign x400_rdcol_1_clock = clock; // @[:@25399.4]
  assign x400_rdcol_1_reset = reset; // @[:@25400.4]
  assign x400_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@25401.4]
  assign x400_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@25402.4]
  assign x400_rdcol_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@25403.4]
  assign RetimeWrapper_10_clock = clock; // @[:@25431.4]
  assign RetimeWrapper_10_reset = reset; // @[:@25432.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25434.4]
  assign RetimeWrapper_10_io_in = {_T_423,_T_424}; // @[package.scala 94:16:@25433.4]
  assign x404_sum_1_clock = clock; // @[:@25440.4]
  assign x404_sum_1_reset = reset; // @[:@25441.4]
  assign x404_sum_1_io_a = x588_sub_1_io_result; // @[Math.scala 151:17:@25442.4]
  assign x404_sum_1_io_b = RetimeWrapper_10_io_out; // @[Math.scala 152:17:@25443.4]
  assign x404_sum_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@25444.4]
  assign RetimeWrapper_11_clock = clock; // @[:@25450.4]
  assign RetimeWrapper_11_reset = reset; // @[:@25451.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25453.4]
  assign RetimeWrapper_11_io_in = x404_sum_1_io_result; // @[package.scala 94:16:@25452.4]
  assign RetimeWrapper_12_clock = clock; // @[:@25459.4]
  assign RetimeWrapper_12_reset = reset; // @[:@25460.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25462.4]
  assign RetimeWrapper_12_io_in = $unsigned(_T_414); // @[package.scala 94:16:@25461.4]
  assign RetimeWrapper_13_clock = clock; // @[:@25468.4]
  assign RetimeWrapper_13_reset = reset; // @[:@25469.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25471.4]
  assign RetimeWrapper_13_io_in = x612_x383_D1_0_number[15:8]; // @[package.scala 94:16:@25470.4]
  assign RetimeWrapper_14_clock = clock; // @[:@25479.4]
  assign RetimeWrapper_14_reset = reset; // @[:@25480.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25482.4]
  assign RetimeWrapper_14_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@25481.4]
  assign RetimeWrapper_15_clock = clock; // @[:@25500.4]
  assign RetimeWrapper_15_reset = reset; // @[:@25501.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25503.4]
  assign RetimeWrapper_15_io_in = __io_result; // @[package.scala 94:16:@25502.4]
  assign RetimeWrapper_16_clock = clock; // @[:@25527.4]
  assign RetimeWrapper_16_reset = reset; // @[:@25528.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25530.4]
  assign RetimeWrapper_16_io_in = x400_rdcol_1_io_result; // @[package.scala 94:16:@25529.4]
  assign RetimeWrapper_17_clock = clock; // @[:@25543.4]
  assign RetimeWrapper_17_reset = reset; // @[:@25544.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25546.4]
  assign RetimeWrapper_17_io_in = $signed(_T_465) < $signed(32'sh0); // @[package.scala 94:16:@25545.4]
  assign RetimeWrapper_18_clock = clock; // @[:@25555.4]
  assign RetimeWrapper_18_reset = reset; // @[:@25556.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25558.4]
  assign RetimeWrapper_18_io_in = x627_x408_D1 | x409; // @[package.scala 94:16:@25557.4]
  assign RetimeWrapper_19_clock = clock; // @[:@25591.4]
  assign RetimeWrapper_19_reset = reset; // @[:@25592.4]
  assign RetimeWrapper_19_io_flow = io_in_x349_TREADY; // @[package.scala 95:18:@25594.4]
  assign RetimeWrapper_19_io_in = _GEN_2 << 9; // @[package.scala 94:16:@25593.4]
  assign RetimeWrapper_20_clock = clock; // @[:@25603.4]
  assign RetimeWrapper_20_reset = reset; // @[:@25604.4]
  assign RetimeWrapper_20_io_flow = io_in_x349_TREADY; // @[package.scala 95:18:@25606.4]
  assign RetimeWrapper_20_io_in = _GEN_3 << 5; // @[package.scala 94:16:@25605.4]
  assign x594_sub_1_clock = clock; // @[:@25613.4]
  assign x594_sub_1_reset = reset; // @[:@25614.4]
  assign x594_sub_1_io_a = _T_528[31:0]; // @[Math.scala 192:17:@25615.4]
  assign x594_sub_1_io_b = _T_534[31:0]; // @[Math.scala 193:17:@25616.4]
  assign x594_sub_1_io_flow = io_in_x349_TREADY; // @[Math.scala 194:20:@25617.4]
  assign RetimeWrapper_21_clock = clock; // @[:@25623.4]
  assign RetimeWrapper_21_reset = reset; // @[:@25624.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25626.4]
  assign RetimeWrapper_21_io_in = {_T_423,_T_424}; // @[package.scala 94:16:@25625.4]
  assign x415_sum_1_clock = clock; // @[:@25632.4]
  assign x415_sum_1_reset = reset; // @[:@25633.4]
  assign x415_sum_1_io_a = x594_sub_1_io_result; // @[Math.scala 151:17:@25634.4]
  assign x415_sum_1_io_b = RetimeWrapper_21_io_out; // @[Math.scala 152:17:@25635.4]
  assign x415_sum_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@25636.4]
  assign RetimeWrapper_22_clock = clock; // @[:@25642.4]
  assign RetimeWrapper_22_reset = reset; // @[:@25643.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25645.4]
  assign RetimeWrapper_22_io_in = $unsigned(_T_509); // @[package.scala 94:16:@25644.4]
  assign RetimeWrapper_23_clock = clock; // @[:@25651.4]
  assign RetimeWrapper_23_reset = reset; // @[:@25652.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25654.4]
  assign RetimeWrapper_23_io_in = ~ x628_x410_D1; // @[package.scala 94:16:@25653.4]
  assign RetimeWrapper_24_clock = clock; // @[:@25660.4]
  assign RetimeWrapper_24_reset = reset; // @[:@25661.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25663.4]
  assign RetimeWrapper_24_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@25662.4]
  assign RetimeWrapper_25_clock = clock; // @[:@25669.4]
  assign RetimeWrapper_25_reset = reset; // @[:@25670.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25672.4]
  assign RetimeWrapper_25_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@25671.4]
  assign RetimeWrapper_26_clock = clock; // @[:@25678.4]
  assign RetimeWrapper_26_reset = reset; // @[:@25679.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25681.4]
  assign RetimeWrapper_26_io_in = $unsigned(_T_414); // @[package.scala 94:16:@25680.4]
  assign RetimeWrapper_27_clock = clock; // @[:@25687.4]
  assign RetimeWrapper_27_reset = reset; // @[:@25688.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25690.4]
  assign RetimeWrapper_27_io_in = x415_sum_1_io_result; // @[package.scala 94:16:@25689.4]
  assign RetimeWrapper_28_clock = clock; // @[:@25699.4]
  assign RetimeWrapper_28_reset = reset; // @[:@25700.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25702.4]
  assign RetimeWrapper_28_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@25701.4]
  assign RetimeWrapper_29_clock = clock; // @[:@25720.4]
  assign RetimeWrapper_29_reset = reset; // @[:@25721.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25723.4]
  assign RetimeWrapper_29_io_in = __1_io_result; // @[package.scala 94:16:@25722.4]
  assign RetimeWrapper_30_clock = clock; // @[:@25739.4]
  assign RetimeWrapper_30_reset = reset; // @[:@25740.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25742.4]
  assign RetimeWrapper_30_io_in = x408 | x418; // @[package.scala 94:16:@25741.4]
  assign RetimeWrapper_31_clock = clock; // @[:@25751.4]
  assign RetimeWrapper_31_reset = reset; // @[:@25752.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25754.4]
  assign RetimeWrapper_31_io_in = {_T_355,_T_356}; // @[package.scala 94:16:@25753.4]
  assign x421_sum_1_clock = clock; // @[:@25760.4]
  assign x421_sum_1_reset = reset; // @[:@25761.4]
  assign x421_sum_1_io_a = x594_sub_1_io_result; // @[Math.scala 151:17:@25762.4]
  assign x421_sum_1_io_b = RetimeWrapper_31_io_out; // @[Math.scala 152:17:@25763.4]
  assign x421_sum_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@25764.4]
  assign RetimeWrapper_32_clock = clock; // @[:@25770.4]
  assign RetimeWrapper_32_reset = reset; // @[:@25771.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25773.4]
  assign RetimeWrapper_32_io_in = x421_sum_1_io_result; // @[package.scala 94:16:@25772.4]
  assign RetimeWrapper_33_clock = clock; // @[:@25779.4]
  assign RetimeWrapper_33_reset = reset; // @[:@25780.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25782.4]
  assign RetimeWrapper_33_io_in = ~ x637_x419_D1; // @[package.scala 94:16:@25781.4]
  assign RetimeWrapper_34_clock = clock; // @[:@25788.4]
  assign RetimeWrapper_34_reset = reset; // @[:@25789.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25791.4]
  assign RetimeWrapper_34_io_in = $unsigned(_T_325); // @[package.scala 94:16:@25790.4]
  assign RetimeWrapper_35_clock = clock; // @[:@25800.4]
  assign RetimeWrapper_35_reset = reset; // @[:@25801.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25803.4]
  assign RetimeWrapper_35_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@25802.4]
  assign x424_rdcol_1_clock = clock; // @[:@25823.4]
  assign x424_rdcol_1_reset = reset; // @[:@25824.4]
  assign x424_rdcol_1_io_a = RetimeWrapper_29_io_out; // @[Math.scala 151:17:@25825.4]
  assign x424_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@25826.4]
  assign x424_rdcol_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@25827.4]
  assign RetimeWrapper_36_clock = clock; // @[:@25843.4]
  assign RetimeWrapper_36_reset = reset; // @[:@25844.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25846.4]
  assign RetimeWrapper_36_io_in = x627_x408_D1 | x425; // @[package.scala 94:16:@25845.4]
  assign RetimeWrapper_37_clock = clock; // @[:@25875.4]
  assign RetimeWrapper_37_reset = reset; // @[:@25876.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25878.4]
  assign RetimeWrapper_37_io_in = {_T_674,_T_675}; // @[package.scala 94:16:@25877.4]
  assign x430_sum_1_clock = clock; // @[:@25884.4]
  assign x430_sum_1_reset = reset; // @[:@25885.4]
  assign x430_sum_1_io_a = x594_sub_1_io_result; // @[Math.scala 151:17:@25886.4]
  assign x430_sum_1_io_b = RetimeWrapper_37_io_out; // @[Math.scala 152:17:@25887.4]
  assign x430_sum_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@25888.4]
  assign RetimeWrapper_38_clock = clock; // @[:@25894.4]
  assign RetimeWrapper_38_reset = reset; // @[:@25895.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25897.4]
  assign RetimeWrapper_38_io_in = x430_sum_1_io_result; // @[package.scala 94:16:@25896.4]
  assign RetimeWrapper_39_clock = clock; // @[:@25903.4]
  assign RetimeWrapper_39_reset = reset; // @[:@25904.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25906.4]
  assign RetimeWrapper_39_io_in = $unsigned(_T_665); // @[package.scala 94:16:@25905.4]
  assign RetimeWrapper_40_clock = clock; // @[:@25912.4]
  assign RetimeWrapper_40_reset = reset; // @[:@25913.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25915.4]
  assign RetimeWrapper_40_io_in = ~ x642_x426_D1; // @[package.scala 94:16:@25914.4]
  assign RetimeWrapper_41_clock = clock; // @[:@25924.4]
  assign RetimeWrapper_41_reset = reset; // @[:@25925.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25927.4]
  assign RetimeWrapper_41_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@25926.4]
  assign x433_rdcol_1_clock = clock; // @[:@25947.4]
  assign x433_rdcol_1_reset = reset; // @[:@25948.4]
  assign x433_rdcol_1_io_a = RetimeWrapper_29_io_out; // @[Math.scala 151:17:@25949.4]
  assign x433_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@25950.4]
  assign x433_rdcol_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@25951.4]
  assign RetimeWrapper_42_clock = clock; // @[:@25967.4]
  assign RetimeWrapper_42_reset = reset; // @[:@25968.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25970.4]
  assign RetimeWrapper_42_io_in = x627_x408_D1 | x434; // @[package.scala 94:16:@25969.4]
  assign RetimeWrapper_43_clock = clock; // @[:@25999.4]
  assign RetimeWrapper_43_reset = reset; // @[:@26000.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26002.4]
  assign RetimeWrapper_43_io_in = {_T_752,_T_753}; // @[package.scala 94:16:@26001.4]
  assign x439_sum_1_clock = clock; // @[:@26008.4]
  assign x439_sum_1_reset = reset; // @[:@26009.4]
  assign x439_sum_1_io_a = x594_sub_1_io_result; // @[Math.scala 151:17:@26010.4]
  assign x439_sum_1_io_b = RetimeWrapper_43_io_out; // @[Math.scala 152:17:@26011.4]
  assign x439_sum_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@26012.4]
  assign RetimeWrapper_44_clock = clock; // @[:@26018.4]
  assign RetimeWrapper_44_reset = reset; // @[:@26019.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26021.4]
  assign RetimeWrapper_44_io_in = ~ x647_x435_D1; // @[package.scala 94:16:@26020.4]
  assign RetimeWrapper_45_clock = clock; // @[:@26027.4]
  assign RetimeWrapper_45_reset = reset; // @[:@26028.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26030.4]
  assign RetimeWrapper_45_io_in = x439_sum_1_io_result; // @[package.scala 94:16:@26029.4]
  assign RetimeWrapper_46_clock = clock; // @[:@26036.4]
  assign RetimeWrapper_46_reset = reset; // @[:@26037.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26039.4]
  assign RetimeWrapper_46_io_in = $unsigned(_T_743); // @[package.scala 94:16:@26038.4]
  assign RetimeWrapper_47_clock = clock; // @[:@26048.4]
  assign RetimeWrapper_47_reset = reset; // @[:@26049.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26051.4]
  assign RetimeWrapper_47_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26050.4]
  assign x442_rdrow_1_clock = clock; // @[:@26073.4]
  assign x442_rdrow_1_reset = reset; // @[:@26074.4]
  assign x442_rdrow_1_io_a = RetimeWrapper_15_io_out; // @[Math.scala 192:17:@26075.4]
  assign x442_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@26076.4]
  assign x442_rdrow_1_io_flow = io_in_x349_TREADY; // @[Math.scala 194:20:@26077.4]
  assign RetimeWrapper_48_clock = clock; // @[:@26104.4]
  assign RetimeWrapper_48_reset = reset; // @[:@26105.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26107.4]
  assign RetimeWrapper_48_io_in = x444 | x409; // @[package.scala 94:16:@26106.4]
  assign RetimeWrapper_49_clock = clock; // @[:@26138.4]
  assign RetimeWrapper_49_reset = reset; // @[:@26139.4]
  assign RetimeWrapper_49_io_flow = io_in_x349_TREADY; // @[package.scala 95:18:@26141.4]
  assign RetimeWrapper_49_io_in = _GEN_4 << 9; // @[package.scala 94:16:@26140.4]
  assign RetimeWrapper_50_clock = clock; // @[:@26150.4]
  assign RetimeWrapper_50_reset = reset; // @[:@26151.4]
  assign RetimeWrapper_50_io_flow = io_in_x349_TREADY; // @[package.scala 95:18:@26153.4]
  assign RetimeWrapper_50_io_in = _GEN_5 << 5; // @[package.scala 94:16:@26152.4]
  assign x601_sub_1_clock = clock; // @[:@26160.4]
  assign x601_sub_1_reset = reset; // @[:@26161.4]
  assign x601_sub_1_io_a = _T_852[31:0]; // @[Math.scala 192:17:@26162.4]
  assign x601_sub_1_io_b = _T_858[31:0]; // @[Math.scala 193:17:@26163.4]
  assign x601_sub_1_io_flow = io_in_x349_TREADY; // @[Math.scala 194:20:@26164.4]
  assign RetimeWrapper_51_clock = clock; // @[:@26170.4]
  assign RetimeWrapper_51_reset = reset; // @[:@26171.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26173.4]
  assign RetimeWrapper_51_io_in = {_T_423,_T_424}; // @[package.scala 94:16:@26172.4]
  assign x450_sum_1_clock = clock; // @[:@26179.4]
  assign x450_sum_1_reset = reset; // @[:@26180.4]
  assign x450_sum_1_io_a = x601_sub_1_io_result; // @[Math.scala 151:17:@26181.4]
  assign x450_sum_1_io_b = RetimeWrapper_51_io_out; // @[Math.scala 152:17:@26182.4]
  assign x450_sum_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@26183.4]
  assign RetimeWrapper_52_clock = clock; // @[:@26189.4]
  assign RetimeWrapper_52_reset = reset; // @[:@26190.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26192.4]
  assign RetimeWrapper_52_io_in = $unsigned(_T_835); // @[package.scala 94:16:@26191.4]
  assign RetimeWrapper_53_clock = clock; // @[:@26198.4]
  assign RetimeWrapper_53_reset = reset; // @[:@26199.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26201.4]
  assign RetimeWrapper_53_io_in = ~ x652_x445_D1; // @[package.scala 94:16:@26200.4]
  assign RetimeWrapper_54_clock = clock; // @[:@26207.4]
  assign RetimeWrapper_54_reset = reset; // @[:@26208.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26210.4]
  assign RetimeWrapper_54_io_in = x450_sum_1_io_result; // @[package.scala 94:16:@26209.4]
  assign RetimeWrapper_55_clock = clock; // @[:@26219.4]
  assign RetimeWrapper_55_reset = reset; // @[:@26220.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26222.4]
  assign RetimeWrapper_55_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26221.4]
  assign RetimeWrapper_56_clock = clock; // @[:@26240.4]
  assign RetimeWrapper_56_reset = reset; // @[:@26241.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26243.4]
  assign RetimeWrapper_56_io_in = $signed(_T_589) < $signed(32'sh0); // @[package.scala 94:16:@26242.4]
  assign RetimeWrapper_57_clock = clock; // @[:@26252.4]
  assign RetimeWrapper_57_reset = reset; // @[:@26253.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26255.4]
  assign RetimeWrapper_57_io_in = x444 | x657_x418_D1; // @[package.scala 94:16:@26254.4]
  assign RetimeWrapper_58_clock = clock; // @[:@26264.4]
  assign RetimeWrapper_58_reset = reset; // @[:@26265.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26267.4]
  assign RetimeWrapper_58_io_in = {_T_355,_T_356}; // @[package.scala 94:16:@26266.4]
  assign x455_sum_1_clock = clock; // @[:@26273.4]
  assign x455_sum_1_reset = reset; // @[:@26274.4]
  assign x455_sum_1_io_a = x601_sub_1_io_result; // @[Math.scala 151:17:@26275.4]
  assign x455_sum_1_io_b = RetimeWrapper_58_io_out; // @[Math.scala 152:17:@26276.4]
  assign x455_sum_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@26277.4]
  assign RetimeWrapper_59_clock = clock; // @[:@26283.4]
  assign RetimeWrapper_59_reset = reset; // @[:@26284.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26286.4]
  assign RetimeWrapper_59_io_in = x455_sum_1_io_result; // @[package.scala 94:16:@26285.4]
  assign RetimeWrapper_60_clock = clock; // @[:@26292.4]
  assign RetimeWrapper_60_reset = reset; // @[:@26293.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26295.4]
  assign RetimeWrapper_60_io_in = ~ x658_x453_D1; // @[package.scala 94:16:@26294.4]
  assign RetimeWrapper_61_clock = clock; // @[:@26304.4]
  assign RetimeWrapper_61_reset = reset; // @[:@26305.4]
  assign RetimeWrapper_61_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26307.4]
  assign RetimeWrapper_61_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26306.4]
  assign RetimeWrapper_62_clock = clock; // @[:@26328.4]
  assign RetimeWrapper_62_reset = reset; // @[:@26329.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26331.4]
  assign RetimeWrapper_62_io_in = x444 | x425; // @[package.scala 94:16:@26330.4]
  assign RetimeWrapper_63_clock = clock; // @[:@26340.4]
  assign RetimeWrapper_63_reset = reset; // @[:@26341.4]
  assign RetimeWrapper_63_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26343.4]
  assign RetimeWrapper_63_io_in = {_T_674,_T_675}; // @[package.scala 94:16:@26342.4]
  assign x460_sum_1_clock = clock; // @[:@26349.4]
  assign x460_sum_1_reset = reset; // @[:@26350.4]
  assign x460_sum_1_io_a = x601_sub_1_io_result; // @[Math.scala 151:17:@26351.4]
  assign x460_sum_1_io_b = RetimeWrapper_63_io_out; // @[Math.scala 152:17:@26352.4]
  assign x460_sum_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@26353.4]
  assign RetimeWrapper_64_clock = clock; // @[:@26359.4]
  assign RetimeWrapper_64_reset = reset; // @[:@26360.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26362.4]
  assign RetimeWrapper_64_io_in = x460_sum_1_io_result; // @[package.scala 94:16:@26361.4]
  assign RetimeWrapper_65_clock = clock; // @[:@26368.4]
  assign RetimeWrapper_65_reset = reset; // @[:@26369.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26371.4]
  assign RetimeWrapper_65_io_in = ~ x662_x458_D1; // @[package.scala 94:16:@26370.4]
  assign RetimeWrapper_66_clock = clock; // @[:@26380.4]
  assign RetimeWrapper_66_reset = reset; // @[:@26381.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26383.4]
  assign RetimeWrapper_66_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26382.4]
  assign RetimeWrapper_67_clock = clock; // @[:@26404.4]
  assign RetimeWrapper_67_reset = reset; // @[:@26405.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26407.4]
  assign RetimeWrapper_67_io_in = x444 | x434; // @[package.scala 94:16:@26406.4]
  assign RetimeWrapper_68_clock = clock; // @[:@26416.4]
  assign RetimeWrapper_68_reset = reset; // @[:@26417.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26419.4]
  assign RetimeWrapper_68_io_in = {_T_752,_T_753}; // @[package.scala 94:16:@26418.4]
  assign x465_sum_1_clock = clock; // @[:@26425.4]
  assign x465_sum_1_reset = reset; // @[:@26426.4]
  assign x465_sum_1_io_a = x601_sub_1_io_result; // @[Math.scala 151:17:@26427.4]
  assign x465_sum_1_io_b = RetimeWrapper_68_io_out; // @[Math.scala 152:17:@26428.4]
  assign x465_sum_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@26429.4]
  assign RetimeWrapper_69_clock = clock; // @[:@26435.4]
  assign RetimeWrapper_69_reset = reset; // @[:@26436.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26438.4]
  assign RetimeWrapper_69_io_in = x465_sum_1_io_result; // @[package.scala 94:16:@26437.4]
  assign RetimeWrapper_70_clock = clock; // @[:@26444.4]
  assign RetimeWrapper_70_reset = reset; // @[:@26445.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26447.4]
  assign RetimeWrapper_70_io_in = ~ x666_x463_D1; // @[package.scala 94:16:@26446.4]
  assign RetimeWrapper_71_clock = clock; // @[:@26456.4]
  assign RetimeWrapper_71_reset = reset; // @[:@26457.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26459.4]
  assign RetimeWrapper_71_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26458.4]
  assign x468_rdrow_1_clock = clock; // @[:@26481.4]
  assign x468_rdrow_1_reset = reset; // @[:@26482.4]
  assign x468_rdrow_1_io_a = RetimeWrapper_15_io_out; // @[Math.scala 192:17:@26483.4]
  assign x468_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@26484.4]
  assign x468_rdrow_1_io_flow = io_in_x349_TREADY; // @[Math.scala 194:20:@26485.4]
  assign RetimeWrapper_72_clock = clock; // @[:@26512.4]
  assign RetimeWrapper_72_reset = reset; // @[:@26513.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26515.4]
  assign RetimeWrapper_72_io_in = x470 | x409; // @[package.scala 94:16:@26514.4]
  assign RetimeWrapper_73_clock = clock; // @[:@26546.4]
  assign RetimeWrapper_73_reset = reset; // @[:@26547.4]
  assign RetimeWrapper_73_io_flow = io_in_x349_TREADY; // @[package.scala 95:18:@26549.4]
  assign RetimeWrapper_73_io_in = _GEN_6 << 9; // @[package.scala 94:16:@26548.4]
  assign RetimeWrapper_74_clock = clock; // @[:@26558.4]
  assign RetimeWrapper_74_reset = reset; // @[:@26559.4]
  assign RetimeWrapper_74_io_flow = io_in_x349_TREADY; // @[package.scala 95:18:@26561.4]
  assign RetimeWrapper_74_io_in = _GEN_7 << 5; // @[package.scala 94:16:@26560.4]
  assign x606_sub_1_clock = clock; // @[:@26568.4]
  assign x606_sub_1_reset = reset; // @[:@26569.4]
  assign x606_sub_1_io_a = _T_1076[31:0]; // @[Math.scala 192:17:@26570.4]
  assign x606_sub_1_io_b = _T_1082[31:0]; // @[Math.scala 193:17:@26571.4]
  assign x606_sub_1_io_flow = io_in_x349_TREADY; // @[Math.scala 194:20:@26572.4]
  assign x476_sum_1_clock = clock; // @[:@26578.4]
  assign x476_sum_1_reset = reset; // @[:@26579.4]
  assign x476_sum_1_io_a = x606_sub_1_io_result; // @[Math.scala 151:17:@26580.4]
  assign x476_sum_1_io_b = RetimeWrapper_51_io_out; // @[Math.scala 152:17:@26581.4]
  assign x476_sum_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@26582.4]
  assign RetimeWrapper_75_clock = clock; // @[:@26588.4]
  assign RetimeWrapper_75_reset = reset; // @[:@26589.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26591.4]
  assign RetimeWrapper_75_io_in = ~ x670_x471_D1; // @[package.scala 94:16:@26590.4]
  assign RetimeWrapper_76_clock = clock; // @[:@26597.4]
  assign RetimeWrapper_76_reset = reset; // @[:@26598.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26600.4]
  assign RetimeWrapper_76_io_in = x476_sum_1_io_result; // @[package.scala 94:16:@26599.4]
  assign RetimeWrapper_77_clock = clock; // @[:@26606.4]
  assign RetimeWrapper_77_reset = reset; // @[:@26607.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26609.4]
  assign RetimeWrapper_77_io_in = $unsigned(_T_1059); // @[package.scala 94:16:@26608.4]
  assign RetimeWrapper_78_clock = clock; // @[:@26618.4]
  assign RetimeWrapper_78_reset = reset; // @[:@26619.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26621.4]
  assign RetimeWrapper_78_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26620.4]
  assign RetimeWrapper_79_clock = clock; // @[:@26642.4]
  assign RetimeWrapper_79_reset = reset; // @[:@26643.4]
  assign RetimeWrapper_79_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26645.4]
  assign RetimeWrapper_79_io_in = x470 | x657_x418_D1; // @[package.scala 94:16:@26644.4]
  assign x481_sum_1_clock = clock; // @[:@26654.4]
  assign x481_sum_1_reset = reset; // @[:@26655.4]
  assign x481_sum_1_io_a = x606_sub_1_io_result; // @[Math.scala 151:17:@26656.4]
  assign x481_sum_1_io_b = RetimeWrapper_58_io_out; // @[Math.scala 152:17:@26657.4]
  assign x481_sum_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@26658.4]
  assign RetimeWrapper_80_clock = clock; // @[:@26664.4]
  assign RetimeWrapper_80_reset = reset; // @[:@26665.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26667.4]
  assign RetimeWrapper_80_io_in = x481_sum_1_io_result; // @[package.scala 94:16:@26666.4]
  assign RetimeWrapper_81_clock = clock; // @[:@26673.4]
  assign RetimeWrapper_81_reset = reset; // @[:@26674.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26676.4]
  assign RetimeWrapper_81_io_in = ~ x674_x479_D1; // @[package.scala 94:16:@26675.4]
  assign RetimeWrapper_82_clock = clock; // @[:@26685.4]
  assign RetimeWrapper_82_reset = reset; // @[:@26686.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26688.4]
  assign RetimeWrapper_82_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26687.4]
  assign RetimeWrapper_83_clock = clock; // @[:@26709.4]
  assign RetimeWrapper_83_reset = reset; // @[:@26710.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26712.4]
  assign RetimeWrapper_83_io_in = x470 | x425; // @[package.scala 94:16:@26711.4]
  assign x486_sum_1_clock = clock; // @[:@26721.4]
  assign x486_sum_1_reset = reset; // @[:@26722.4]
  assign x486_sum_1_io_a = x606_sub_1_io_result; // @[Math.scala 151:17:@26723.4]
  assign x486_sum_1_io_b = RetimeWrapper_63_io_out; // @[Math.scala 152:17:@26724.4]
  assign x486_sum_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@26725.4]
  assign RetimeWrapper_84_clock = clock; // @[:@26731.4]
  assign RetimeWrapper_84_reset = reset; // @[:@26732.4]
  assign RetimeWrapper_84_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26734.4]
  assign RetimeWrapper_84_io_in = ~ x677_x484_D1; // @[package.scala 94:16:@26733.4]
  assign RetimeWrapper_85_clock = clock; // @[:@26740.4]
  assign RetimeWrapper_85_reset = reset; // @[:@26741.4]
  assign RetimeWrapper_85_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26743.4]
  assign RetimeWrapper_85_io_in = x486_sum_1_io_result; // @[package.scala 94:16:@26742.4]
  assign RetimeWrapper_86_clock = clock; // @[:@26752.4]
  assign RetimeWrapper_86_reset = reset; // @[:@26753.4]
  assign RetimeWrapper_86_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26755.4]
  assign RetimeWrapper_86_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26754.4]
  assign RetimeWrapper_87_clock = clock; // @[:@26776.4]
  assign RetimeWrapper_87_reset = reset; // @[:@26777.4]
  assign RetimeWrapper_87_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26779.4]
  assign RetimeWrapper_87_io_in = x470 | x434; // @[package.scala 94:16:@26778.4]
  assign x491_sum_1_clock = clock; // @[:@26788.4]
  assign x491_sum_1_reset = reset; // @[:@26789.4]
  assign x491_sum_1_io_a = x606_sub_1_io_result; // @[Math.scala 151:17:@26790.4]
  assign x491_sum_1_io_b = RetimeWrapper_68_io_out; // @[Math.scala 152:17:@26791.4]
  assign x491_sum_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@26792.4]
  assign RetimeWrapper_88_clock = clock; // @[:@26798.4]
  assign RetimeWrapper_88_reset = reset; // @[:@26799.4]
  assign RetimeWrapper_88_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26801.4]
  assign RetimeWrapper_88_io_in = ~ x680_x489_D1; // @[package.scala 94:16:@26800.4]
  assign RetimeWrapper_89_clock = clock; // @[:@26807.4]
  assign RetimeWrapper_89_reset = reset; // @[:@26808.4]
  assign RetimeWrapper_89_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26810.4]
  assign RetimeWrapper_89_io_in = x491_sum_1_io_result; // @[package.scala 94:16:@26809.4]
  assign RetimeWrapper_90_clock = clock; // @[:@26819.4]
  assign RetimeWrapper_90_reset = reset; // @[:@26820.4]
  assign RetimeWrapper_90_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26822.4]
  assign RetimeWrapper_90_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26821.4]
  assign x499_x15_1_io_a = x385_lb_0_io_rPort_1_output_0; // @[Math.scala 151:17:@26867.4]
  assign x499_x15_1_io_b = _T_1225[7:0]; // @[Math.scala 152:17:@26868.4]
  assign x500_x16_1_io_a = x385_lb_0_io_rPort_8_output_0; // @[Math.scala 151:17:@26879.4]
  assign x500_x16_1_io_b = _T_1229[7:0]; // @[Math.scala 152:17:@26880.4]
  assign x501_x15_1_io_a = _T_1233[7:0]; // @[Math.scala 151:17:@26889.4]
  assign x501_x15_1_io_b = _T_1237[7:0]; // @[Math.scala 152:17:@26890.4]
  assign x502_x16_1_io_a = x385_lb_0_io_rPort_7_output_0; // @[Math.scala 151:17:@26899.4]
  assign x502_x16_1_io_b = _T_1241[7:0]; // @[Math.scala 152:17:@26900.4]
  assign x503_x15_1_io_a = x499_x15_1_io_result; // @[Math.scala 151:17:@26909.4]
  assign x503_x15_1_io_b = x500_x16_1_io_result; // @[Math.scala 152:17:@26910.4]
  assign x504_x16_1_io_a = x501_x15_1_io_result; // @[Math.scala 151:17:@26919.4]
  assign x504_x16_1_io_b = x502_x16_1_io_result; // @[Math.scala 152:17:@26920.4]
  assign x505_x15_1_io_a = x503_x15_1_io_result; // @[Math.scala 151:17:@26929.4]
  assign x505_x15_1_io_b = x504_x16_1_io_result; // @[Math.scala 152:17:@26930.4]
  assign x506_sum_1_clock = clock; // @[:@26937.4]
  assign x506_sum_1_reset = reset; // @[:@26938.4]
  assign x506_sum_1_io_a = x505_x15_1_io_result; // @[Math.scala 151:17:@26939.4]
  assign x506_sum_1_io_b = x385_lb_0_io_rPort_9_output_0; // @[Math.scala 152:17:@26940.4]
  assign x506_sum_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@26941.4]
  assign x513_x15_1_io_a = x385_lb_0_io_rPort_11_output_0; // @[Math.scala 151:17:@26981.4]
  assign x513_x15_1_io_b = _T_1281[7:0]; // @[Math.scala 152:17:@26982.4]
  assign x514_x16_1_io_a = x385_lb_0_io_rPort_0_output_0; // @[Math.scala 151:17:@26991.4]
  assign x514_x16_1_io_b = _T_1285[7:0]; // @[Math.scala 152:17:@26992.4]
  assign x515_x15_1_io_a = _T_1289[7:0]; // @[Math.scala 151:17:@27001.4]
  assign x515_x15_1_io_b = _T_1293[7:0]; // @[Math.scala 152:17:@27002.4]
  assign x516_x16_1_io_a = x385_lb_0_io_rPort_10_output_0; // @[Math.scala 151:17:@27011.4]
  assign x516_x16_1_io_b = _T_1297[7:0]; // @[Math.scala 152:17:@27012.4]
  assign x517_x15_1_io_a = x513_x15_1_io_result; // @[Math.scala 151:17:@27021.4]
  assign x517_x15_1_io_b = x514_x16_1_io_result; // @[Math.scala 152:17:@27022.4]
  assign x518_x16_1_io_a = x515_x15_1_io_result; // @[Math.scala 151:17:@27031.4]
  assign x518_x16_1_io_b = x516_x16_1_io_result; // @[Math.scala 152:17:@27032.4]
  assign x519_x15_1_io_a = x517_x15_1_io_result; // @[Math.scala 151:17:@27041.4]
  assign x519_x15_1_io_b = x518_x16_1_io_result; // @[Math.scala 152:17:@27042.4]
  assign x520_sum_1_clock = clock; // @[:@27049.4]
  assign x520_sum_1_reset = reset; // @[:@27050.4]
  assign x520_sum_1_io_a = x519_x15_1_io_result; // @[Math.scala 151:17:@27051.4]
  assign x520_sum_1_io_b = x385_lb_0_io_rPort_2_output_0; // @[Math.scala 152:17:@27052.4]
  assign x520_sum_1_io_flow = io_in_x349_TREADY; // @[Math.scala 153:20:@27053.4]
  assign RetimeWrapper_91_clock = clock; // @[:@27072.4]
  assign RetimeWrapper_91_reset = reset; // @[:@27073.4]
  assign RetimeWrapper_91_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27075.4]
  assign RetimeWrapper_91_io_in = {x507_number,x521_number}; // @[package.scala 94:16:@27074.4]
  assign RetimeWrapper_92_clock = clock; // @[:@27081.4]
  assign RetimeWrapper_92_reset = reset; // @[:@27082.4]
  assign RetimeWrapper_92_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27084.4]
  assign RetimeWrapper_92_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@27083.4]
  assign RetimeWrapper_93_clock = clock; // @[:@27090.4]
  assign RetimeWrapper_93_reset = reset; // @[:@27091.4]
  assign RetimeWrapper_93_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27093.4]
  assign RetimeWrapper_93_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@27092.4]
  assign RetimeWrapper_94_clock = clock; // @[:@27099.4]
  assign RetimeWrapper_94_reset = reset; // @[:@27100.4]
  assign RetimeWrapper_94_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27102.4]
  assign RetimeWrapper_94_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27101.4]
endmodule
module x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1( // @[:@27120.2]
  input          clock, // @[:@27121.4]
  input          reset, // @[:@27122.4]
  input          io_in_x348_TVALID, // @[:@27123.4]
  output         io_in_x348_TREADY, // @[:@27123.4]
  input  [255:0] io_in_x348_TDATA, // @[:@27123.4]
  input  [7:0]   io_in_x348_TID, // @[:@27123.4]
  input  [7:0]   io_in_x348_TDEST, // @[:@27123.4]
  output         io_in_x349_TVALID, // @[:@27123.4]
  input          io_in_x349_TREADY, // @[:@27123.4]
  output [255:0] io_in_x349_TDATA, // @[:@27123.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@27123.4]
  input          io_sigsIn_smChildAcks_0, // @[:@27123.4]
  output         io_sigsOut_smDoneIn_0, // @[:@27123.4]
  input          io_rr // @[:@27123.4]
);
  wire  x378_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@27157.4]
  wire  x378_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@27157.4]
  wire  x378_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@27157.4]
  wire  x378_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@27157.4]
  wire [12:0] x378_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@27157.4]
  wire [12:0] x378_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@27157.4]
  wire  x378_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@27157.4]
  wire  x378_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@27157.4]
  wire  x378_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@27157.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 32:18:@27217.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 32:18:@27217.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 32:18:@27217.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 32:18:@27217.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 32:18:@27217.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 32:18:@27217.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 32:18:@27217.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 32:18:@27217.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 32:18:@27217.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 32:18:@27217.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 32:18:@27217.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 32:18:@27217.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@27245.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@27245.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@27245.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@27245.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@27245.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@27287.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@27287.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@27287.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@27287.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@27287.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@27295.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@27295.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@27295.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@27295.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@27295.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 600:24:@27329.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 600:24:@27329.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x348_TREADY; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 600:24:@27329.4]
  wire [255:0] x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x348_TDATA; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 600:24:@27329.4]
  wire [7:0] x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x348_TID; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 600:24:@27329.4]
  wire [7:0] x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x348_TDEST; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 600:24:@27329.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x349_TVALID; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 600:24:@27329.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x349_TREADY; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 600:24:@27329.4]
  wire [255:0] x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x349_TDATA; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 600:24:@27329.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 600:24:@27329.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 600:24:@27329.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 600:24:@27329.4]
  wire [31:0] x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 600:24:@27329.4]
  wire [31:0] x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 600:24:@27329.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 600:24:@27329.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 600:24:@27329.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 600:24:@27329.4]
  wire  _T_240; // @[package.scala 96:25:@27250.4 package.scala 96:25:@27251.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x527_outr_UnitPipe.scala 69:66:@27256.4]
  wire  _T_253; // @[package.scala 96:25:@27292.4 package.scala 96:25:@27293.4]
  wire  _T_259; // @[package.scala 96:25:@27300.4 package.scala 96:25:@27301.4]
  wire  _T_262; // @[SpatialBlocks.scala 138:93:@27303.4]
  wire  x526_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@27304.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:36:@27312.4]
  wire  _T_265; // @[SpatialBlocks.scala 157:78:@27313.4]
  wire  _T_272; // @[SpatialBlocks.scala 159:58:@27325.4]
  x356_ctrchain x378_ctrchain ( // @[SpatialBlocks.scala 37:22:@27157.4]
    .clock(x378_ctrchain_clock),
    .reset(x378_ctrchain_reset),
    .io_input_reset(x378_ctrchain_io_input_reset),
    .io_input_enable(x378_ctrchain_io_input_enable),
    .io_output_counts_1(x378_ctrchain_io_output_counts_1),
    .io_output_counts_0(x378_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x378_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x378_ctrchain_io_output_oobs_1),
    .io_output_done(x378_ctrchain_io_output_done)
  );
  x526_inr_Foreach_SAMPLER_BOX_sm x526_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 32:18:@27217.4]
    .clock(x526_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x526_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x526_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x526_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x526_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x526_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x526_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x526_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x526_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x526_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x526_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x526_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@27245.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@27287.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@27295.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1 x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 600:24:@27329.4]
    .clock(x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x348_TREADY(x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x348_TREADY),
    .io_in_x348_TDATA(x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x348_TDATA),
    .io_in_x348_TID(x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x348_TID),
    .io_in_x348_TDEST(x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x348_TDEST),
    .io_in_x349_TVALID(x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x349_TVALID),
    .io_in_x349_TREADY(x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x349_TREADY),
    .io_in_x349_TDATA(x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x349_TDATA),
    .io_sigsIn_backpressure(x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_240 = RetimeWrapper_io_out; // @[package.scala 96:25:@27250.4 package.scala 96:25:@27251.4]
  assign x526_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x348_TVALID | x526_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x527_outr_UnitPipe.scala 69:66:@27256.4]
  assign _T_253 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@27292.4 package.scala 96:25:@27293.4]
  assign _T_259 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@27300.4 package.scala 96:25:@27301.4]
  assign _T_262 = ~ _T_259; // @[SpatialBlocks.scala 138:93:@27303.4]
  assign x526_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_253 & _T_262; // @[SpatialBlocks.scala 138:90:@27304.4]
  assign _T_264 = x526_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@27312.4]
  assign _T_265 = ~ x526_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@27313.4]
  assign _T_272 = x526_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@27325.4]
  assign io_in_x348_TREADY = x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x348_TREADY; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 48:23:@27387.4]
  assign io_in_x349_TVALID = x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x349_TVALID; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 49:23:@27397.4]
  assign io_in_x349_TDATA = x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x349_TDATA; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 49:23:@27395.4]
  assign io_sigsOut_smDoneIn_0 = x526_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@27310.4]
  assign x378_ctrchain_clock = clock; // @[:@27158.4]
  assign x378_ctrchain_reset = reset; // @[:@27159.4]
  assign x378_ctrchain_io_input_reset = x526_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@27328.4]
  assign x378_ctrchain_io_input_enable = _T_272 & x526_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@27280.4 SpatialBlocks.scala 159:42:@27327.4]
  assign x526_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@27218.4]
  assign x526_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@27219.4]
  assign x526_inr_Foreach_SAMPLER_BOX_sm_io_enable = x526_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x526_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@27307.4]
  assign x526_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_240 : 1'h0; // @[sm_x527_outr_UnitPipe.scala 67:50:@27253.4]
  assign x526_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@27309.4]
  assign x526_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x349_TREADY | x526_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@27281.4]
  assign x526_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x527_outr_UnitPipe.scala 71:48:@27259.4]
  assign RetimeWrapper_clock = clock; // @[:@27246.4]
  assign RetimeWrapper_reset = reset; // @[:@27247.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@27249.4]
  assign RetimeWrapper_io_in = x378_ctrchain_io_output_done; // @[package.scala 94:16:@27248.4]
  assign RetimeWrapper_1_clock = clock; // @[:@27288.4]
  assign RetimeWrapper_1_reset = reset; // @[:@27289.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@27291.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@27290.4]
  assign RetimeWrapper_2_clock = clock; // @[:@27296.4]
  assign RetimeWrapper_2_reset = reset; // @[:@27297.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@27299.4]
  assign RetimeWrapper_2_io_in = x526_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@27298.4]
  assign x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@27330.4]
  assign x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@27331.4]
  assign x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x348_TDATA = io_in_x348_TDATA; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 48:23:@27386.4]
  assign x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x348_TID = io_in_x348_TID; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 48:23:@27382.4]
  assign x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x348_TDEST = io_in_x348_TDEST; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 48:23:@27381.4]
  assign x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x349_TREADY = io_in_x349_TREADY; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 49:23:@27396.4]
  assign x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x349_TREADY | x526_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 605:22:@27414.4]
  assign x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_264 & _T_265; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 605:22:@27412.4]
  assign x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x526_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 605:22:@27410.4]
  assign x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x378_ctrchain_io_output_counts_1[12]}},x378_ctrchain_io_output_counts_1}; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 605:22:@27405.4]
  assign x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x378_ctrchain_io_output_counts_0[12]}},x378_ctrchain_io_output_counts_0}; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 605:22:@27404.4]
  assign x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x378_ctrchain_io_output_oobs_0; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 605:22:@27402.4]
  assign x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x378_ctrchain_io_output_oobs_1; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 605:22:@27403.4]
  assign x526_inr_Foreach_SAMPLER_BOX_kernelx526_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x526_inr_Foreach_SAMPLER_BOX.scala 604:18:@27398.4]
endmodule
module x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1( // @[:@27428.2]
  input          clock, // @[:@27429.4]
  input          reset, // @[:@27430.4]
  input          io_in_x348_TVALID, // @[:@27431.4]
  output         io_in_x348_TREADY, // @[:@27431.4]
  input  [255:0] io_in_x348_TDATA, // @[:@27431.4]
  input  [7:0]   io_in_x348_TID, // @[:@27431.4]
  input  [7:0]   io_in_x348_TDEST, // @[:@27431.4]
  output         io_in_x349_TVALID, // @[:@27431.4]
  input          io_in_x349_TREADY, // @[:@27431.4]
  output [255:0] io_in_x349_TDATA, // @[:@27431.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@27431.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@27431.4]
  input          io_sigsIn_smChildAcks_0, // @[:@27431.4]
  input          io_sigsIn_smChildAcks_1, // @[:@27431.4]
  output         io_sigsOut_smDoneIn_0, // @[:@27431.4]
  output         io_sigsOut_smDoneIn_1, // @[:@27431.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@27431.4]
  output         io_sigsOut_smCtrCopyDone_1, // @[:@27431.4]
  input          io_rr // @[:@27431.4]
);
  wire  x351_fifoinraw_0_clock; // @[m_x351_fifoinraw_0.scala 27:17:@27445.4]
  wire  x351_fifoinraw_0_reset; // @[m_x351_fifoinraw_0.scala 27:17:@27445.4]
  wire  x352_fifoinpacked_0_clock; // @[m_x352_fifoinpacked_0.scala 27:17:@27469.4]
  wire  x352_fifoinpacked_0_reset; // @[m_x352_fifoinpacked_0.scala 27:17:@27469.4]
  wire  x352_fifoinpacked_0_io_wPort_0_en_0; // @[m_x352_fifoinpacked_0.scala 27:17:@27469.4]
  wire  x352_fifoinpacked_0_io_full; // @[m_x352_fifoinpacked_0.scala 27:17:@27469.4]
  wire  x352_fifoinpacked_0_io_active_0_in; // @[m_x352_fifoinpacked_0.scala 27:17:@27469.4]
  wire  x352_fifoinpacked_0_io_active_0_out; // @[m_x352_fifoinpacked_0.scala 27:17:@27469.4]
  wire  x353_fifooutraw_0_clock; // @[m_x353_fifooutraw_0.scala 27:17:@27493.4]
  wire  x353_fifooutraw_0_reset; // @[m_x353_fifooutraw_0.scala 27:17:@27493.4]
  wire  x356_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@27517.4]
  wire  x356_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@27517.4]
  wire  x356_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@27517.4]
  wire  x356_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@27517.4]
  wire [12:0] x356_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@27517.4]
  wire [12:0] x356_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@27517.4]
  wire  x356_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@27517.4]
  wire  x356_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@27517.4]
  wire  x356_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@27517.4]
  wire  x374_inr_Foreach_sm_clock; // @[sm_x374_inr_Foreach.scala 32:18:@27577.4]
  wire  x374_inr_Foreach_sm_reset; // @[sm_x374_inr_Foreach.scala 32:18:@27577.4]
  wire  x374_inr_Foreach_sm_io_enable; // @[sm_x374_inr_Foreach.scala 32:18:@27577.4]
  wire  x374_inr_Foreach_sm_io_done; // @[sm_x374_inr_Foreach.scala 32:18:@27577.4]
  wire  x374_inr_Foreach_sm_io_doneLatch; // @[sm_x374_inr_Foreach.scala 32:18:@27577.4]
  wire  x374_inr_Foreach_sm_io_ctrDone; // @[sm_x374_inr_Foreach.scala 32:18:@27577.4]
  wire  x374_inr_Foreach_sm_io_datapathEn; // @[sm_x374_inr_Foreach.scala 32:18:@27577.4]
  wire  x374_inr_Foreach_sm_io_ctrInc; // @[sm_x374_inr_Foreach.scala 32:18:@27577.4]
  wire  x374_inr_Foreach_sm_io_ctrRst; // @[sm_x374_inr_Foreach.scala 32:18:@27577.4]
  wire  x374_inr_Foreach_sm_io_parentAck; // @[sm_x374_inr_Foreach.scala 32:18:@27577.4]
  wire  x374_inr_Foreach_sm_io_backpressure; // @[sm_x374_inr_Foreach.scala 32:18:@27577.4]
  wire  x374_inr_Foreach_sm_io_break; // @[sm_x374_inr_Foreach.scala 32:18:@27577.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@27605.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@27605.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@27605.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@27605.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@27605.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@27651.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@27651.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@27651.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@27651.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@27651.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@27659.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@27659.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@27659.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@27659.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@27659.4]
  wire  x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_clock; // @[sm_x374_inr_Foreach.scala 106:24:@27694.4]
  wire  x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_reset; // @[sm_x374_inr_Foreach.scala 106:24:@27694.4]
  wire  x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_in_x352_fifoinpacked_0_wPort_0_en_0; // @[sm_x374_inr_Foreach.scala 106:24:@27694.4]
  wire  x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_in_x352_fifoinpacked_0_full; // @[sm_x374_inr_Foreach.scala 106:24:@27694.4]
  wire  x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_in_x352_fifoinpacked_0_active_0_in; // @[sm_x374_inr_Foreach.scala 106:24:@27694.4]
  wire  x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_in_x352_fifoinpacked_0_active_0_out; // @[sm_x374_inr_Foreach.scala 106:24:@27694.4]
  wire  x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x374_inr_Foreach.scala 106:24:@27694.4]
  wire  x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x374_inr_Foreach.scala 106:24:@27694.4]
  wire  x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x374_inr_Foreach.scala 106:24:@27694.4]
  wire [31:0] x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x374_inr_Foreach.scala 106:24:@27694.4]
  wire [31:0] x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x374_inr_Foreach.scala 106:24:@27694.4]
  wire  x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x374_inr_Foreach.scala 106:24:@27694.4]
  wire  x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x374_inr_Foreach.scala 106:24:@27694.4]
  wire  x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_rr; // @[sm_x374_inr_Foreach.scala 106:24:@27694.4]
  wire  x527_outr_UnitPipe_sm_clock; // @[sm_x527_outr_UnitPipe.scala 32:18:@27826.4]
  wire  x527_outr_UnitPipe_sm_reset; // @[sm_x527_outr_UnitPipe.scala 32:18:@27826.4]
  wire  x527_outr_UnitPipe_sm_io_enable; // @[sm_x527_outr_UnitPipe.scala 32:18:@27826.4]
  wire  x527_outr_UnitPipe_sm_io_done; // @[sm_x527_outr_UnitPipe.scala 32:18:@27826.4]
  wire  x527_outr_UnitPipe_sm_io_rst; // @[sm_x527_outr_UnitPipe.scala 32:18:@27826.4]
  wire  x527_outr_UnitPipe_sm_io_ctrDone; // @[sm_x527_outr_UnitPipe.scala 32:18:@27826.4]
  wire  x527_outr_UnitPipe_sm_io_ctrInc; // @[sm_x527_outr_UnitPipe.scala 32:18:@27826.4]
  wire  x527_outr_UnitPipe_sm_io_parentAck; // @[sm_x527_outr_UnitPipe.scala 32:18:@27826.4]
  wire  x527_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x527_outr_UnitPipe.scala 32:18:@27826.4]
  wire  x527_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x527_outr_UnitPipe.scala 32:18:@27826.4]
  wire  x527_outr_UnitPipe_sm_io_childAck_0; // @[sm_x527_outr_UnitPipe.scala 32:18:@27826.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@27883.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@27883.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@27883.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@27883.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@27883.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@27891.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@27891.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@27891.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@27891.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@27891.4]
  wire  x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_clock; // @[sm_x527_outr_UnitPipe.scala 76:24:@27921.4]
  wire  x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_reset; // @[sm_x527_outr_UnitPipe.scala 76:24:@27921.4]
  wire  x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x348_TVALID; // @[sm_x527_outr_UnitPipe.scala 76:24:@27921.4]
  wire  x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x348_TREADY; // @[sm_x527_outr_UnitPipe.scala 76:24:@27921.4]
  wire [255:0] x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x348_TDATA; // @[sm_x527_outr_UnitPipe.scala 76:24:@27921.4]
  wire [7:0] x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x348_TID; // @[sm_x527_outr_UnitPipe.scala 76:24:@27921.4]
  wire [7:0] x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x348_TDEST; // @[sm_x527_outr_UnitPipe.scala 76:24:@27921.4]
  wire  x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x349_TVALID; // @[sm_x527_outr_UnitPipe.scala 76:24:@27921.4]
  wire  x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x349_TREADY; // @[sm_x527_outr_UnitPipe.scala 76:24:@27921.4]
  wire [255:0] x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x349_TDATA; // @[sm_x527_outr_UnitPipe.scala 76:24:@27921.4]
  wire  x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x527_outr_UnitPipe.scala 76:24:@27921.4]
  wire  x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x527_outr_UnitPipe.scala 76:24:@27921.4]
  wire  x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x527_outr_UnitPipe.scala 76:24:@27921.4]
  wire  x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_rr; // @[sm_x527_outr_UnitPipe.scala 76:24:@27921.4]
  wire  _T_254; // @[package.scala 96:25:@27610.4 package.scala 96:25:@27611.4]
  wire  _T_260; // @[implicits.scala 47:10:@27614.4]
  wire  _T_261; // @[sm_x528_outr_UnitPipe.scala 70:41:@27615.4]
  wire  _T_262; // @[sm_x528_outr_UnitPipe.scala 70:78:@27616.4]
  wire  _T_263; // @[sm_x528_outr_UnitPipe.scala 70:76:@27617.4]
  wire  _T_275; // @[package.scala 96:25:@27656.4 package.scala 96:25:@27657.4]
  wire  _T_281; // @[package.scala 96:25:@27664.4 package.scala 96:25:@27665.4]
  wire  _T_284; // @[SpatialBlocks.scala 138:93:@27667.4]
  wire  _T_286; // @[SpatialBlocks.scala 157:36:@27676.4]
  wire  _T_287; // @[SpatialBlocks.scala 157:78:@27677.4]
  wire  _T_354; // @[package.scala 100:49:@27854.4]
  reg  _T_357; // @[package.scala 48:56:@27855.4]
  reg [31:0] _RAND_0;
  wire  _T_371; // @[package.scala 96:25:@27888.4 package.scala 96:25:@27889.4]
  wire  _T_377; // @[package.scala 96:25:@27896.4 package.scala 96:25:@27897.4]
  wire  _T_380; // @[SpatialBlocks.scala 138:93:@27899.4]
  x351_fifoinraw_0 x351_fifoinraw_0 ( // @[m_x351_fifoinraw_0.scala 27:17:@27445.4]
    .clock(x351_fifoinraw_0_clock),
    .reset(x351_fifoinraw_0_reset)
  );
  x352_fifoinpacked_0 x352_fifoinpacked_0 ( // @[m_x352_fifoinpacked_0.scala 27:17:@27469.4]
    .clock(x352_fifoinpacked_0_clock),
    .reset(x352_fifoinpacked_0_reset),
    .io_wPort_0_en_0(x352_fifoinpacked_0_io_wPort_0_en_0),
    .io_full(x352_fifoinpacked_0_io_full),
    .io_active_0_in(x352_fifoinpacked_0_io_active_0_in),
    .io_active_0_out(x352_fifoinpacked_0_io_active_0_out)
  );
  x351_fifoinraw_0 x353_fifooutraw_0 ( // @[m_x353_fifooutraw_0.scala 27:17:@27493.4]
    .clock(x353_fifooutraw_0_clock),
    .reset(x353_fifooutraw_0_reset)
  );
  x356_ctrchain x356_ctrchain ( // @[SpatialBlocks.scala 37:22:@27517.4]
    .clock(x356_ctrchain_clock),
    .reset(x356_ctrchain_reset),
    .io_input_reset(x356_ctrchain_io_input_reset),
    .io_input_enable(x356_ctrchain_io_input_enable),
    .io_output_counts_1(x356_ctrchain_io_output_counts_1),
    .io_output_counts_0(x356_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x356_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x356_ctrchain_io_output_oobs_1),
    .io_output_done(x356_ctrchain_io_output_done)
  );
  x374_inr_Foreach_sm x374_inr_Foreach_sm ( // @[sm_x374_inr_Foreach.scala 32:18:@27577.4]
    .clock(x374_inr_Foreach_sm_clock),
    .reset(x374_inr_Foreach_sm_reset),
    .io_enable(x374_inr_Foreach_sm_io_enable),
    .io_done(x374_inr_Foreach_sm_io_done),
    .io_doneLatch(x374_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x374_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x374_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x374_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x374_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x374_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x374_inr_Foreach_sm_io_backpressure),
    .io_break(x374_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@27605.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@27651.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@27659.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x374_inr_Foreach_kernelx374_inr_Foreach_concrete1 x374_inr_Foreach_kernelx374_inr_Foreach_concrete1 ( // @[sm_x374_inr_Foreach.scala 106:24:@27694.4]
    .clock(x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_clock),
    .reset(x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_reset),
    .io_in_x352_fifoinpacked_0_wPort_0_en_0(x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_in_x352_fifoinpacked_0_wPort_0_en_0),
    .io_in_x352_fifoinpacked_0_full(x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_in_x352_fifoinpacked_0_full),
    .io_in_x352_fifoinpacked_0_active_0_in(x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_in_x352_fifoinpacked_0_active_0_in),
    .io_in_x352_fifoinpacked_0_active_0_out(x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_in_x352_fifoinpacked_0_active_0_out),
    .io_sigsIn_backpressure(x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_rr)
  );
  RootController_sm x527_outr_UnitPipe_sm ( // @[sm_x527_outr_UnitPipe.scala 32:18:@27826.4]
    .clock(x527_outr_UnitPipe_sm_clock),
    .reset(x527_outr_UnitPipe_sm_reset),
    .io_enable(x527_outr_UnitPipe_sm_io_enable),
    .io_done(x527_outr_UnitPipe_sm_io_done),
    .io_rst(x527_outr_UnitPipe_sm_io_rst),
    .io_ctrDone(x527_outr_UnitPipe_sm_io_ctrDone),
    .io_ctrInc(x527_outr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x527_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x527_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x527_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x527_outr_UnitPipe_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@27883.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@27891.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1 x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1 ( // @[sm_x527_outr_UnitPipe.scala 76:24:@27921.4]
    .clock(x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_clock),
    .reset(x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_reset),
    .io_in_x348_TVALID(x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x348_TVALID),
    .io_in_x348_TREADY(x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x348_TREADY),
    .io_in_x348_TDATA(x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x348_TDATA),
    .io_in_x348_TID(x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x348_TID),
    .io_in_x348_TDEST(x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x348_TDEST),
    .io_in_x349_TVALID(x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x349_TVALID),
    .io_in_x349_TREADY(x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x349_TREADY),
    .io_in_x349_TDATA(x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x349_TDATA),
    .io_sigsIn_smEnableOuts_0(x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_254 = RetimeWrapper_io_out; // @[package.scala 96:25:@27610.4 package.scala 96:25:@27611.4]
  assign _T_260 = x352_fifoinpacked_0_io_full; // @[implicits.scala 47:10:@27614.4]
  assign _T_261 = ~ _T_260; // @[sm_x528_outr_UnitPipe.scala 70:41:@27615.4]
  assign _T_262 = ~ x352_fifoinpacked_0_io_active_0_out; // @[sm_x528_outr_UnitPipe.scala 70:78:@27616.4]
  assign _T_263 = _T_261 | _T_262; // @[sm_x528_outr_UnitPipe.scala 70:76:@27617.4]
  assign _T_275 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@27656.4 package.scala 96:25:@27657.4]
  assign _T_281 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@27664.4 package.scala 96:25:@27665.4]
  assign _T_284 = ~ _T_281; // @[SpatialBlocks.scala 138:93:@27667.4]
  assign _T_286 = x374_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@27676.4]
  assign _T_287 = ~ x374_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@27677.4]
  assign _T_354 = x527_outr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@27854.4]
  assign _T_371 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@27888.4 package.scala 96:25:@27889.4]
  assign _T_377 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@27896.4 package.scala 96:25:@27897.4]
  assign _T_380 = ~ _T_377; // @[SpatialBlocks.scala 138:93:@27899.4]
  assign io_in_x348_TREADY = x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x348_TREADY; // @[sm_x527_outr_UnitPipe.scala 48:23:@27977.4]
  assign io_in_x349_TVALID = x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x349_TVALID; // @[sm_x527_outr_UnitPipe.scala 49:23:@27987.4]
  assign io_in_x349_TDATA = x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x349_TDATA; // @[sm_x527_outr_UnitPipe.scala 49:23:@27985.4]
  assign io_sigsOut_smDoneIn_0 = x374_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@27674.4]
  assign io_sigsOut_smDoneIn_1 = x527_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@27906.4]
  assign io_sigsOut_smCtrCopyDone_0 = x374_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@27693.4]
  assign io_sigsOut_smCtrCopyDone_1 = x527_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@27920.4]
  assign x351_fifoinraw_0_clock = clock; // @[:@27446.4]
  assign x351_fifoinraw_0_reset = reset; // @[:@27447.4]
  assign x352_fifoinpacked_0_clock = clock; // @[:@27470.4]
  assign x352_fifoinpacked_0_reset = reset; // @[:@27471.4]
  assign x352_fifoinpacked_0_io_wPort_0_en_0 = x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_in_x352_fifoinpacked_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@27754.4]
  assign x352_fifoinpacked_0_io_active_0_in = x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_in_x352_fifoinpacked_0_active_0_in; // @[MemInterfaceType.scala 167:86:@27753.4]
  assign x353_fifooutraw_0_clock = clock; // @[:@27494.4]
  assign x353_fifooutraw_0_reset = reset; // @[:@27495.4]
  assign x356_ctrchain_clock = clock; // @[:@27518.4]
  assign x356_ctrchain_reset = reset; // @[:@27519.4]
  assign x356_ctrchain_io_input_reset = x374_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@27692.4]
  assign x356_ctrchain_io_input_enable = x374_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@27644.4 SpatialBlocks.scala 159:42:@27691.4]
  assign x374_inr_Foreach_sm_clock = clock; // @[:@27578.4]
  assign x374_inr_Foreach_sm_reset = reset; // @[:@27579.4]
  assign x374_inr_Foreach_sm_io_enable = _T_275 & _T_284; // @[SpatialBlocks.scala 140:18:@27671.4]
  assign x374_inr_Foreach_sm_io_ctrDone = io_rr ? _T_254 : 1'h0; // @[sm_x528_outr_UnitPipe.scala 69:38:@27613.4]
  assign x374_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@27673.4]
  assign x374_inr_Foreach_sm_io_backpressure = _T_263 | x374_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@27645.4]
  assign x374_inr_Foreach_sm_io_break = 1'h0; // @[sm_x528_outr_UnitPipe.scala 73:36:@27623.4]
  assign RetimeWrapper_clock = clock; // @[:@27606.4]
  assign RetimeWrapper_reset = reset; // @[:@27607.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@27609.4]
  assign RetimeWrapper_io_in = x356_ctrchain_io_output_done; // @[package.scala 94:16:@27608.4]
  assign RetimeWrapper_1_clock = clock; // @[:@27652.4]
  assign RetimeWrapper_1_reset = reset; // @[:@27653.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@27655.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@27654.4]
  assign RetimeWrapper_2_clock = clock; // @[:@27660.4]
  assign RetimeWrapper_2_reset = reset; // @[:@27661.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@27663.4]
  assign RetimeWrapper_2_io_in = x374_inr_Foreach_sm_io_done; // @[package.scala 94:16:@27662.4]
  assign x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_clock = clock; // @[:@27695.4]
  assign x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_reset = reset; // @[:@27696.4]
  assign x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_in_x352_fifoinpacked_0_full = x352_fifoinpacked_0_io_full; // @[MemInterfaceType.scala 159:15:@27748.4]
  assign x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_in_x352_fifoinpacked_0_active_0_out = x352_fifoinpacked_0_io_active_0_out; // @[MemInterfaceType.scala 158:75:@27747.4]
  assign x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_263 | x374_inr_Foreach_sm_io_doneLatch; // @[sm_x374_inr_Foreach.scala 111:22:@27777.4]
  assign x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_286 & _T_287; // @[sm_x374_inr_Foreach.scala 111:22:@27775.4]
  assign x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_break = x374_inr_Foreach_sm_io_break; // @[sm_x374_inr_Foreach.scala 111:22:@27773.4]
  assign x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x356_ctrchain_io_output_counts_1[12]}},x356_ctrchain_io_output_counts_1}; // @[sm_x374_inr_Foreach.scala 111:22:@27768.4]
  assign x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x356_ctrchain_io_output_counts_0[12]}},x356_ctrchain_io_output_counts_0}; // @[sm_x374_inr_Foreach.scala 111:22:@27767.4]
  assign x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x356_ctrchain_io_output_oobs_0; // @[sm_x374_inr_Foreach.scala 111:22:@27765.4]
  assign x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x356_ctrchain_io_output_oobs_1; // @[sm_x374_inr_Foreach.scala 111:22:@27766.4]
  assign x374_inr_Foreach_kernelx374_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x374_inr_Foreach.scala 110:18:@27761.4]
  assign x527_outr_UnitPipe_sm_clock = clock; // @[:@27827.4]
  assign x527_outr_UnitPipe_sm_reset = reset; // @[:@27828.4]
  assign x527_outr_UnitPipe_sm_io_enable = _T_371 & _T_380; // @[SpatialBlocks.scala 140:18:@27903.4]
  assign x527_outr_UnitPipe_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 134:15:@27878.4]
  assign x527_outr_UnitPipe_sm_io_ctrDone = x527_outr_UnitPipe_sm_io_ctrInc & _T_357; // @[sm_x528_outr_UnitPipe.scala 78:40:@27858.4]
  assign x527_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@27905.4]
  assign x527_outr_UnitPipe_sm_io_doneIn_0 = x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@27875.4]
  assign RetimeWrapper_3_clock = clock; // @[:@27884.4]
  assign RetimeWrapper_3_reset = reset; // @[:@27885.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@27887.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@27886.4]
  assign RetimeWrapper_4_clock = clock; // @[:@27892.4]
  assign RetimeWrapper_4_reset = reset; // @[:@27893.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@27895.4]
  assign RetimeWrapper_4_io_in = x527_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@27894.4]
  assign x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_clock = clock; // @[:@27922.4]
  assign x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_reset = reset; // @[:@27923.4]
  assign x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x348_TVALID = io_in_x348_TVALID; // @[sm_x527_outr_UnitPipe.scala 48:23:@27978.4]
  assign x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x348_TDATA = io_in_x348_TDATA; // @[sm_x527_outr_UnitPipe.scala 48:23:@27976.4]
  assign x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x348_TID = io_in_x348_TID; // @[sm_x527_outr_UnitPipe.scala 48:23:@27972.4]
  assign x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x348_TDEST = io_in_x348_TDEST; // @[sm_x527_outr_UnitPipe.scala 48:23:@27971.4]
  assign x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_in_x349_TREADY = io_in_x349_TREADY; // @[sm_x527_outr_UnitPipe.scala 49:23:@27986.4]
  assign x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x527_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x527_outr_UnitPipe.scala 81:22:@27996.4]
  assign x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x527_outr_UnitPipe_sm_io_childAck_0; // @[sm_x527_outr_UnitPipe.scala 81:22:@27994.4]
  assign x527_outr_UnitPipe_kernelx527_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x527_outr_UnitPipe.scala 80:18:@27988.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_357 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_357 <= 1'h0;
    end else begin
      _T_357 <= _T_354;
    end
  end
endmodule
module x550_outr_UnitPipe_sm( // @[:@28485.2]
  input   clock, // @[:@28486.4]
  input   reset, // @[:@28487.4]
  input   io_enable, // @[:@28488.4]
  output  io_done, // @[:@28488.4]
  input   io_parentAck, // @[:@28488.4]
  input   io_doneIn_0, // @[:@28488.4]
  input   io_doneIn_1, // @[:@28488.4]
  input   io_doneIn_2, // @[:@28488.4]
  output  io_enableOut_0, // @[:@28488.4]
  output  io_enableOut_1, // @[:@28488.4]
  output  io_enableOut_2, // @[:@28488.4]
  output  io_childAck_0, // @[:@28488.4]
  output  io_childAck_1, // @[:@28488.4]
  output  io_childAck_2, // @[:@28488.4]
  input   io_ctrCopyDone_0, // @[:@28488.4]
  input   io_ctrCopyDone_1, // @[:@28488.4]
  input   io_ctrCopyDone_2 // @[:@28488.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@28491.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@28491.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@28491.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@28491.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@28491.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@28491.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@28494.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@28494.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@28494.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@28494.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@28494.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@28494.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@28497.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@28497.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@28497.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@28497.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@28497.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@28497.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@28500.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@28500.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@28500.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@28500.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@28500.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@28500.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@28503.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@28503.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@28503.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@28503.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@28503.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@28503.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@28506.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@28506.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@28506.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@28506.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@28506.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@28506.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@28547.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@28547.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@28547.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@28547.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@28547.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@28547.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@28550.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@28550.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@28550.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@28550.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@28550.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@28550.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@28553.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@28553.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@28553.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@28553.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@28553.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@28553.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@28604.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@28604.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@28604.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@28604.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@28604.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@28618.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@28618.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@28618.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@28618.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@28618.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@28636.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@28636.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@28636.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@28636.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@28636.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@28673.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@28673.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@28673.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@28673.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@28673.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@28687.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@28687.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@28687.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@28687.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@28687.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@28705.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@28705.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@28705.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@28705.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@28705.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@28742.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@28742.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@28742.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@28742.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@28742.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@28756.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@28756.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@28756.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@28756.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@28756.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@28774.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@28774.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@28774.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@28774.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@28774.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@28831.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@28831.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@28831.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@28831.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@28831.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@28848.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@28848.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@28848.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@28848.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@28848.4]
  wire  _T_77; // @[Controllers.scala 80:47:@28509.4]
  wire  allDone; // @[Controllers.scala 80:47:@28510.4]
  wire  _T_151; // @[Controllers.scala 165:35:@28588.4]
  wire  _T_153; // @[Controllers.scala 165:60:@28589.4]
  wire  _T_154; // @[Controllers.scala 165:58:@28590.4]
  wire  _T_156; // @[Controllers.scala 165:76:@28591.4]
  wire  _T_157; // @[Controllers.scala 165:74:@28592.4]
  wire  _T_161; // @[Controllers.scala 165:109:@28595.4]
  wire  _T_164; // @[Controllers.scala 165:141:@28597.4]
  wire  _T_172; // @[package.scala 96:25:@28609.4 package.scala 96:25:@28610.4]
  wire  _T_176; // @[Controllers.scala 167:54:@28612.4]
  wire  _T_177; // @[Controllers.scala 167:52:@28613.4]
  wire  _T_184; // @[package.scala 96:25:@28623.4 package.scala 96:25:@28624.4]
  wire  _T_202; // @[package.scala 96:25:@28641.4 package.scala 96:25:@28642.4]
  wire  _T_206; // @[Controllers.scala 169:67:@28644.4]
  wire  _T_207; // @[Controllers.scala 169:86:@28645.4]
  wire  _T_219; // @[Controllers.scala 165:35:@28657.4]
  wire  _T_221; // @[Controllers.scala 165:60:@28658.4]
  wire  _T_222; // @[Controllers.scala 165:58:@28659.4]
  wire  _T_224; // @[Controllers.scala 165:76:@28660.4]
  wire  _T_225; // @[Controllers.scala 165:74:@28661.4]
  wire  _T_229; // @[Controllers.scala 165:109:@28664.4]
  wire  _T_232; // @[Controllers.scala 165:141:@28666.4]
  wire  _T_240; // @[package.scala 96:25:@28678.4 package.scala 96:25:@28679.4]
  wire  _T_244; // @[Controllers.scala 167:54:@28681.4]
  wire  _T_245; // @[Controllers.scala 167:52:@28682.4]
  wire  _T_252; // @[package.scala 96:25:@28692.4 package.scala 96:25:@28693.4]
  wire  _T_270; // @[package.scala 96:25:@28710.4 package.scala 96:25:@28711.4]
  wire  _T_274; // @[Controllers.scala 169:67:@28713.4]
  wire  _T_275; // @[Controllers.scala 169:86:@28714.4]
  wire  _T_287; // @[Controllers.scala 165:35:@28726.4]
  wire  _T_289; // @[Controllers.scala 165:60:@28727.4]
  wire  _T_290; // @[Controllers.scala 165:58:@28728.4]
  wire  _T_292; // @[Controllers.scala 165:76:@28729.4]
  wire  _T_293; // @[Controllers.scala 165:74:@28730.4]
  wire  _T_297; // @[Controllers.scala 165:109:@28733.4]
  wire  _T_300; // @[Controllers.scala 165:141:@28735.4]
  wire  _T_308; // @[package.scala 96:25:@28747.4 package.scala 96:25:@28748.4]
  wire  _T_312; // @[Controllers.scala 167:54:@28750.4]
  wire  _T_313; // @[Controllers.scala 167:52:@28751.4]
  wire  _T_320; // @[package.scala 96:25:@28761.4 package.scala 96:25:@28762.4]
  wire  _T_338; // @[package.scala 96:25:@28779.4 package.scala 96:25:@28780.4]
  wire  _T_342; // @[Controllers.scala 169:67:@28782.4]
  wire  _T_343; // @[Controllers.scala 169:86:@28783.4]
  wire  _T_358; // @[Controllers.scala 213:68:@28801.4]
  wire  _T_360; // @[Controllers.scala 213:90:@28803.4]
  wire  _T_362; // @[Controllers.scala 213:132:@28805.4]
  wire  _T_366; // @[Controllers.scala 213:68:@28810.4]
  wire  _T_368; // @[Controllers.scala 213:90:@28812.4]
  wire  _T_374; // @[Controllers.scala 213:68:@28818.4]
  wire  _T_376; // @[Controllers.scala 213:90:@28820.4]
  wire  _T_383; // @[package.scala 100:49:@28826.4]
  reg  _T_386; // @[package.scala 48:56:@28827.4]
  reg [31:0] _RAND_0;
  wire  _T_387; // @[package.scala 100:41:@28829.4]
  reg  _T_400; // @[package.scala 48:56:@28845.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@28491.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@28494.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@28497.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@28500.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@28503.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@28506.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@28547.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@28550.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@28553.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@28604.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@28618.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@28636.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@28673.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@28687.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@28705.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@28742.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@28756.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@28774.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@28831.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@28848.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@28509.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@28510.4]
  assign _T_151 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@28588.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@28589.4]
  assign _T_154 = _T_151 & _T_153; // @[Controllers.scala 165:58:@28590.4]
  assign _T_156 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@28591.4]
  assign _T_157 = _T_154 & _T_156; // @[Controllers.scala 165:74:@28592.4]
  assign _T_161 = _T_157 & io_enable; // @[Controllers.scala 165:109:@28595.4]
  assign _T_164 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@28597.4]
  assign _T_172 = RetimeWrapper_io_out; // @[package.scala 96:25:@28609.4 package.scala 96:25:@28610.4]
  assign _T_176 = _T_172 == 1'h0; // @[Controllers.scala 167:54:@28612.4]
  assign _T_177 = io_doneIn_0 | _T_176; // @[Controllers.scala 167:52:@28613.4]
  assign _T_184 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@28623.4 package.scala 96:25:@28624.4]
  assign _T_202 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@28641.4 package.scala 96:25:@28642.4]
  assign _T_206 = _T_202 == 1'h0; // @[Controllers.scala 169:67:@28644.4]
  assign _T_207 = _T_206 & io_enable; // @[Controllers.scala 169:86:@28645.4]
  assign _T_219 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@28657.4]
  assign _T_221 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@28658.4]
  assign _T_222 = _T_219 & _T_221; // @[Controllers.scala 165:58:@28659.4]
  assign _T_224 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@28660.4]
  assign _T_225 = _T_222 & _T_224; // @[Controllers.scala 165:74:@28661.4]
  assign _T_229 = _T_225 & io_enable; // @[Controllers.scala 165:109:@28664.4]
  assign _T_232 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@28666.4]
  assign _T_240 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@28678.4 package.scala 96:25:@28679.4]
  assign _T_244 = _T_240 == 1'h0; // @[Controllers.scala 167:54:@28681.4]
  assign _T_245 = io_doneIn_1 | _T_244; // @[Controllers.scala 167:52:@28682.4]
  assign _T_252 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@28692.4 package.scala 96:25:@28693.4]
  assign _T_270 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@28710.4 package.scala 96:25:@28711.4]
  assign _T_274 = _T_270 == 1'h0; // @[Controllers.scala 169:67:@28713.4]
  assign _T_275 = _T_274 & io_enable; // @[Controllers.scala 169:86:@28714.4]
  assign _T_287 = ~ iterDone_2_io_output; // @[Controllers.scala 165:35:@28726.4]
  assign _T_289 = io_doneIn_2 == 1'h0; // @[Controllers.scala 165:60:@28727.4]
  assign _T_290 = _T_287 & _T_289; // @[Controllers.scala 165:58:@28728.4]
  assign _T_292 = done_2_io_output == 1'h0; // @[Controllers.scala 165:76:@28729.4]
  assign _T_293 = _T_290 & _T_292; // @[Controllers.scala 165:74:@28730.4]
  assign _T_297 = _T_293 & io_enable; // @[Controllers.scala 165:109:@28733.4]
  assign _T_300 = io_ctrCopyDone_2 == 1'h0; // @[Controllers.scala 165:141:@28735.4]
  assign _T_308 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@28747.4 package.scala 96:25:@28748.4]
  assign _T_312 = _T_308 == 1'h0; // @[Controllers.scala 167:54:@28750.4]
  assign _T_313 = io_doneIn_2 | _T_312; // @[Controllers.scala 167:52:@28751.4]
  assign _T_320 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@28761.4 package.scala 96:25:@28762.4]
  assign _T_338 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@28779.4 package.scala 96:25:@28780.4]
  assign _T_342 = _T_338 == 1'h0; // @[Controllers.scala 169:67:@28782.4]
  assign _T_343 = _T_342 & io_enable; // @[Controllers.scala 169:86:@28783.4]
  assign _T_358 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@28801.4]
  assign _T_360 = _T_358 & _T_151; // @[Controllers.scala 213:90:@28803.4]
  assign _T_362 = ~ allDone; // @[Controllers.scala 213:132:@28805.4]
  assign _T_366 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@28810.4]
  assign _T_368 = _T_366 & _T_219; // @[Controllers.scala 213:90:@28812.4]
  assign _T_374 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@28818.4]
  assign _T_376 = _T_374 & _T_287; // @[Controllers.scala 213:90:@28820.4]
  assign _T_383 = allDone == 1'h0; // @[package.scala 100:49:@28826.4]
  assign _T_387 = allDone & _T_386; // @[package.scala 100:41:@28829.4]
  assign io_done = RetimeWrapper_10_io_out; // @[Controllers.scala 245:13:@28855.4]
  assign io_enableOut_0 = _T_360 & _T_362; // @[Controllers.scala 213:55:@28809.4]
  assign io_enableOut_1 = _T_368 & _T_362; // @[Controllers.scala 213:55:@28817.4]
  assign io_enableOut_2 = _T_376 & _T_362; // @[Controllers.scala 213:55:@28825.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@28796.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@28798.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@28800.4]
  assign active_0_clock = clock; // @[:@28492.4]
  assign active_0_reset = reset; // @[:@28493.4]
  assign active_0_io_input_set = _T_161 & _T_164; // @[Controllers.scala 165:32:@28599.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@28603.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@28513.4]
  assign active_1_clock = clock; // @[:@28495.4]
  assign active_1_reset = reset; // @[:@28496.4]
  assign active_1_io_input_set = _T_229 & _T_232; // @[Controllers.scala 165:32:@28668.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@28672.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@28514.4]
  assign active_2_clock = clock; // @[:@28498.4]
  assign active_2_reset = reset; // @[:@28499.4]
  assign active_2_io_input_set = _T_297 & _T_300; // @[Controllers.scala 165:32:@28737.4]
  assign active_2_io_input_reset = io_ctrCopyDone_2 | io_parentAck; // @[Controllers.scala 166:34:@28741.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@28515.4]
  assign done_0_clock = clock; // @[:@28501.4]
  assign done_0_reset = reset; // @[:@28502.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_207; // @[Controllers.scala 169:30:@28649.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@28527.4 Controllers.scala 170:32:@28656.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@28516.4]
  assign done_1_clock = clock; // @[:@28504.4]
  assign done_1_reset = reset; // @[:@28505.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_275; // @[Controllers.scala 169:30:@28718.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@28536.4 Controllers.scala 170:32:@28725.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@28517.4]
  assign done_2_clock = clock; // @[:@28507.4]
  assign done_2_reset = reset; // @[:@28508.4]
  assign done_2_io_input_set = io_ctrCopyDone_2 | _T_343; // @[Controllers.scala 169:30:@28787.4]
  assign done_2_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@28545.4 Controllers.scala 170:32:@28794.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@28518.4]
  assign iterDone_0_clock = clock; // @[:@28548.4]
  assign iterDone_0_reset = reset; // @[:@28549.4]
  assign iterDone_0_io_input_set = _T_177 & io_enable; // @[Controllers.scala 167:34:@28617.4]
  assign iterDone_0_io_input_reset = _T_184 | io_parentAck; // @[Controllers.scala 92:37:@28567.4 Controllers.scala 168:36:@28633.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@28556.4]
  assign iterDone_1_clock = clock; // @[:@28551.4]
  assign iterDone_1_reset = reset; // @[:@28552.4]
  assign iterDone_1_io_input_set = _T_245 & io_enable; // @[Controllers.scala 167:34:@28686.4]
  assign iterDone_1_io_input_reset = _T_252 | io_parentAck; // @[Controllers.scala 92:37:@28576.4 Controllers.scala 168:36:@28702.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@28557.4]
  assign iterDone_2_clock = clock; // @[:@28554.4]
  assign iterDone_2_reset = reset; // @[:@28555.4]
  assign iterDone_2_io_input_set = _T_313 & io_enable; // @[Controllers.scala 167:34:@28755.4]
  assign iterDone_2_io_input_reset = _T_320 | io_parentAck; // @[Controllers.scala 92:37:@28585.4 Controllers.scala 168:36:@28771.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@28558.4]
  assign RetimeWrapper_clock = clock; // @[:@28605.4]
  assign RetimeWrapper_reset = reset; // @[:@28606.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@28608.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@28607.4]
  assign RetimeWrapper_1_clock = clock; // @[:@28619.4]
  assign RetimeWrapper_1_reset = reset; // @[:@28620.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@28622.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@28621.4]
  assign RetimeWrapper_2_clock = clock; // @[:@28637.4]
  assign RetimeWrapper_2_reset = reset; // @[:@28638.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@28640.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@28639.4]
  assign RetimeWrapper_3_clock = clock; // @[:@28674.4]
  assign RetimeWrapper_3_reset = reset; // @[:@28675.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@28677.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@28676.4]
  assign RetimeWrapper_4_clock = clock; // @[:@28688.4]
  assign RetimeWrapper_4_reset = reset; // @[:@28689.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@28691.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@28690.4]
  assign RetimeWrapper_5_clock = clock; // @[:@28706.4]
  assign RetimeWrapper_5_reset = reset; // @[:@28707.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@28709.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@28708.4]
  assign RetimeWrapper_6_clock = clock; // @[:@28743.4]
  assign RetimeWrapper_6_reset = reset; // @[:@28744.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@28746.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@28745.4]
  assign RetimeWrapper_7_clock = clock; // @[:@28757.4]
  assign RetimeWrapper_7_reset = reset; // @[:@28758.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@28760.4]
  assign RetimeWrapper_7_io_in = io_doneIn_2; // @[package.scala 94:16:@28759.4]
  assign RetimeWrapper_8_clock = clock; // @[:@28775.4]
  assign RetimeWrapper_8_reset = reset; // @[:@28776.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@28778.4]
  assign RetimeWrapper_8_io_in = 1'h1; // @[package.scala 94:16:@28777.4]
  assign RetimeWrapper_9_clock = clock; // @[:@28832.4]
  assign RetimeWrapper_9_reset = reset; // @[:@28833.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@28835.4]
  assign RetimeWrapper_9_io_in = _T_387 | io_parentAck; // @[package.scala 94:16:@28834.4]
  assign RetimeWrapper_10_clock = clock; // @[:@28849.4]
  assign RetimeWrapper_10_reset = reset; // @[:@28850.4]
  assign RetimeWrapper_10_io_flow = io_enable; // @[package.scala 95:18:@28852.4]
  assign RetimeWrapper_10_io_in = allDone & _T_400; // @[package.scala 94:16:@28851.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_386 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_400 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_386 <= 1'h0;
    end else begin
      _T_386 <= _T_383;
    end
    if (reset) begin
      _T_400 <= 1'h0;
    end else begin
      _T_400 <= _T_383;
    end
  end
endmodule
module x536_inr_UnitPipe_sm( // @[:@29028.2]
  input   clock, // @[:@29029.4]
  input   reset, // @[:@29030.4]
  input   io_enable, // @[:@29031.4]
  output  io_done, // @[:@29031.4]
  output  io_doneLatch, // @[:@29031.4]
  input   io_ctrDone, // @[:@29031.4]
  output  io_datapathEn, // @[:@29031.4]
  output  io_ctrInc, // @[:@29031.4]
  input   io_parentAck, // @[:@29031.4]
  input   io_backpressure // @[:@29031.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@29033.4]
  wire  active_reset; // @[Controllers.scala 261:22:@29033.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@29033.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@29033.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@29033.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@29033.4]
  wire  done_clock; // @[Controllers.scala 262:20:@29036.4]
  wire  done_reset; // @[Controllers.scala 262:20:@29036.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@29036.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@29036.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@29036.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@29036.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@29090.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@29090.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@29090.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@29090.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@29090.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@29098.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@29098.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@29098.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@29098.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@29098.4]
  wire  _T_80; // @[Controllers.scala 264:48:@29041.4]
  wire  _T_81; // @[Controllers.scala 264:46:@29042.4]
  wire  _T_82; // @[Controllers.scala 264:62:@29043.4]
  wire  _T_83; // @[Controllers.scala 264:60:@29044.4]
  wire  _T_100; // @[package.scala 100:49:@29061.4]
  reg  _T_103; // @[package.scala 48:56:@29062.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 100:49:@29070.4]
  wire  _T_116; // @[Controllers.scala 283:41:@29078.4]
  wire  _T_117; // @[Controllers.scala 283:59:@29079.4]
  wire  _T_119; // @[Controllers.scala 284:37:@29082.4]
  reg  _T_125; // @[package.scala 48:56:@29086.4]
  reg [31:0] _RAND_1;
  reg  _T_142; // @[Controllers.scala 291:31:@29108.4]
  reg [31:0] _RAND_2;
  reg  _T_149; // @[package.scala 48:56:@29111.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:41:@29113.4]
  wire  _T_152; // @[Controllers.scala 292:61:@29114.4]
  wire  _T_153; // @[Controllers.scala 292:24:@29115.4]
  SRFF active ( // @[Controllers.scala 261:22:@29033.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@29036.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@29090.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@29098.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@29041.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@29042.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@29043.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@29044.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@29061.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 100:49:@29070.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@29078.4]
  assign _T_117 = _T_116 & io_enable; // @[Controllers.scala 283:59:@29079.4]
  assign _T_119 = active_io_output & io_enable; // @[Controllers.scala 284:37:@29082.4]
  assign _T_150 = done_io_output & _T_149; // @[package.scala 100:41:@29113.4]
  assign _T_152 = _T_150 ? 1'h1 : _T_142; // @[Controllers.scala 292:61:@29114.4]
  assign _T_153 = io_parentAck ? 1'h0 : _T_152; // @[Controllers.scala 292:24:@29115.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@29089.4]
  assign io_doneLatch = _T_142; // @[Controllers.scala 293:18:@29117.4]
  assign io_datapathEn = _T_117 & io_backpressure; // @[Controllers.scala 283:21:@29081.4]
  assign io_ctrInc = _T_119 & io_backpressure; // @[Controllers.scala 284:17:@29084.4]
  assign active_clock = clock; // @[:@29034.4]
  assign active_reset = reset; // @[:@29035.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@29046.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@29050.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@29051.4]
  assign done_clock = clock; // @[:@29037.4]
  assign done_reset = reset; // @[:@29038.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@29066.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@29059.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@29060.4]
  assign RetimeWrapper_clock = clock; // @[:@29091.4]
  assign RetimeWrapper_reset = reset; // @[:@29092.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@29094.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@29093.4]
  assign RetimeWrapper_1_clock = clock; // @[:@29099.4]
  assign RetimeWrapper_1_reset = reset; // @[:@29100.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@29102.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 94:16:@29101.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_125 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_142 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_149 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_142 <= 1'h0;
      end else begin
        if (_T_150) begin
          _T_142 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_108;
    end
  end
endmodule
module x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1( // @[:@29192.2]
  output        io_in_x529_valid, // @[:@29195.4]
  output [63:0] io_in_x529_bits_addr, // @[:@29195.4]
  output [31:0] io_in_x529_bits_size, // @[:@29195.4]
  input  [63:0] io_in_x346_outdram_number, // @[:@29195.4]
  input         io_sigsIn_backpressure, // @[:@29195.4]
  input         io_sigsIn_datapathEn, // @[:@29195.4]
  input         io_rr // @[:@29195.4]
);
  wire [96:0] x533_tuple; // @[Cat.scala 30:58:@29209.4]
  wire  _T_135; // @[implicits.scala 55:10:@29212.4]
  assign x533_tuple = {33'h1fa400,io_in_x346_outdram_number}; // @[Cat.scala 30:58:@29209.4]
  assign _T_135 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@29212.4]
  assign io_in_x529_valid = _T_135 & io_sigsIn_backpressure; // @[sm_x536_inr_UnitPipe.scala 65:18:@29215.4]
  assign io_in_x529_bits_addr = x533_tuple[63:0]; // @[sm_x536_inr_UnitPipe.scala 66:22:@29217.4]
  assign io_in_x529_bits_size = x533_tuple[95:64]; // @[sm_x536_inr_UnitPipe.scala 67:22:@29219.4]
endmodule
module FF_13( // @[:@29221.2]
  input         clock, // @[:@29222.4]
  input         reset, // @[:@29223.4]
  output [22:0] io_rPort_0_output_0, // @[:@29224.4]
  input  [22:0] io_wPort_0_data_0, // @[:@29224.4]
  input         io_wPort_0_reset, // @[:@29224.4]
  input         io_wPort_0_en_0 // @[:@29224.4]
);
  reg [22:0] ff; // @[MemPrimitives.scala 311:19:@29239.4]
  reg [31:0] _RAND_0;
  wire [22:0] _T_68; // @[MemPrimitives.scala 315:32:@29241.4]
  wire [22:0] _T_69; // @[MemPrimitives.scala 315:12:@29242.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 315:32:@29241.4]
  assign _T_69 = io_wPort_0_reset ? 23'h0 : _T_68; // @[MemPrimitives.scala 315:12:@29242.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 316:34:@29244.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[22:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 23'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 23'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_5( // @[:@29259.2]
  input         clock, // @[:@29260.4]
  input         reset, // @[:@29261.4]
  input         io_input_reset, // @[:@29262.4]
  input         io_input_enable, // @[:@29262.4]
  output [22:0] io_output_count_0, // @[:@29262.4]
  output        io_output_oobs_0, // @[:@29262.4]
  output        io_output_done // @[:@29262.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@29275.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@29275.4]
  wire [22:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@29275.4]
  wire [22:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@29275.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@29275.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@29275.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@29291.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@29291.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@29291.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@29291.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@29291.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@29291.4]
  wire  _T_36; // @[Counter.scala 264:45:@29294.4]
  wire [22:0] _T_48; // @[Counter.scala 287:52:@29319.4]
  wire [23:0] _T_50; // @[Counter.scala 291:33:@29320.4]
  wire [22:0] _T_51; // @[Counter.scala 291:33:@29321.4]
  wire [22:0] _T_52; // @[Counter.scala 291:33:@29322.4]
  wire  _T_57; // @[Counter.scala 293:18:@29324.4]
  wire [22:0] _T_68; // @[Counter.scala 299:115:@29332.4]
  wire [22:0] _T_71; // @[Counter.scala 299:152:@29335.4]
  wire [22:0] _T_72; // @[Counter.scala 299:74:@29336.4]
  wire  _T_75; // @[Counter.scala 322:102:@29340.4]
  wire  _T_77; // @[Counter.scala 322:130:@29341.4]
  FF_13 bases_0 ( // @[Counter.scala 261:53:@29275.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@29291.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@29294.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@29319.4]
  assign _T_50 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@29320.4]
  assign _T_51 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@29321.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@29322.4]
  assign _T_57 = $signed(_T_52) >= $signed(23'sh1fa400); // @[Counter.scala 293:18:@29324.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@29332.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@29335.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@29336.4]
  assign _T_75 = $signed(_T_48) < $signed(23'sh0); // @[Counter.scala 322:102:@29340.4]
  assign _T_77 = $signed(_T_48) >= $signed(23'sh1fa400); // @[Counter.scala 322:130:@29341.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@29339.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@29343.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@29345.4]
  assign bases_0_clock = clock; // @[:@29276.4]
  assign bases_0_reset = reset; // @[:@29277.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 23'h0 : _T_72; // @[Counter.scala 299:31:@29338.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@29317.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@29318.4]
  assign SRFF_clock = clock; // @[:@29292.4]
  assign SRFF_reset = reset; // @[:@29293.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@29296.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@29298.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@29299.4]
endmodule
module x538_ctrchain( // @[:@29350.2]
  input         clock, // @[:@29351.4]
  input         reset, // @[:@29352.4]
  input         io_input_reset, // @[:@29353.4]
  input         io_input_enable, // @[:@29353.4]
  output [22:0] io_output_counts_0, // @[:@29353.4]
  output        io_output_oobs_0, // @[:@29353.4]
  output        io_output_done // @[:@29353.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@29355.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@29355.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@29355.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@29355.4]
  wire [22:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@29355.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@29355.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@29355.4]
  reg  wasDone; // @[Counter.scala 542:24:@29364.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 546:69:@29370.4]
  wire  _T_47; // @[Counter.scala 546:80:@29371.4]
  reg  doneLatch; // @[Counter.scala 550:26:@29376.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 551:48:@29377.4]
  wire  _T_55; // @[Counter.scala 551:19:@29378.4]
  SingleCounter_5 ctrs_0 ( // @[Counter.scala 513:46:@29355.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 546:69:@29370.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 546:80:@29371.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@29377.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 551:19:@29378.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@29380.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@29382.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 546:18:@29373.4]
  assign ctrs_0_clock = clock; // @[:@29356.4]
  assign ctrs_0_reset = reset; // @[:@29357.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@29361.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@29362.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x545_inr_Foreach_sm( // @[:@29570.2]
  input   clock, // @[:@29571.4]
  input   reset, // @[:@29572.4]
  input   io_enable, // @[:@29573.4]
  output  io_done, // @[:@29573.4]
  output  io_doneLatch, // @[:@29573.4]
  input   io_ctrDone, // @[:@29573.4]
  output  io_datapathEn, // @[:@29573.4]
  output  io_ctrInc, // @[:@29573.4]
  output  io_ctrRst, // @[:@29573.4]
  input   io_parentAck, // @[:@29573.4]
  input   io_backpressure, // @[:@29573.4]
  input   io_break // @[:@29573.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@29575.4]
  wire  active_reset; // @[Controllers.scala 261:22:@29575.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@29575.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@29575.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@29575.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@29575.4]
  wire  done_clock; // @[Controllers.scala 262:20:@29578.4]
  wire  done_reset; // @[Controllers.scala 262:20:@29578.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@29578.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@29578.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@29578.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@29578.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@29612.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@29612.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@29612.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@29612.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@29612.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@29634.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@29634.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@29634.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@29634.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@29634.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@29646.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@29646.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@29646.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@29646.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@29646.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@29654.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@29654.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@29654.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@29654.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@29654.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@29670.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@29670.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@29670.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@29670.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@29670.4]
  wire  _T_80; // @[Controllers.scala 264:48:@29583.4]
  wire  _T_81; // @[Controllers.scala 264:46:@29584.4]
  wire  _T_82; // @[Controllers.scala 264:62:@29585.4]
  wire  _T_83; // @[Controllers.scala 264:60:@29586.4]
  wire  _T_100; // @[package.scala 100:49:@29603.4]
  reg  _T_103; // @[package.scala 48:56:@29604.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@29617.4 package.scala 96:25:@29618.4]
  wire  _T_110; // @[package.scala 100:49:@29619.4]
  reg  _T_113; // @[package.scala 48:56:@29620.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@29622.4]
  wire  _T_118; // @[Controllers.scala 283:41:@29627.4]
  wire  _T_119; // @[Controllers.scala 283:59:@29628.4]
  wire  _T_121; // @[Controllers.scala 284:37:@29631.4]
  wire  _T_124; // @[package.scala 96:25:@29639.4 package.scala 96:25:@29640.4]
  wire  _T_126; // @[package.scala 100:49:@29641.4]
  reg  _T_129; // @[package.scala 48:56:@29642.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@29664.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@29666.4]
  reg  _T_153; // @[package.scala 48:56:@29667.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@29675.4 package.scala 96:25:@29676.4]
  wire  _T_158; // @[Controllers.scala 292:61:@29677.4]
  wire  _T_159; // @[Controllers.scala 292:24:@29678.4]
  SRFF active ( // @[Controllers.scala 261:22:@29575.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@29578.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@29612.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@29634.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@29646.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@29654.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@29670.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@29583.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@29584.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@29585.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@29586.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@29603.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@29617.4 package.scala 96:25:@29618.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@29619.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@29622.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@29627.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@29628.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@29631.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@29639.4 package.scala 96:25:@29640.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@29641.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@29666.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@29675.4 package.scala 96:25:@29676.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@29677.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@29678.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@29645.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@29680.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@29630.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@29633.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@29625.4]
  assign active_clock = clock; // @[:@29576.4]
  assign active_reset = reset; // @[:@29577.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@29588.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@29592.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@29593.4]
  assign done_clock = clock; // @[:@29579.4]
  assign done_reset = reset; // @[:@29580.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@29608.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@29601.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@29602.4]
  assign RetimeWrapper_clock = clock; // @[:@29613.4]
  assign RetimeWrapper_reset = reset; // @[:@29614.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@29616.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@29615.4]
  assign RetimeWrapper_1_clock = clock; // @[:@29635.4]
  assign RetimeWrapper_1_reset = reset; // @[:@29636.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@29638.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@29637.4]
  assign RetimeWrapper_2_clock = clock; // @[:@29647.4]
  assign RetimeWrapper_2_reset = reset; // @[:@29648.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@29650.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@29649.4]
  assign RetimeWrapper_3_clock = clock; // @[:@29655.4]
  assign RetimeWrapper_3_reset = reset; // @[:@29656.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@29658.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@29657.4]
  assign RetimeWrapper_4_clock = clock; // @[:@29671.4]
  assign RetimeWrapper_4_reset = reset; // @[:@29672.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@29674.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@29673.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x545_inr_Foreach_kernelx545_inr_Foreach_concrete1( // @[:@29892.2]
  input         clock, // @[:@29893.4]
  input         reset, // @[:@29894.4]
  output        io_in_x530_valid, // @[:@29895.4]
  output [7:0]  io_in_x530_bits_wdata_0, // @[:@29895.4]
  output        io_in_x530_bits_wstrb, // @[:@29895.4]
  output [20:0] io_in_x350_outbuf_0_rPort_0_ofs_0, // @[:@29895.4]
  output        io_in_x350_outbuf_0_rPort_0_en_0, // @[:@29895.4]
  output        io_in_x350_outbuf_0_rPort_0_backpressure, // @[:@29895.4]
  input  [7:0]  io_in_x350_outbuf_0_rPort_0_output_0, // @[:@29895.4]
  input         io_sigsIn_backpressure, // @[:@29895.4]
  input         io_sigsIn_datapathEn, // @[:@29895.4]
  input         io_sigsIn_break, // @[:@29895.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@29895.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@29895.4]
  input         io_rr // @[:@29895.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@29922.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@29922.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@29951.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@29951.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@29951.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@29951.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@29951.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@29960.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@29960.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@29960.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@29960.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@29960.4]
  wire  b540; // @[sm_x545_inr_Foreach.scala 62:18:@29930.4]
  wire  _T_274; // @[sm_x545_inr_Foreach.scala 67:129:@29934.4]
  wire  _T_278; // @[implicits.scala 55:10:@29937.4]
  wire  _T_279; // @[sm_x545_inr_Foreach.scala 67:146:@29938.4]
  wire [8:0] x543_tuple; // @[Cat.scala 30:58:@29948.4]
  wire  _T_290; // @[package.scala 96:25:@29965.4 package.scala 96:25:@29966.4]
  wire  _T_292; // @[implicits.scala 55:10:@29967.4]
  wire  x685_b540_D2; // @[package.scala 96:25:@29956.4 package.scala 96:25:@29957.4]
  wire  _T_293; // @[sm_x545_inr_Foreach.scala 74:112:@29968.4]
  wire [31:0] b539_number; // @[Math.scala 712:22:@29927.4 Math.scala 713:14:@29928.4]
  _ _ ( // @[Math.scala 709:24:@29922.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@29951.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@29960.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign b540 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x545_inr_Foreach.scala 62:18:@29930.4]
  assign _T_274 = ~ io_sigsIn_break; // @[sm_x545_inr_Foreach.scala 67:129:@29934.4]
  assign _T_278 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@29937.4]
  assign _T_279 = _T_274 & _T_278; // @[sm_x545_inr_Foreach.scala 67:146:@29938.4]
  assign x543_tuple = {1'h1,io_in_x350_outbuf_0_rPort_0_output_0}; // @[Cat.scala 30:58:@29948.4]
  assign _T_290 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@29965.4 package.scala 96:25:@29966.4]
  assign _T_292 = io_rr ? _T_290 : 1'h0; // @[implicits.scala 55:10:@29967.4]
  assign x685_b540_D2 = RetimeWrapper_io_out; // @[package.scala 96:25:@29956.4 package.scala 96:25:@29957.4]
  assign _T_293 = _T_292 & x685_b540_D2; // @[sm_x545_inr_Foreach.scala 74:112:@29968.4]
  assign b539_number = __io_result; // @[Math.scala 712:22:@29927.4 Math.scala 713:14:@29928.4]
  assign io_in_x530_valid = _T_293 & io_sigsIn_backpressure; // @[sm_x545_inr_Foreach.scala 74:18:@29970.4]
  assign io_in_x530_bits_wdata_0 = x543_tuple[7:0]; // @[sm_x545_inr_Foreach.scala 75:26:@29972.4]
  assign io_in_x530_bits_wstrb = x543_tuple[8]; // @[sm_x545_inr_Foreach.scala 76:23:@29974.4]
  assign io_in_x350_outbuf_0_rPort_0_ofs_0 = b539_number[20:0]; // @[MemInterfaceType.scala 107:54:@29941.4]
  assign io_in_x350_outbuf_0_rPort_0_en_0 = _T_279 & b540; // @[MemInterfaceType.scala 110:79:@29943.4]
  assign io_in_x350_outbuf_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@29942.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@29925.4]
  assign RetimeWrapper_clock = clock; // @[:@29952.4]
  assign RetimeWrapper_reset = reset; // @[:@29953.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29955.4]
  assign RetimeWrapper_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@29954.4]
  assign RetimeWrapper_1_clock = clock; // @[:@29961.4]
  assign RetimeWrapper_1_reset = reset; // @[:@29962.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29964.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@29963.4]
endmodule
module x549_inr_UnitPipe_sm( // @[:@30130.2]
  input   clock, // @[:@30131.4]
  input   reset, // @[:@30132.4]
  input   io_enable, // @[:@30133.4]
  output  io_done, // @[:@30133.4]
  output  io_doneLatch, // @[:@30133.4]
  input   io_ctrDone, // @[:@30133.4]
  output  io_datapathEn, // @[:@30133.4]
  output  io_ctrInc, // @[:@30133.4]
  input   io_parentAck // @[:@30133.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@30135.4]
  wire  active_reset; // @[Controllers.scala 261:22:@30135.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@30135.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@30135.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@30135.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@30135.4]
  wire  done_clock; // @[Controllers.scala 262:20:@30138.4]
  wire  done_reset; // @[Controllers.scala 262:20:@30138.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@30138.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@30138.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@30138.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@30138.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@30172.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@30172.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@30172.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@30172.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@30172.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@30194.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@30194.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@30194.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@30194.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@30194.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@30206.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@30206.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@30206.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@30206.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@30206.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@30214.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@30214.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@30214.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@30214.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@30214.4]
  wire  _T_80; // @[Controllers.scala 264:48:@30143.4]
  wire  _T_81; // @[Controllers.scala 264:46:@30144.4]
  wire  _T_82; // @[Controllers.scala 264:62:@30145.4]
  wire  _T_100; // @[package.scala 100:49:@30163.4]
  reg  _T_103; // @[package.scala 48:56:@30164.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@30187.4]
  wire  _T_124; // @[package.scala 96:25:@30199.4 package.scala 96:25:@30200.4]
  wire  _T_126; // @[package.scala 100:49:@30201.4]
  reg  _T_129; // @[package.scala 48:56:@30202.4]
  reg [31:0] _RAND_1;
  reg  _T_146; // @[Controllers.scala 291:31:@30224.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@30226.4]
  reg  _T_153; // @[package.scala 48:56:@30227.4]
  reg [31:0] _RAND_3;
  wire  _T_154; // @[package.scala 100:41:@30229.4]
  wire  _T_156; // @[Controllers.scala 292:61:@30230.4]
  wire  _T_157; // @[Controllers.scala 292:24:@30231.4]
  SRFF active ( // @[Controllers.scala 261:22:@30135.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@30138.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@30172.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@30194.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@30206.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@30214.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@30143.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@30144.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@30145.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@30163.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@30187.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@30199.4 package.scala 96:25:@30200.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@30201.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@30226.4]
  assign _T_154 = done_io_output & _T_153; // @[package.scala 100:41:@30229.4]
  assign _T_156 = _T_154 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@30230.4]
  assign _T_157 = io_parentAck ? 1'h0 : _T_156; // @[Controllers.scala 292:24:@30231.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@30205.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@30233.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@30190.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@30193.4]
  assign active_clock = clock; // @[:@30136.4]
  assign active_reset = reset; // @[:@30137.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@30148.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@30152.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@30153.4]
  assign done_clock = clock; // @[:@30139.4]
  assign done_reset = reset; // @[:@30140.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@30168.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@30161.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@30162.4]
  assign RetimeWrapper_clock = clock; // @[:@30173.4]
  assign RetimeWrapper_reset = reset; // @[:@30174.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@30176.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@30175.4]
  assign RetimeWrapper_1_clock = clock; // @[:@30195.4]
  assign RetimeWrapper_1_reset = reset; // @[:@30196.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@30198.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@30197.4]
  assign RetimeWrapper_2_clock = clock; // @[:@30207.4]
  assign RetimeWrapper_2_reset = reset; // @[:@30208.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@30210.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@30209.4]
  assign RetimeWrapper_3_clock = clock; // @[:@30215.4]
  assign RetimeWrapper_3_reset = reset; // @[:@30216.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@30218.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@30217.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_154) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x549_inr_UnitPipe_kernelx549_inr_UnitPipe_concrete1( // @[:@30308.2]
  output  io_in_x531_ready, // @[:@30311.4]
  input   io_sigsIn_datapathEn // @[:@30311.4]
);
  assign io_in_x531_ready = io_sigsIn_datapathEn; // @[sm_x549_inr_UnitPipe.scala 57:18:@30323.4]
endmodule
module x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1( // @[:@30326.2]
  input         clock, // @[:@30327.4]
  input         reset, // @[:@30328.4]
  input         io_in_x529_ready, // @[:@30329.4]
  output        io_in_x529_valid, // @[:@30329.4]
  output [63:0] io_in_x529_bits_addr, // @[:@30329.4]
  output [31:0] io_in_x529_bits_size, // @[:@30329.4]
  input         io_in_x530_ready, // @[:@30329.4]
  output        io_in_x530_valid, // @[:@30329.4]
  output [7:0]  io_in_x530_bits_wdata_0, // @[:@30329.4]
  output        io_in_x530_bits_wstrb, // @[:@30329.4]
  output [20:0] io_in_x350_outbuf_0_rPort_0_ofs_0, // @[:@30329.4]
  output        io_in_x350_outbuf_0_rPort_0_en_0, // @[:@30329.4]
  output        io_in_x350_outbuf_0_rPort_0_backpressure, // @[:@30329.4]
  input  [7:0]  io_in_x350_outbuf_0_rPort_0_output_0, // @[:@30329.4]
  output        io_in_x531_ready, // @[:@30329.4]
  input         io_in_x531_valid, // @[:@30329.4]
  input  [63:0] io_in_x346_outdram_number, // @[:@30329.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@30329.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@30329.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@30329.4]
  input         io_sigsIn_smChildAcks_0, // @[:@30329.4]
  input         io_sigsIn_smChildAcks_1, // @[:@30329.4]
  input         io_sigsIn_smChildAcks_2, // @[:@30329.4]
  output        io_sigsOut_smDoneIn_0, // @[:@30329.4]
  output        io_sigsOut_smDoneIn_1, // @[:@30329.4]
  output        io_sigsOut_smDoneIn_2, // @[:@30329.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@30329.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@30329.4]
  output        io_sigsOut_smCtrCopyDone_2, // @[:@30329.4]
  input         io_rr // @[:@30329.4]
);
  wire  x536_inr_UnitPipe_sm_clock; // @[sm_x536_inr_UnitPipe.scala 33:18:@30396.4]
  wire  x536_inr_UnitPipe_sm_reset; // @[sm_x536_inr_UnitPipe.scala 33:18:@30396.4]
  wire  x536_inr_UnitPipe_sm_io_enable; // @[sm_x536_inr_UnitPipe.scala 33:18:@30396.4]
  wire  x536_inr_UnitPipe_sm_io_done; // @[sm_x536_inr_UnitPipe.scala 33:18:@30396.4]
  wire  x536_inr_UnitPipe_sm_io_doneLatch; // @[sm_x536_inr_UnitPipe.scala 33:18:@30396.4]
  wire  x536_inr_UnitPipe_sm_io_ctrDone; // @[sm_x536_inr_UnitPipe.scala 33:18:@30396.4]
  wire  x536_inr_UnitPipe_sm_io_datapathEn; // @[sm_x536_inr_UnitPipe.scala 33:18:@30396.4]
  wire  x536_inr_UnitPipe_sm_io_ctrInc; // @[sm_x536_inr_UnitPipe.scala 33:18:@30396.4]
  wire  x536_inr_UnitPipe_sm_io_parentAck; // @[sm_x536_inr_UnitPipe.scala 33:18:@30396.4]
  wire  x536_inr_UnitPipe_sm_io_backpressure; // @[sm_x536_inr_UnitPipe.scala 33:18:@30396.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@30453.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@30453.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@30453.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@30453.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@30453.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@30461.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@30461.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@30461.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@30461.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@30461.4]
  wire  x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_in_x529_valid; // @[sm_x536_inr_UnitPipe.scala 69:24:@30491.4]
  wire [63:0] x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_in_x529_bits_addr; // @[sm_x536_inr_UnitPipe.scala 69:24:@30491.4]
  wire [31:0] x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_in_x529_bits_size; // @[sm_x536_inr_UnitPipe.scala 69:24:@30491.4]
  wire [63:0] x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_in_x346_outdram_number; // @[sm_x536_inr_UnitPipe.scala 69:24:@30491.4]
  wire  x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x536_inr_UnitPipe.scala 69:24:@30491.4]
  wire  x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x536_inr_UnitPipe.scala 69:24:@30491.4]
  wire  x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_rr; // @[sm_x536_inr_UnitPipe.scala 69:24:@30491.4]
  wire  x538_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@30559.4]
  wire  x538_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@30559.4]
  wire  x538_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@30559.4]
  wire  x538_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@30559.4]
  wire [22:0] x538_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@30559.4]
  wire  x538_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@30559.4]
  wire  x538_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@30559.4]
  wire  x545_inr_Foreach_sm_clock; // @[sm_x545_inr_Foreach.scala 33:18:@30612.4]
  wire  x545_inr_Foreach_sm_reset; // @[sm_x545_inr_Foreach.scala 33:18:@30612.4]
  wire  x545_inr_Foreach_sm_io_enable; // @[sm_x545_inr_Foreach.scala 33:18:@30612.4]
  wire  x545_inr_Foreach_sm_io_done; // @[sm_x545_inr_Foreach.scala 33:18:@30612.4]
  wire  x545_inr_Foreach_sm_io_doneLatch; // @[sm_x545_inr_Foreach.scala 33:18:@30612.4]
  wire  x545_inr_Foreach_sm_io_ctrDone; // @[sm_x545_inr_Foreach.scala 33:18:@30612.4]
  wire  x545_inr_Foreach_sm_io_datapathEn; // @[sm_x545_inr_Foreach.scala 33:18:@30612.4]
  wire  x545_inr_Foreach_sm_io_ctrInc; // @[sm_x545_inr_Foreach.scala 33:18:@30612.4]
  wire  x545_inr_Foreach_sm_io_ctrRst; // @[sm_x545_inr_Foreach.scala 33:18:@30612.4]
  wire  x545_inr_Foreach_sm_io_parentAck; // @[sm_x545_inr_Foreach.scala 33:18:@30612.4]
  wire  x545_inr_Foreach_sm_io_backpressure; // @[sm_x545_inr_Foreach.scala 33:18:@30612.4]
  wire  x545_inr_Foreach_sm_io_break; // @[sm_x545_inr_Foreach.scala 33:18:@30612.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@30640.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@30640.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@30640.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@30640.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@30640.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@30680.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@30680.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@30680.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@30680.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@30680.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@30688.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@30688.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@30688.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@30688.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@30688.4]
  wire  x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_clock; // @[sm_x545_inr_Foreach.scala 78:24:@30723.4]
  wire  x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_reset; // @[sm_x545_inr_Foreach.scala 78:24:@30723.4]
  wire  x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x530_valid; // @[sm_x545_inr_Foreach.scala 78:24:@30723.4]
  wire [7:0] x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x530_bits_wdata_0; // @[sm_x545_inr_Foreach.scala 78:24:@30723.4]
  wire  x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x530_bits_wstrb; // @[sm_x545_inr_Foreach.scala 78:24:@30723.4]
  wire [20:0] x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x350_outbuf_0_rPort_0_ofs_0; // @[sm_x545_inr_Foreach.scala 78:24:@30723.4]
  wire  x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x350_outbuf_0_rPort_0_en_0; // @[sm_x545_inr_Foreach.scala 78:24:@30723.4]
  wire  x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x350_outbuf_0_rPort_0_backpressure; // @[sm_x545_inr_Foreach.scala 78:24:@30723.4]
  wire [7:0] x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x350_outbuf_0_rPort_0_output_0; // @[sm_x545_inr_Foreach.scala 78:24:@30723.4]
  wire  x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x545_inr_Foreach.scala 78:24:@30723.4]
  wire  x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x545_inr_Foreach.scala 78:24:@30723.4]
  wire  x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x545_inr_Foreach.scala 78:24:@30723.4]
  wire [31:0] x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x545_inr_Foreach.scala 78:24:@30723.4]
  wire  x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x545_inr_Foreach.scala 78:24:@30723.4]
  wire  x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_rr; // @[sm_x545_inr_Foreach.scala 78:24:@30723.4]
  wire  x549_inr_UnitPipe_sm_clock; // @[sm_x549_inr_UnitPipe.scala 32:18:@30843.4]
  wire  x549_inr_UnitPipe_sm_reset; // @[sm_x549_inr_UnitPipe.scala 32:18:@30843.4]
  wire  x549_inr_UnitPipe_sm_io_enable; // @[sm_x549_inr_UnitPipe.scala 32:18:@30843.4]
  wire  x549_inr_UnitPipe_sm_io_done; // @[sm_x549_inr_UnitPipe.scala 32:18:@30843.4]
  wire  x549_inr_UnitPipe_sm_io_doneLatch; // @[sm_x549_inr_UnitPipe.scala 32:18:@30843.4]
  wire  x549_inr_UnitPipe_sm_io_ctrDone; // @[sm_x549_inr_UnitPipe.scala 32:18:@30843.4]
  wire  x549_inr_UnitPipe_sm_io_datapathEn; // @[sm_x549_inr_UnitPipe.scala 32:18:@30843.4]
  wire  x549_inr_UnitPipe_sm_io_ctrInc; // @[sm_x549_inr_UnitPipe.scala 32:18:@30843.4]
  wire  x549_inr_UnitPipe_sm_io_parentAck; // @[sm_x549_inr_UnitPipe.scala 32:18:@30843.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@30900.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@30900.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@30900.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@30900.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@30900.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@30908.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@30908.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@30908.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@30908.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@30908.4]
  wire  x549_inr_UnitPipe_kernelx549_inr_UnitPipe_concrete1_io_in_x531_ready; // @[sm_x549_inr_UnitPipe.scala 60:24:@30938.4]
  wire  x549_inr_UnitPipe_kernelx549_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x549_inr_UnitPipe.scala 60:24:@30938.4]
  wire  _T_359; // @[package.scala 100:49:@30424.4]
  reg  _T_362; // @[package.scala 48:56:@30425.4]
  reg [31:0] _RAND_0;
  wire  _T_375; // @[package.scala 96:25:@30458.4 package.scala 96:25:@30459.4]
  wire  _T_381; // @[package.scala 96:25:@30466.4 package.scala 96:25:@30467.4]
  wire  _T_384; // @[SpatialBlocks.scala 138:93:@30469.4]
  wire  _T_454; // @[package.scala 96:25:@30645.4 package.scala 96:25:@30646.4]
  wire  _T_468; // @[package.scala 96:25:@30685.4 package.scala 96:25:@30686.4]
  wire  _T_474; // @[package.scala 96:25:@30693.4 package.scala 96:25:@30694.4]
  wire  _T_477; // @[SpatialBlocks.scala 138:93:@30696.4]
  wire  _T_479; // @[SpatialBlocks.scala 157:36:@30705.4]
  wire  _T_480; // @[SpatialBlocks.scala 157:78:@30706.4]
  wire  _T_547; // @[package.scala 100:49:@30871.4]
  reg  _T_550; // @[package.scala 48:56:@30872.4]
  reg [31:0] _RAND_1;
  wire  x549_inr_UnitPipe_sigsIn_forwardpressure; // @[sm_x550_outr_UnitPipe.scala 101:55:@30878.4]
  wire  _T_563; // @[package.scala 96:25:@30905.4 package.scala 96:25:@30906.4]
  wire  _T_569; // @[package.scala 96:25:@30913.4 package.scala 96:25:@30914.4]
  wire  _T_572; // @[SpatialBlocks.scala 138:93:@30916.4]
  wire  x549_inr_UnitPipe_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@30917.4]
  x536_inr_UnitPipe_sm x536_inr_UnitPipe_sm ( // @[sm_x536_inr_UnitPipe.scala 33:18:@30396.4]
    .clock(x536_inr_UnitPipe_sm_clock),
    .reset(x536_inr_UnitPipe_sm_reset),
    .io_enable(x536_inr_UnitPipe_sm_io_enable),
    .io_done(x536_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x536_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x536_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x536_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x536_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x536_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x536_inr_UnitPipe_sm_io_backpressure)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@30453.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@30461.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1 x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1 ( // @[sm_x536_inr_UnitPipe.scala 69:24:@30491.4]
    .io_in_x529_valid(x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_in_x529_valid),
    .io_in_x529_bits_addr(x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_in_x529_bits_addr),
    .io_in_x529_bits_size(x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_in_x529_bits_size),
    .io_in_x346_outdram_number(x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_in_x346_outdram_number),
    .io_sigsIn_backpressure(x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_rr(x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_rr)
  );
  x538_ctrchain x538_ctrchain ( // @[SpatialBlocks.scala 37:22:@30559.4]
    .clock(x538_ctrchain_clock),
    .reset(x538_ctrchain_reset),
    .io_input_reset(x538_ctrchain_io_input_reset),
    .io_input_enable(x538_ctrchain_io_input_enable),
    .io_output_counts_0(x538_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x538_ctrchain_io_output_oobs_0),
    .io_output_done(x538_ctrchain_io_output_done)
  );
  x545_inr_Foreach_sm x545_inr_Foreach_sm ( // @[sm_x545_inr_Foreach.scala 33:18:@30612.4]
    .clock(x545_inr_Foreach_sm_clock),
    .reset(x545_inr_Foreach_sm_reset),
    .io_enable(x545_inr_Foreach_sm_io_enable),
    .io_done(x545_inr_Foreach_sm_io_done),
    .io_doneLatch(x545_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x545_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x545_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x545_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x545_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x545_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x545_inr_Foreach_sm_io_backpressure),
    .io_break(x545_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@30640.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@30680.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@30688.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x545_inr_Foreach_kernelx545_inr_Foreach_concrete1 x545_inr_Foreach_kernelx545_inr_Foreach_concrete1 ( // @[sm_x545_inr_Foreach.scala 78:24:@30723.4]
    .clock(x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_clock),
    .reset(x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_reset),
    .io_in_x530_valid(x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x530_valid),
    .io_in_x530_bits_wdata_0(x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x530_bits_wdata_0),
    .io_in_x530_bits_wstrb(x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x530_bits_wstrb),
    .io_in_x350_outbuf_0_rPort_0_ofs_0(x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x350_outbuf_0_rPort_0_ofs_0),
    .io_in_x350_outbuf_0_rPort_0_en_0(x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x350_outbuf_0_rPort_0_en_0),
    .io_in_x350_outbuf_0_rPort_0_backpressure(x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x350_outbuf_0_rPort_0_backpressure),
    .io_in_x350_outbuf_0_rPort_0_output_0(x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x350_outbuf_0_rPort_0_output_0),
    .io_sigsIn_backpressure(x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_rr)
  );
  x549_inr_UnitPipe_sm x549_inr_UnitPipe_sm ( // @[sm_x549_inr_UnitPipe.scala 32:18:@30843.4]
    .clock(x549_inr_UnitPipe_sm_clock),
    .reset(x549_inr_UnitPipe_sm_reset),
    .io_enable(x549_inr_UnitPipe_sm_io_enable),
    .io_done(x549_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x549_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x549_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x549_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x549_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x549_inr_UnitPipe_sm_io_parentAck)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@30900.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@30908.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x549_inr_UnitPipe_kernelx549_inr_UnitPipe_concrete1 x549_inr_UnitPipe_kernelx549_inr_UnitPipe_concrete1 ( // @[sm_x549_inr_UnitPipe.scala 60:24:@30938.4]
    .io_in_x531_ready(x549_inr_UnitPipe_kernelx549_inr_UnitPipe_concrete1_io_in_x531_ready),
    .io_sigsIn_datapathEn(x549_inr_UnitPipe_kernelx549_inr_UnitPipe_concrete1_io_sigsIn_datapathEn)
  );
  assign _T_359 = x536_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@30424.4]
  assign _T_375 = RetimeWrapper_io_out; // @[package.scala 96:25:@30458.4 package.scala 96:25:@30459.4]
  assign _T_381 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@30466.4 package.scala 96:25:@30467.4]
  assign _T_384 = ~ _T_381; // @[SpatialBlocks.scala 138:93:@30469.4]
  assign _T_454 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@30645.4 package.scala 96:25:@30646.4]
  assign _T_468 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@30685.4 package.scala 96:25:@30686.4]
  assign _T_474 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@30693.4 package.scala 96:25:@30694.4]
  assign _T_477 = ~ _T_474; // @[SpatialBlocks.scala 138:93:@30696.4]
  assign _T_479 = x545_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@30705.4]
  assign _T_480 = ~ x545_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@30706.4]
  assign _T_547 = x549_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@30871.4]
  assign x549_inr_UnitPipe_sigsIn_forwardpressure = io_in_x531_valid | x549_inr_UnitPipe_sm_io_doneLatch; // @[sm_x550_outr_UnitPipe.scala 101:55:@30878.4]
  assign _T_563 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@30905.4 package.scala 96:25:@30906.4]
  assign _T_569 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@30913.4 package.scala 96:25:@30914.4]
  assign _T_572 = ~ _T_569; // @[SpatialBlocks.scala 138:93:@30916.4]
  assign x549_inr_UnitPipe_sigsIn_baseEn = _T_563 & _T_572; // @[SpatialBlocks.scala 138:90:@30917.4]
  assign io_in_x529_valid = x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_in_x529_valid; // @[sm_x536_inr_UnitPipe.scala 49:23:@30529.4]
  assign io_in_x529_bits_addr = x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_in_x529_bits_addr; // @[sm_x536_inr_UnitPipe.scala 49:23:@30528.4]
  assign io_in_x529_bits_size = x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_in_x529_bits_size; // @[sm_x536_inr_UnitPipe.scala 49:23:@30527.4]
  assign io_in_x530_valid = x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x530_valid; // @[sm_x545_inr_Foreach.scala 49:23:@30773.4]
  assign io_in_x530_bits_wdata_0 = x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x530_bits_wdata_0; // @[sm_x545_inr_Foreach.scala 49:23:@30772.4]
  assign io_in_x530_bits_wstrb = x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x530_bits_wstrb; // @[sm_x545_inr_Foreach.scala 49:23:@30771.4]
  assign io_in_x350_outbuf_0_rPort_0_ofs_0 = x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x350_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@30778.4]
  assign io_in_x350_outbuf_0_rPort_0_en_0 = x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x350_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@30777.4]
  assign io_in_x350_outbuf_0_rPort_0_backpressure = x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x350_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@30776.4]
  assign io_in_x531_ready = x549_inr_UnitPipe_kernelx549_inr_UnitPipe_concrete1_io_in_x531_ready; // @[sm_x549_inr_UnitPipe.scala 46:23:@30974.4]
  assign io_sigsOut_smDoneIn_0 = x536_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@30476.4]
  assign io_sigsOut_smDoneIn_1 = x545_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@30703.4]
  assign io_sigsOut_smDoneIn_2 = x549_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@30923.4]
  assign io_sigsOut_smCtrCopyDone_0 = x536_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@30490.4]
  assign io_sigsOut_smCtrCopyDone_1 = x545_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@30722.4]
  assign io_sigsOut_smCtrCopyDone_2 = x549_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@30937.4]
  assign x536_inr_UnitPipe_sm_clock = clock; // @[:@30397.4]
  assign x536_inr_UnitPipe_sm_reset = reset; // @[:@30398.4]
  assign x536_inr_UnitPipe_sm_io_enable = _T_375 & _T_384; // @[SpatialBlocks.scala 140:18:@30473.4]
  assign x536_inr_UnitPipe_sm_io_ctrDone = x536_inr_UnitPipe_sm_io_ctrInc & _T_362; // @[sm_x550_outr_UnitPipe.scala 77:39:@30428.4]
  assign x536_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@30475.4]
  assign x536_inr_UnitPipe_sm_io_backpressure = io_in_x529_ready | x536_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@30447.4]
  assign RetimeWrapper_clock = clock; // @[:@30454.4]
  assign RetimeWrapper_reset = reset; // @[:@30455.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@30457.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@30456.4]
  assign RetimeWrapper_1_clock = clock; // @[:@30462.4]
  assign RetimeWrapper_1_reset = reset; // @[:@30463.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@30465.4]
  assign RetimeWrapper_1_io_in = x536_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@30464.4]
  assign x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_in_x346_outdram_number = io_in_x346_outdram_number; // @[sm_x536_inr_UnitPipe.scala 50:31:@30531.4]
  assign x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x529_ready | x536_inr_UnitPipe_sm_io_doneLatch; // @[sm_x536_inr_UnitPipe.scala 74:22:@30546.4]
  assign x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x536_inr_UnitPipe_sm_io_datapathEn; // @[sm_x536_inr_UnitPipe.scala 74:22:@30544.4]
  assign x536_inr_UnitPipe_kernelx536_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x536_inr_UnitPipe.scala 73:18:@30532.4]
  assign x538_ctrchain_clock = clock; // @[:@30560.4]
  assign x538_ctrchain_reset = reset; // @[:@30561.4]
  assign x538_ctrchain_io_input_reset = x545_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@30721.4]
  assign x538_ctrchain_io_input_enable = x545_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@30673.4 SpatialBlocks.scala 159:42:@30720.4]
  assign x545_inr_Foreach_sm_clock = clock; // @[:@30613.4]
  assign x545_inr_Foreach_sm_reset = reset; // @[:@30614.4]
  assign x545_inr_Foreach_sm_io_enable = _T_468 & _T_477; // @[SpatialBlocks.scala 140:18:@30700.4]
  assign x545_inr_Foreach_sm_io_ctrDone = io_rr ? _T_454 : 1'h0; // @[sm_x550_outr_UnitPipe.scala 90:38:@30648.4]
  assign x545_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@30702.4]
  assign x545_inr_Foreach_sm_io_backpressure = io_in_x530_ready | x545_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@30674.4]
  assign x545_inr_Foreach_sm_io_break = 1'h0; // @[sm_x550_outr_UnitPipe.scala 94:36:@30654.4]
  assign RetimeWrapper_2_clock = clock; // @[:@30641.4]
  assign RetimeWrapper_2_reset = reset; // @[:@30642.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@30644.4]
  assign RetimeWrapper_2_io_in = x538_ctrchain_io_output_done; // @[package.scala 94:16:@30643.4]
  assign RetimeWrapper_3_clock = clock; // @[:@30681.4]
  assign RetimeWrapper_3_reset = reset; // @[:@30682.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@30684.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@30683.4]
  assign RetimeWrapper_4_clock = clock; // @[:@30689.4]
  assign RetimeWrapper_4_reset = reset; // @[:@30690.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@30692.4]
  assign RetimeWrapper_4_io_in = x545_inr_Foreach_sm_io_done; // @[package.scala 94:16:@30691.4]
  assign x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_clock = clock; // @[:@30724.4]
  assign x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_reset = reset; // @[:@30725.4]
  assign x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_in_x350_outbuf_0_rPort_0_output_0 = io_in_x350_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@30775.4]
  assign x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x530_ready | x545_inr_Foreach_sm_io_doneLatch; // @[sm_x545_inr_Foreach.scala 83:22:@30794.4]
  assign x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_479 & _T_480; // @[sm_x545_inr_Foreach.scala 83:22:@30792.4]
  assign x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_sigsIn_break = x545_inr_Foreach_sm_io_break; // @[sm_x545_inr_Foreach.scala 83:22:@30790.4]
  assign x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{9{x538_ctrchain_io_output_counts_0[22]}},x538_ctrchain_io_output_counts_0}; // @[sm_x545_inr_Foreach.scala 83:22:@30785.4]
  assign x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x538_ctrchain_io_output_oobs_0; // @[sm_x545_inr_Foreach.scala 83:22:@30784.4]
  assign x545_inr_Foreach_kernelx545_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x545_inr_Foreach.scala 82:18:@30780.4]
  assign x549_inr_UnitPipe_sm_clock = clock; // @[:@30844.4]
  assign x549_inr_UnitPipe_sm_reset = reset; // @[:@30845.4]
  assign x549_inr_UnitPipe_sm_io_enable = x549_inr_UnitPipe_sigsIn_baseEn & x549_inr_UnitPipe_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@30920.4]
  assign x549_inr_UnitPipe_sm_io_ctrDone = x549_inr_UnitPipe_sm_io_ctrInc & _T_550; // @[sm_x550_outr_UnitPipe.scala 99:39:@30875.4]
  assign x549_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 142:21:@30922.4]
  assign RetimeWrapper_5_clock = clock; // @[:@30901.4]
  assign RetimeWrapper_5_reset = reset; // @[:@30902.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@30904.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@30903.4]
  assign RetimeWrapper_6_clock = clock; // @[:@30909.4]
  assign RetimeWrapper_6_reset = reset; // @[:@30910.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@30912.4]
  assign RetimeWrapper_6_io_in = x549_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@30911.4]
  assign x549_inr_UnitPipe_kernelx549_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x549_inr_UnitPipe_sm_io_datapathEn; // @[sm_x549_inr_UnitPipe.scala 65:22:@30987.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_362 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_550 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_362 <= 1'h0;
    end else begin
      _T_362 <= _T_359;
    end
    if (reset) begin
      _T_550 <= 1'h0;
    end else begin
      _T_550 <= _T_547;
    end
  end
endmodule
module x607_kernelx607_concrete1( // @[:@31003.2]
  input          clock, // @[:@31004.4]
  input          reset, // @[:@31005.4]
  input          io_in_x348_TVALID, // @[:@31006.4]
  output         io_in_x348_TREADY, // @[:@31006.4]
  input  [255:0] io_in_x348_TDATA, // @[:@31006.4]
  input  [7:0]   io_in_x348_TID, // @[:@31006.4]
  input  [7:0]   io_in_x348_TDEST, // @[:@31006.4]
  input          io_in_x529_ready, // @[:@31006.4]
  output         io_in_x529_valid, // @[:@31006.4]
  output [63:0]  io_in_x529_bits_addr, // @[:@31006.4]
  output [31:0]  io_in_x529_bits_size, // @[:@31006.4]
  output         io_in_x349_TVALID, // @[:@31006.4]
  input          io_in_x349_TREADY, // @[:@31006.4]
  output [255:0] io_in_x349_TDATA, // @[:@31006.4]
  input          io_in_x530_ready, // @[:@31006.4]
  output         io_in_x530_valid, // @[:@31006.4]
  output [7:0]   io_in_x530_bits_wdata_0, // @[:@31006.4]
  output         io_in_x530_bits_wstrb, // @[:@31006.4]
  output [20:0]  io_in_x350_outbuf_0_rPort_0_ofs_0, // @[:@31006.4]
  output         io_in_x350_outbuf_0_rPort_0_en_0, // @[:@31006.4]
  output         io_in_x350_outbuf_0_rPort_0_backpressure, // @[:@31006.4]
  input  [7:0]   io_in_x350_outbuf_0_rPort_0_output_0, // @[:@31006.4]
  output         io_in_x531_ready, // @[:@31006.4]
  input          io_in_x531_valid, // @[:@31006.4]
  input  [63:0]  io_in_x346_outdram_number, // @[:@31006.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@31006.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@31006.4]
  input          io_sigsIn_smChildAcks_0, // @[:@31006.4]
  input          io_sigsIn_smChildAcks_1, // @[:@31006.4]
  output         io_sigsOut_smDoneIn_0, // @[:@31006.4]
  output         io_sigsOut_smDoneIn_1, // @[:@31006.4]
  input          io_rr // @[:@31006.4]
);
  wire  x528_outr_UnitPipe_sm_clock; // @[sm_x528_outr_UnitPipe.scala 32:18:@31079.4]
  wire  x528_outr_UnitPipe_sm_reset; // @[sm_x528_outr_UnitPipe.scala 32:18:@31079.4]
  wire  x528_outr_UnitPipe_sm_io_enable; // @[sm_x528_outr_UnitPipe.scala 32:18:@31079.4]
  wire  x528_outr_UnitPipe_sm_io_done; // @[sm_x528_outr_UnitPipe.scala 32:18:@31079.4]
  wire  x528_outr_UnitPipe_sm_io_parentAck; // @[sm_x528_outr_UnitPipe.scala 32:18:@31079.4]
  wire  x528_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x528_outr_UnitPipe.scala 32:18:@31079.4]
  wire  x528_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x528_outr_UnitPipe.scala 32:18:@31079.4]
  wire  x528_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x528_outr_UnitPipe.scala 32:18:@31079.4]
  wire  x528_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x528_outr_UnitPipe.scala 32:18:@31079.4]
  wire  x528_outr_UnitPipe_sm_io_childAck_0; // @[sm_x528_outr_UnitPipe.scala 32:18:@31079.4]
  wire  x528_outr_UnitPipe_sm_io_childAck_1; // @[sm_x528_outr_UnitPipe.scala 32:18:@31079.4]
  wire  x528_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x528_outr_UnitPipe.scala 32:18:@31079.4]
  wire  x528_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x528_outr_UnitPipe.scala 32:18:@31079.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@31141.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@31141.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@31141.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@31141.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@31141.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@31149.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@31149.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@31149.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@31149.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@31149.4]
  wire  x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_clock; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire  x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_reset; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire  x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x348_TVALID; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire  x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x348_TREADY; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire [255:0] x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x348_TDATA; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire [7:0] x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x348_TID; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire [7:0] x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x348_TDEST; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire  x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x349_TVALID; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire  x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x349_TREADY; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire [255:0] x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x349_TDATA; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire  x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire  x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire  x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire  x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire  x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire  x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire  x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire  x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire  x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_rr; // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
  wire  x550_outr_UnitPipe_sm_clock; // @[sm_x550_outr_UnitPipe.scala 36:18:@31358.4]
  wire  x550_outr_UnitPipe_sm_reset; // @[sm_x550_outr_UnitPipe.scala 36:18:@31358.4]
  wire  x550_outr_UnitPipe_sm_io_enable; // @[sm_x550_outr_UnitPipe.scala 36:18:@31358.4]
  wire  x550_outr_UnitPipe_sm_io_done; // @[sm_x550_outr_UnitPipe.scala 36:18:@31358.4]
  wire  x550_outr_UnitPipe_sm_io_parentAck; // @[sm_x550_outr_UnitPipe.scala 36:18:@31358.4]
  wire  x550_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x550_outr_UnitPipe.scala 36:18:@31358.4]
  wire  x550_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x550_outr_UnitPipe.scala 36:18:@31358.4]
  wire  x550_outr_UnitPipe_sm_io_doneIn_2; // @[sm_x550_outr_UnitPipe.scala 36:18:@31358.4]
  wire  x550_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x550_outr_UnitPipe.scala 36:18:@31358.4]
  wire  x550_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x550_outr_UnitPipe.scala 36:18:@31358.4]
  wire  x550_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x550_outr_UnitPipe.scala 36:18:@31358.4]
  wire  x550_outr_UnitPipe_sm_io_childAck_0; // @[sm_x550_outr_UnitPipe.scala 36:18:@31358.4]
  wire  x550_outr_UnitPipe_sm_io_childAck_1; // @[sm_x550_outr_UnitPipe.scala 36:18:@31358.4]
  wire  x550_outr_UnitPipe_sm_io_childAck_2; // @[sm_x550_outr_UnitPipe.scala 36:18:@31358.4]
  wire  x550_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x550_outr_UnitPipe.scala 36:18:@31358.4]
  wire  x550_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x550_outr_UnitPipe.scala 36:18:@31358.4]
  wire  x550_outr_UnitPipe_sm_io_ctrCopyDone_2; // @[sm_x550_outr_UnitPipe.scala 36:18:@31358.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@31430.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@31430.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@31430.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@31430.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@31430.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@31438.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@31438.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@31438.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@31438.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@31438.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_clock; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_reset; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x529_ready; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x529_valid; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire [63:0] x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x529_bits_addr; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire [31:0] x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x529_bits_size; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x530_ready; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x530_valid; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire [7:0] x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x530_bits_wdata_0; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x530_bits_wstrb; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire [20:0] x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x350_outbuf_0_rPort_0_ofs_0; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x350_outbuf_0_rPort_0_en_0; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x350_outbuf_0_rPort_0_backpressure; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire [7:0] x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x350_outbuf_0_rPort_0_output_0; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x531_ready; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x531_valid; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire [63:0] x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x346_outdram_number; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_rr; // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
  wire  _T_408; // @[package.scala 96:25:@31146.4 package.scala 96:25:@31147.4]
  wire  _T_414; // @[package.scala 96:25:@31154.4 package.scala 96:25:@31155.4]
  wire  _T_417; // @[SpatialBlocks.scala 138:93:@31157.4]
  wire  _T_508; // @[package.scala 96:25:@31435.4 package.scala 96:25:@31436.4]
  wire  _T_514; // @[package.scala 96:25:@31443.4 package.scala 96:25:@31444.4]
  wire  _T_517; // @[SpatialBlocks.scala 138:93:@31446.4]
  x528_outr_UnitPipe_sm x528_outr_UnitPipe_sm ( // @[sm_x528_outr_UnitPipe.scala 32:18:@31079.4]
    .clock(x528_outr_UnitPipe_sm_clock),
    .reset(x528_outr_UnitPipe_sm_reset),
    .io_enable(x528_outr_UnitPipe_sm_io_enable),
    .io_done(x528_outr_UnitPipe_sm_io_done),
    .io_parentAck(x528_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x528_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x528_outr_UnitPipe_sm_io_doneIn_1),
    .io_enableOut_0(x528_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x528_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x528_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x528_outr_UnitPipe_sm_io_childAck_1),
    .io_ctrCopyDone_0(x528_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x528_outr_UnitPipe_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@31141.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@31149.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1 x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1 ( // @[sm_x528_outr_UnitPipe.scala 87:24:@31180.4]
    .clock(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_clock),
    .reset(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_reset),
    .io_in_x348_TVALID(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x348_TVALID),
    .io_in_x348_TREADY(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x348_TREADY),
    .io_in_x348_TDATA(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x348_TDATA),
    .io_in_x348_TID(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x348_TID),
    .io_in_x348_TDEST(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x348_TDEST),
    .io_in_x349_TVALID(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x349_TVALID),
    .io_in_x349_TREADY(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x349_TREADY),
    .io_in_x349_TDATA(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x349_TDATA),
    .io_sigsIn_smEnableOuts_0(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_rr)
  );
  x550_outr_UnitPipe_sm x550_outr_UnitPipe_sm ( // @[sm_x550_outr_UnitPipe.scala 36:18:@31358.4]
    .clock(x550_outr_UnitPipe_sm_clock),
    .reset(x550_outr_UnitPipe_sm_reset),
    .io_enable(x550_outr_UnitPipe_sm_io_enable),
    .io_done(x550_outr_UnitPipe_sm_io_done),
    .io_parentAck(x550_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x550_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x550_outr_UnitPipe_sm_io_doneIn_1),
    .io_doneIn_2(x550_outr_UnitPipe_sm_io_doneIn_2),
    .io_enableOut_0(x550_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x550_outr_UnitPipe_sm_io_enableOut_1),
    .io_enableOut_2(x550_outr_UnitPipe_sm_io_enableOut_2),
    .io_childAck_0(x550_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x550_outr_UnitPipe_sm_io_childAck_1),
    .io_childAck_2(x550_outr_UnitPipe_sm_io_childAck_2),
    .io_ctrCopyDone_0(x550_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x550_outr_UnitPipe_sm_io_ctrCopyDone_1),
    .io_ctrCopyDone_2(x550_outr_UnitPipe_sm_io_ctrCopyDone_2)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@31430.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@31438.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1 x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1 ( // @[sm_x550_outr_UnitPipe.scala 108:24:@31470.4]
    .clock(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_clock),
    .reset(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_reset),
    .io_in_x529_ready(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x529_ready),
    .io_in_x529_valid(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x529_valid),
    .io_in_x529_bits_addr(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x529_bits_addr),
    .io_in_x529_bits_size(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x529_bits_size),
    .io_in_x530_ready(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x530_ready),
    .io_in_x530_valid(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x530_valid),
    .io_in_x530_bits_wdata_0(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x530_bits_wdata_0),
    .io_in_x530_bits_wstrb(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x530_bits_wstrb),
    .io_in_x350_outbuf_0_rPort_0_ofs_0(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x350_outbuf_0_rPort_0_ofs_0),
    .io_in_x350_outbuf_0_rPort_0_en_0(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x350_outbuf_0_rPort_0_en_0),
    .io_in_x350_outbuf_0_rPort_0_backpressure(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x350_outbuf_0_rPort_0_backpressure),
    .io_in_x350_outbuf_0_rPort_0_output_0(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x350_outbuf_0_rPort_0_output_0),
    .io_in_x531_ready(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x531_ready),
    .io_in_x531_valid(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x531_valid),
    .io_in_x346_outdram_number(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x346_outdram_number),
    .io_sigsIn_smEnableOuts_0(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smCtrCopyDone_0(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_sigsOut_smCtrCopyDone_2(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2),
    .io_rr(x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_408 = RetimeWrapper_io_out; // @[package.scala 96:25:@31146.4 package.scala 96:25:@31147.4]
  assign _T_414 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@31154.4 package.scala 96:25:@31155.4]
  assign _T_417 = ~ _T_414; // @[SpatialBlocks.scala 138:93:@31157.4]
  assign _T_508 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@31435.4 package.scala 96:25:@31436.4]
  assign _T_514 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@31443.4 package.scala 96:25:@31444.4]
  assign _T_517 = ~ _T_514; // @[SpatialBlocks.scala 138:93:@31446.4]
  assign io_in_x348_TREADY = x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x348_TREADY; // @[sm_x528_outr_UnitPipe.scala 48:23:@31248.4]
  assign io_in_x529_valid = x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x529_valid; // @[sm_x550_outr_UnitPipe.scala 58:23:@31552.4]
  assign io_in_x529_bits_addr = x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x529_bits_addr; // @[sm_x550_outr_UnitPipe.scala 58:23:@31551.4]
  assign io_in_x529_bits_size = x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x529_bits_size; // @[sm_x550_outr_UnitPipe.scala 58:23:@31550.4]
  assign io_in_x349_TVALID = x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x349_TVALID; // @[sm_x528_outr_UnitPipe.scala 49:23:@31258.4]
  assign io_in_x349_TDATA = x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x349_TDATA; // @[sm_x528_outr_UnitPipe.scala 49:23:@31256.4]
  assign io_in_x530_valid = x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x530_valid; // @[sm_x550_outr_UnitPipe.scala 59:23:@31556.4]
  assign io_in_x530_bits_wdata_0 = x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x530_bits_wdata_0; // @[sm_x550_outr_UnitPipe.scala 59:23:@31555.4]
  assign io_in_x530_bits_wstrb = x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x530_bits_wstrb; // @[sm_x550_outr_UnitPipe.scala 59:23:@31554.4]
  assign io_in_x350_outbuf_0_rPort_0_ofs_0 = x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x350_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@31561.4]
  assign io_in_x350_outbuf_0_rPort_0_en_0 = x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x350_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@31560.4]
  assign io_in_x350_outbuf_0_rPort_0_backpressure = x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x350_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@31559.4]
  assign io_in_x531_ready = x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x531_ready; // @[sm_x550_outr_UnitPipe.scala 61:23:@31565.4]
  assign io_sigsOut_smDoneIn_0 = x528_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@31164.4]
  assign io_sigsOut_smDoneIn_1 = x550_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@31453.4]
  assign x528_outr_UnitPipe_sm_clock = clock; // @[:@31080.4]
  assign x528_outr_UnitPipe_sm_reset = reset; // @[:@31081.4]
  assign x528_outr_UnitPipe_sm_io_enable = _T_408 & _T_417; // @[SpatialBlocks.scala 140:18:@31161.4]
  assign x528_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@31163.4]
  assign x528_outr_UnitPipe_sm_io_doneIn_0 = x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@31131.4]
  assign x528_outr_UnitPipe_sm_io_doneIn_1 = x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@31132.4]
  assign x528_outr_UnitPipe_sm_io_ctrCopyDone_0 = x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@31178.4]
  assign x528_outr_UnitPipe_sm_io_ctrCopyDone_1 = x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@31179.4]
  assign RetimeWrapper_clock = clock; // @[:@31142.4]
  assign RetimeWrapper_reset = reset; // @[:@31143.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@31145.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@31144.4]
  assign RetimeWrapper_1_clock = clock; // @[:@31150.4]
  assign RetimeWrapper_1_reset = reset; // @[:@31151.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@31153.4]
  assign RetimeWrapper_1_io_in = x528_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@31152.4]
  assign x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_clock = clock; // @[:@31181.4]
  assign x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_reset = reset; // @[:@31182.4]
  assign x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x348_TVALID = io_in_x348_TVALID; // @[sm_x528_outr_UnitPipe.scala 48:23:@31249.4]
  assign x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x348_TDATA = io_in_x348_TDATA; // @[sm_x528_outr_UnitPipe.scala 48:23:@31247.4]
  assign x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x348_TID = io_in_x348_TID; // @[sm_x528_outr_UnitPipe.scala 48:23:@31243.4]
  assign x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x348_TDEST = io_in_x348_TDEST; // @[sm_x528_outr_UnitPipe.scala 48:23:@31242.4]
  assign x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_in_x349_TREADY = io_in_x349_TREADY; // @[sm_x528_outr_UnitPipe.scala 49:23:@31257.4]
  assign x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x528_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x528_outr_UnitPipe.scala 92:22:@31274.4]
  assign x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x528_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x528_outr_UnitPipe.scala 92:22:@31275.4]
  assign x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x528_outr_UnitPipe_sm_io_childAck_0; // @[sm_x528_outr_UnitPipe.scala 92:22:@31270.4]
  assign x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x528_outr_UnitPipe_sm_io_childAck_1; // @[sm_x528_outr_UnitPipe.scala 92:22:@31271.4]
  assign x528_outr_UnitPipe_kernelx528_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x528_outr_UnitPipe.scala 91:18:@31259.4]
  assign x550_outr_UnitPipe_sm_clock = clock; // @[:@31359.4]
  assign x550_outr_UnitPipe_sm_reset = reset; // @[:@31360.4]
  assign x550_outr_UnitPipe_sm_io_enable = _T_508 & _T_517; // @[SpatialBlocks.scala 140:18:@31450.4]
  assign x550_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@31452.4]
  assign x550_outr_UnitPipe_sm_io_doneIn_0 = x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@31418.4]
  assign x550_outr_UnitPipe_sm_io_doneIn_1 = x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@31419.4]
  assign x550_outr_UnitPipe_sm_io_doneIn_2 = x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:67:@31420.4]
  assign x550_outr_UnitPipe_sm_io_ctrCopyDone_0 = x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@31467.4]
  assign x550_outr_UnitPipe_sm_io_ctrCopyDone_1 = x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@31468.4]
  assign x550_outr_UnitPipe_sm_io_ctrCopyDone_2 = x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[SpatialBlocks.scala 161:90:@31469.4]
  assign RetimeWrapper_2_clock = clock; // @[:@31431.4]
  assign RetimeWrapper_2_reset = reset; // @[:@31432.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@31434.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@31433.4]
  assign RetimeWrapper_3_clock = clock; // @[:@31439.4]
  assign RetimeWrapper_3_reset = reset; // @[:@31440.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@31442.4]
  assign RetimeWrapper_3_io_in = x550_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@31441.4]
  assign x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_clock = clock; // @[:@31471.4]
  assign x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_reset = reset; // @[:@31472.4]
  assign x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x529_ready = io_in_x529_ready; // @[sm_x550_outr_UnitPipe.scala 58:23:@31553.4]
  assign x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x530_ready = io_in_x530_ready; // @[sm_x550_outr_UnitPipe.scala 59:23:@31557.4]
  assign x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x350_outbuf_0_rPort_0_output_0 = io_in_x350_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@31558.4]
  assign x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x531_valid = io_in_x531_valid; // @[sm_x550_outr_UnitPipe.scala 61:23:@31564.4]
  assign x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_in_x346_outdram_number = io_in_x346_outdram_number; // @[sm_x550_outr_UnitPipe.scala 62:31:@31566.4]
  assign x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x550_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x550_outr_UnitPipe.scala 113:22:@31589.4]
  assign x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x550_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x550_outr_UnitPipe.scala 113:22:@31590.4]
  assign x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2 = x550_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x550_outr_UnitPipe.scala 113:22:@31591.4]
  assign x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x550_outr_UnitPipe_sm_io_childAck_0; // @[sm_x550_outr_UnitPipe.scala 113:22:@31583.4]
  assign x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x550_outr_UnitPipe_sm_io_childAck_1; // @[sm_x550_outr_UnitPipe.scala 113:22:@31584.4]
  assign x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2 = x550_outr_UnitPipe_sm_io_childAck_2; // @[sm_x550_outr_UnitPipe.scala 113:22:@31585.4]
  assign x550_outr_UnitPipe_kernelx550_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x550_outr_UnitPipe.scala 112:18:@31567.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@31619.2]
  input          clock, // @[:@31620.4]
  input          reset, // @[:@31621.4]
  input          io_in_x348_TVALID, // @[:@31622.4]
  output         io_in_x348_TREADY, // @[:@31622.4]
  input  [255:0] io_in_x348_TDATA, // @[:@31622.4]
  input  [7:0]   io_in_x348_TID, // @[:@31622.4]
  input  [7:0]   io_in_x348_TDEST, // @[:@31622.4]
  input          io_in_x529_ready, // @[:@31622.4]
  output         io_in_x529_valid, // @[:@31622.4]
  output [63:0]  io_in_x529_bits_addr, // @[:@31622.4]
  output [31:0]  io_in_x529_bits_size, // @[:@31622.4]
  output         io_in_x349_TVALID, // @[:@31622.4]
  input          io_in_x349_TREADY, // @[:@31622.4]
  output [255:0] io_in_x349_TDATA, // @[:@31622.4]
  input          io_in_x530_ready, // @[:@31622.4]
  output         io_in_x530_valid, // @[:@31622.4]
  output [7:0]   io_in_x530_bits_wdata_0, // @[:@31622.4]
  output         io_in_x530_bits_wstrb, // @[:@31622.4]
  output         io_in_x531_ready, // @[:@31622.4]
  input          io_in_x531_valid, // @[:@31622.4]
  input  [63:0]  io_in_x346_outdram_number, // @[:@31622.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@31622.4]
  input          io_sigsIn_smChildAcks_0, // @[:@31622.4]
  output         io_sigsOut_smDoneIn_0, // @[:@31622.4]
  input          io_rr // @[:@31622.4]
);
  wire  x350_outbuf_0_clock; // @[m_x350_outbuf_0.scala 27:17:@31632.4]
  wire  x350_outbuf_0_reset; // @[m_x350_outbuf_0.scala 27:17:@31632.4]
  wire [20:0] x350_outbuf_0_io_rPort_0_ofs_0; // @[m_x350_outbuf_0.scala 27:17:@31632.4]
  wire  x350_outbuf_0_io_rPort_0_en_0; // @[m_x350_outbuf_0.scala 27:17:@31632.4]
  wire  x350_outbuf_0_io_rPort_0_backpressure; // @[m_x350_outbuf_0.scala 27:17:@31632.4]
  wire [7:0] x350_outbuf_0_io_rPort_0_output_0; // @[m_x350_outbuf_0.scala 27:17:@31632.4]
  wire  x607_sm_clock; // @[sm_x607.scala 37:18:@31690.4]
  wire  x607_sm_reset; // @[sm_x607.scala 37:18:@31690.4]
  wire  x607_sm_io_enable; // @[sm_x607.scala 37:18:@31690.4]
  wire  x607_sm_io_done; // @[sm_x607.scala 37:18:@31690.4]
  wire  x607_sm_io_ctrDone; // @[sm_x607.scala 37:18:@31690.4]
  wire  x607_sm_io_ctrInc; // @[sm_x607.scala 37:18:@31690.4]
  wire  x607_sm_io_parentAck; // @[sm_x607.scala 37:18:@31690.4]
  wire  x607_sm_io_doneIn_0; // @[sm_x607.scala 37:18:@31690.4]
  wire  x607_sm_io_doneIn_1; // @[sm_x607.scala 37:18:@31690.4]
  wire  x607_sm_io_enableOut_0; // @[sm_x607.scala 37:18:@31690.4]
  wire  x607_sm_io_enableOut_1; // @[sm_x607.scala 37:18:@31690.4]
  wire  x607_sm_io_childAck_0; // @[sm_x607.scala 37:18:@31690.4]
  wire  x607_sm_io_childAck_1; // @[sm_x607.scala 37:18:@31690.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@31757.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@31757.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@31757.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@31757.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@31757.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@31765.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@31765.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@31765.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@31765.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@31765.4]
  wire  x607_kernelx607_concrete1_clock; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_reset; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_in_x348_TVALID; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_in_x348_TREADY; // @[sm_x607.scala 102:24:@31794.4]
  wire [255:0] x607_kernelx607_concrete1_io_in_x348_TDATA; // @[sm_x607.scala 102:24:@31794.4]
  wire [7:0] x607_kernelx607_concrete1_io_in_x348_TID; // @[sm_x607.scala 102:24:@31794.4]
  wire [7:0] x607_kernelx607_concrete1_io_in_x348_TDEST; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_in_x529_ready; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_in_x529_valid; // @[sm_x607.scala 102:24:@31794.4]
  wire [63:0] x607_kernelx607_concrete1_io_in_x529_bits_addr; // @[sm_x607.scala 102:24:@31794.4]
  wire [31:0] x607_kernelx607_concrete1_io_in_x529_bits_size; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_in_x349_TVALID; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_in_x349_TREADY; // @[sm_x607.scala 102:24:@31794.4]
  wire [255:0] x607_kernelx607_concrete1_io_in_x349_TDATA; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_in_x530_ready; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_in_x530_valid; // @[sm_x607.scala 102:24:@31794.4]
  wire [7:0] x607_kernelx607_concrete1_io_in_x530_bits_wdata_0; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_in_x530_bits_wstrb; // @[sm_x607.scala 102:24:@31794.4]
  wire [20:0] x607_kernelx607_concrete1_io_in_x350_outbuf_0_rPort_0_ofs_0; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_in_x350_outbuf_0_rPort_0_en_0; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_in_x350_outbuf_0_rPort_0_backpressure; // @[sm_x607.scala 102:24:@31794.4]
  wire [7:0] x607_kernelx607_concrete1_io_in_x350_outbuf_0_rPort_0_output_0; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_in_x531_ready; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_in_x531_valid; // @[sm_x607.scala 102:24:@31794.4]
  wire [63:0] x607_kernelx607_concrete1_io_in_x346_outdram_number; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x607.scala 102:24:@31794.4]
  wire  x607_kernelx607_concrete1_io_rr; // @[sm_x607.scala 102:24:@31794.4]
  wire  _T_266; // @[package.scala 100:49:@31723.4]
  reg  _T_269; // @[package.scala 48:56:@31724.4]
  reg [31:0] _RAND_0;
  wire  _T_283; // @[package.scala 96:25:@31762.4 package.scala 96:25:@31763.4]
  wire  _T_289; // @[package.scala 96:25:@31770.4 package.scala 96:25:@31771.4]
  wire  _T_292; // @[SpatialBlocks.scala 138:93:@31773.4]
  x350_outbuf_0 x350_outbuf_0 ( // @[m_x350_outbuf_0.scala 27:17:@31632.4]
    .clock(x350_outbuf_0_clock),
    .reset(x350_outbuf_0_reset),
    .io_rPort_0_ofs_0(x350_outbuf_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x350_outbuf_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x350_outbuf_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x350_outbuf_0_io_rPort_0_output_0)
  );
  x607_sm x607_sm ( // @[sm_x607.scala 37:18:@31690.4]
    .clock(x607_sm_clock),
    .reset(x607_sm_reset),
    .io_enable(x607_sm_io_enable),
    .io_done(x607_sm_io_done),
    .io_ctrDone(x607_sm_io_ctrDone),
    .io_ctrInc(x607_sm_io_ctrInc),
    .io_parentAck(x607_sm_io_parentAck),
    .io_doneIn_0(x607_sm_io_doneIn_0),
    .io_doneIn_1(x607_sm_io_doneIn_1),
    .io_enableOut_0(x607_sm_io_enableOut_0),
    .io_enableOut_1(x607_sm_io_enableOut_1),
    .io_childAck_0(x607_sm_io_childAck_0),
    .io_childAck_1(x607_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@31757.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@31765.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x607_kernelx607_concrete1 x607_kernelx607_concrete1 ( // @[sm_x607.scala 102:24:@31794.4]
    .clock(x607_kernelx607_concrete1_clock),
    .reset(x607_kernelx607_concrete1_reset),
    .io_in_x348_TVALID(x607_kernelx607_concrete1_io_in_x348_TVALID),
    .io_in_x348_TREADY(x607_kernelx607_concrete1_io_in_x348_TREADY),
    .io_in_x348_TDATA(x607_kernelx607_concrete1_io_in_x348_TDATA),
    .io_in_x348_TID(x607_kernelx607_concrete1_io_in_x348_TID),
    .io_in_x348_TDEST(x607_kernelx607_concrete1_io_in_x348_TDEST),
    .io_in_x529_ready(x607_kernelx607_concrete1_io_in_x529_ready),
    .io_in_x529_valid(x607_kernelx607_concrete1_io_in_x529_valid),
    .io_in_x529_bits_addr(x607_kernelx607_concrete1_io_in_x529_bits_addr),
    .io_in_x529_bits_size(x607_kernelx607_concrete1_io_in_x529_bits_size),
    .io_in_x349_TVALID(x607_kernelx607_concrete1_io_in_x349_TVALID),
    .io_in_x349_TREADY(x607_kernelx607_concrete1_io_in_x349_TREADY),
    .io_in_x349_TDATA(x607_kernelx607_concrete1_io_in_x349_TDATA),
    .io_in_x530_ready(x607_kernelx607_concrete1_io_in_x530_ready),
    .io_in_x530_valid(x607_kernelx607_concrete1_io_in_x530_valid),
    .io_in_x530_bits_wdata_0(x607_kernelx607_concrete1_io_in_x530_bits_wdata_0),
    .io_in_x530_bits_wstrb(x607_kernelx607_concrete1_io_in_x530_bits_wstrb),
    .io_in_x350_outbuf_0_rPort_0_ofs_0(x607_kernelx607_concrete1_io_in_x350_outbuf_0_rPort_0_ofs_0),
    .io_in_x350_outbuf_0_rPort_0_en_0(x607_kernelx607_concrete1_io_in_x350_outbuf_0_rPort_0_en_0),
    .io_in_x350_outbuf_0_rPort_0_backpressure(x607_kernelx607_concrete1_io_in_x350_outbuf_0_rPort_0_backpressure),
    .io_in_x350_outbuf_0_rPort_0_output_0(x607_kernelx607_concrete1_io_in_x350_outbuf_0_rPort_0_output_0),
    .io_in_x531_ready(x607_kernelx607_concrete1_io_in_x531_ready),
    .io_in_x531_valid(x607_kernelx607_concrete1_io_in_x531_valid),
    .io_in_x346_outdram_number(x607_kernelx607_concrete1_io_in_x346_outdram_number),
    .io_sigsIn_smEnableOuts_0(x607_kernelx607_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x607_kernelx607_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x607_kernelx607_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x607_kernelx607_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x607_kernelx607_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x607_kernelx607_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(x607_kernelx607_concrete1_io_rr)
  );
  assign _T_266 = x607_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@31723.4]
  assign _T_283 = RetimeWrapper_io_out; // @[package.scala 96:25:@31762.4 package.scala 96:25:@31763.4]
  assign _T_289 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@31770.4 package.scala 96:25:@31771.4]
  assign _T_292 = ~ _T_289; // @[SpatialBlocks.scala 138:93:@31773.4]
  assign io_in_x348_TREADY = x607_kernelx607_concrete1_io_in_x348_TREADY; // @[sm_x607.scala 63:23:@31880.4]
  assign io_in_x529_valid = x607_kernelx607_concrete1_io_in_x529_valid; // @[sm_x607.scala 64:23:@31884.4]
  assign io_in_x529_bits_addr = x607_kernelx607_concrete1_io_in_x529_bits_addr; // @[sm_x607.scala 64:23:@31883.4]
  assign io_in_x529_bits_size = x607_kernelx607_concrete1_io_in_x529_bits_size; // @[sm_x607.scala 64:23:@31882.4]
  assign io_in_x349_TVALID = x607_kernelx607_concrete1_io_in_x349_TVALID; // @[sm_x607.scala 65:23:@31894.4]
  assign io_in_x349_TDATA = x607_kernelx607_concrete1_io_in_x349_TDATA; // @[sm_x607.scala 65:23:@31892.4]
  assign io_in_x530_valid = x607_kernelx607_concrete1_io_in_x530_valid; // @[sm_x607.scala 66:23:@31897.4]
  assign io_in_x530_bits_wdata_0 = x607_kernelx607_concrete1_io_in_x530_bits_wdata_0; // @[sm_x607.scala 66:23:@31896.4]
  assign io_in_x530_bits_wstrb = x607_kernelx607_concrete1_io_in_x530_bits_wstrb; // @[sm_x607.scala 66:23:@31895.4]
  assign io_in_x531_ready = x607_kernelx607_concrete1_io_in_x531_ready; // @[sm_x607.scala 68:23:@31906.4]
  assign io_sigsOut_smDoneIn_0 = x607_sm_io_done; // @[SpatialBlocks.scala 156:53:@31780.4]
  assign x350_outbuf_0_clock = clock; // @[:@31633.4]
  assign x350_outbuf_0_reset = reset; // @[:@31634.4]
  assign x350_outbuf_0_io_rPort_0_ofs_0 = x607_kernelx607_concrete1_io_in_x350_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@31902.4]
  assign x350_outbuf_0_io_rPort_0_en_0 = x607_kernelx607_concrete1_io_in_x350_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@31901.4]
  assign x350_outbuf_0_io_rPort_0_backpressure = x607_kernelx607_concrete1_io_in_x350_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@31900.4]
  assign x607_sm_clock = clock; // @[:@31691.4]
  assign x607_sm_reset = reset; // @[:@31692.4]
  assign x607_sm_io_enable = _T_283 & _T_292; // @[SpatialBlocks.scala 140:18:@31777.4]
  assign x607_sm_io_ctrDone = x607_sm_io_ctrInc & _T_269; // @[sm_RootController.scala 82:26:@31727.4]
  assign x607_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@31779.4]
  assign x607_sm_io_doneIn_0 = x607_kernelx607_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@31747.4]
  assign x607_sm_io_doneIn_1 = x607_kernelx607_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@31748.4]
  assign RetimeWrapper_clock = clock; // @[:@31758.4]
  assign RetimeWrapper_reset = reset; // @[:@31759.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@31761.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@31760.4]
  assign RetimeWrapper_1_clock = clock; // @[:@31766.4]
  assign RetimeWrapper_1_reset = reset; // @[:@31767.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@31769.4]
  assign RetimeWrapper_1_io_in = x607_sm_io_done; // @[package.scala 94:16:@31768.4]
  assign x607_kernelx607_concrete1_clock = clock; // @[:@31795.4]
  assign x607_kernelx607_concrete1_reset = reset; // @[:@31796.4]
  assign x607_kernelx607_concrete1_io_in_x348_TVALID = io_in_x348_TVALID; // @[sm_x607.scala 63:23:@31881.4]
  assign x607_kernelx607_concrete1_io_in_x348_TDATA = io_in_x348_TDATA; // @[sm_x607.scala 63:23:@31879.4]
  assign x607_kernelx607_concrete1_io_in_x348_TID = io_in_x348_TID; // @[sm_x607.scala 63:23:@31875.4]
  assign x607_kernelx607_concrete1_io_in_x348_TDEST = io_in_x348_TDEST; // @[sm_x607.scala 63:23:@31874.4]
  assign x607_kernelx607_concrete1_io_in_x529_ready = io_in_x529_ready; // @[sm_x607.scala 64:23:@31885.4]
  assign x607_kernelx607_concrete1_io_in_x349_TREADY = io_in_x349_TREADY; // @[sm_x607.scala 65:23:@31893.4]
  assign x607_kernelx607_concrete1_io_in_x530_ready = io_in_x530_ready; // @[sm_x607.scala 66:23:@31898.4]
  assign x607_kernelx607_concrete1_io_in_x350_outbuf_0_rPort_0_output_0 = x350_outbuf_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@31899.4]
  assign x607_kernelx607_concrete1_io_in_x531_valid = io_in_x531_valid; // @[sm_x607.scala 68:23:@31905.4]
  assign x607_kernelx607_concrete1_io_in_x346_outdram_number = io_in_x346_outdram_number; // @[sm_x607.scala 69:31:@31907.4]
  assign x607_kernelx607_concrete1_io_sigsIn_smEnableOuts_0 = x607_sm_io_enableOut_0; // @[sm_x607.scala 107:22:@31918.4]
  assign x607_kernelx607_concrete1_io_sigsIn_smEnableOuts_1 = x607_sm_io_enableOut_1; // @[sm_x607.scala 107:22:@31919.4]
  assign x607_kernelx607_concrete1_io_sigsIn_smChildAcks_0 = x607_sm_io_childAck_0; // @[sm_x607.scala 107:22:@31914.4]
  assign x607_kernelx607_concrete1_io_sigsIn_smChildAcks_1 = x607_sm_io_childAck_1; // @[sm_x607.scala 107:22:@31915.4]
  assign x607_kernelx607_concrete1_io_rr = io_rr; // @[sm_x607.scala 106:18:@31908.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_269 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_269 <= 1'h0;
    end else begin
      _T_269 <= _T_266;
    end
  end
endmodule
module AccelUnit( // @[:@31941.2]
  input          clock, // @[:@31942.4]
  input          reset, // @[:@31943.4]
  input          io_enable, // @[:@31944.4]
  output         io_done, // @[:@31944.4]
  input          io_reset, // @[:@31944.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@31944.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@31944.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@31944.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@31944.4]
  output         io_memStreams_loads_0_data_ready, // @[:@31944.4]
  input          io_memStreams_loads_0_data_valid, // @[:@31944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@31944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@31944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@31944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@31944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@31944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@31944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@31944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@31944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@31944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@31944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@31944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@31944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@31944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@31944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@31944.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@31944.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@31944.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@31944.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@31944.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@31944.4]
  input          io_memStreams_stores_0_data_ready, // @[:@31944.4]
  output         io_memStreams_stores_0_data_valid, // @[:@31944.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_0, // @[:@31944.4]
  output         io_memStreams_stores_0_data_bits_wstrb, // @[:@31944.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@31944.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@31944.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@31944.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@31944.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@31944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@31944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@31944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@31944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@31944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@31944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@31944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@31944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@31944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@31944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@31944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@31944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@31944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@31944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@31944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@31944.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@31944.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@31944.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@31944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@31944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@31944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@31944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@31944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@31944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@31944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@31944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@31944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@31944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@31944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@31944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@31944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@31944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@31944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@31944.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@31944.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@31944.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@31944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@31944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@31944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@31944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@31944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@31944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@31944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@31944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@31944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@31944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@31944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@31944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@31944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@31944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@31944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@31944.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@31944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@31944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@31944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@31944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@31944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@31944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@31944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@31944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@31944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@31944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@31944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@31944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@31944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@31944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@31944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@31944.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@31944.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@31944.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@31944.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@31944.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@31944.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@31944.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@31944.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@31944.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@31944.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@31944.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@31944.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@31944.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@31944.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@31944.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@31944.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@31944.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@31944.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@31944.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@31944.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@31944.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@31944.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@31944.4]
  output         io_heap_0_req_valid, // @[:@31944.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@31944.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@31944.4]
  input          io_heap_0_resp_valid, // @[:@31944.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@31944.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@31944.4]
  input  [63:0]  io_argIns_0, // @[:@31944.4]
  input  [63:0]  io_argIns_1, // @[:@31944.4]
  input          io_argOuts_0_port_ready, // @[:@31944.4]
  output         io_argOuts_0_port_valid, // @[:@31944.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@31944.4]
  input  [63:0]  io_argOuts_0_echo // @[:@31944.4]
);
  wire  SingleCounter_clock; // @[Main.scala 40:32:@32092.4]
  wire  SingleCounter_reset; // @[Main.scala 40:32:@32092.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 40:32:@32092.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 40:32:@32092.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@32110.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@32110.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@32110.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@32110.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@32110.4]
  wire  SRFF_clock; // @[Main.scala 44:28:@32119.4]
  wire  SRFF_reset; // @[Main.scala 44:28:@32119.4]
  wire  SRFF_io_input_set; // @[Main.scala 44:28:@32119.4]
  wire  SRFF_io_input_reset; // @[Main.scala 44:28:@32119.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 44:28:@32119.4]
  wire  SRFF_io_output; // @[Main.scala 44:28:@32119.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 36:18:@32158.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 36:18:@32158.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 36:18:@32158.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 36:18:@32158.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 36:18:@32158.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 36:18:@32158.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 36:18:@32158.4]
  wire  RootController_sm_io_parentAck; // @[sm_RootController.scala 36:18:@32158.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 36:18:@32158.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 36:18:@32158.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 36:18:@32158.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32190.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32190.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32190.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@32190.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@32190.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 91:24:@32252.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 91:24:@32252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x348_TVALID; // @[sm_RootController.scala 91:24:@32252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x348_TREADY; // @[sm_RootController.scala 91:24:@32252.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x348_TDATA; // @[sm_RootController.scala 91:24:@32252.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x348_TID; // @[sm_RootController.scala 91:24:@32252.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x348_TDEST; // @[sm_RootController.scala 91:24:@32252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x529_ready; // @[sm_RootController.scala 91:24:@32252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x529_valid; // @[sm_RootController.scala 91:24:@32252.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x529_bits_addr; // @[sm_RootController.scala 91:24:@32252.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x529_bits_size; // @[sm_RootController.scala 91:24:@32252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x349_TVALID; // @[sm_RootController.scala 91:24:@32252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x349_TREADY; // @[sm_RootController.scala 91:24:@32252.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x349_TDATA; // @[sm_RootController.scala 91:24:@32252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x530_ready; // @[sm_RootController.scala 91:24:@32252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x530_valid; // @[sm_RootController.scala 91:24:@32252.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x530_bits_wdata_0; // @[sm_RootController.scala 91:24:@32252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x530_bits_wstrb; // @[sm_RootController.scala 91:24:@32252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x531_ready; // @[sm_RootController.scala 91:24:@32252.4]
  wire  RootController_kernelRootController_concrete1_io_in_x531_valid; // @[sm_RootController.scala 91:24:@32252.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x346_outdram_number; // @[sm_RootController.scala 91:24:@32252.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 91:24:@32252.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 91:24:@32252.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 91:24:@32252.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 91:24:@32252.4]
  wire  _T_599; // @[package.scala 96:25:@32115.4 package.scala 96:25:@32116.4]
  wire  _T_664; // @[Main.scala 46:50:@32186.4]
  wire  _T_665; // @[Main.scala 46:59:@32187.4]
  wire  _T_677; // @[package.scala 100:49:@32207.4]
  reg  _T_680; // @[package.scala 48:56:@32208.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 40:32:@32092.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@32110.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 44:28:@32119.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 36:18:@32158.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_parentAck(RootController_sm_io_parentAck),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@32190.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 91:24:@32252.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x348_TVALID(RootController_kernelRootController_concrete1_io_in_x348_TVALID),
    .io_in_x348_TREADY(RootController_kernelRootController_concrete1_io_in_x348_TREADY),
    .io_in_x348_TDATA(RootController_kernelRootController_concrete1_io_in_x348_TDATA),
    .io_in_x348_TID(RootController_kernelRootController_concrete1_io_in_x348_TID),
    .io_in_x348_TDEST(RootController_kernelRootController_concrete1_io_in_x348_TDEST),
    .io_in_x529_ready(RootController_kernelRootController_concrete1_io_in_x529_ready),
    .io_in_x529_valid(RootController_kernelRootController_concrete1_io_in_x529_valid),
    .io_in_x529_bits_addr(RootController_kernelRootController_concrete1_io_in_x529_bits_addr),
    .io_in_x529_bits_size(RootController_kernelRootController_concrete1_io_in_x529_bits_size),
    .io_in_x349_TVALID(RootController_kernelRootController_concrete1_io_in_x349_TVALID),
    .io_in_x349_TREADY(RootController_kernelRootController_concrete1_io_in_x349_TREADY),
    .io_in_x349_TDATA(RootController_kernelRootController_concrete1_io_in_x349_TDATA),
    .io_in_x530_ready(RootController_kernelRootController_concrete1_io_in_x530_ready),
    .io_in_x530_valid(RootController_kernelRootController_concrete1_io_in_x530_valid),
    .io_in_x530_bits_wdata_0(RootController_kernelRootController_concrete1_io_in_x530_bits_wdata_0),
    .io_in_x530_bits_wstrb(RootController_kernelRootController_concrete1_io_in_x530_bits_wstrb),
    .io_in_x531_ready(RootController_kernelRootController_concrete1_io_in_x531_ready),
    .io_in_x531_valid(RootController_kernelRootController_concrete1_io_in_x531_valid),
    .io_in_x346_outdram_number(RootController_kernelRootController_concrete1_io_in_x346_outdram_number),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@32115.4 package.scala 96:25:@32116.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 46:50:@32186.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 46:59:@32187.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@32207.4]
  assign io_done = SRFF_io_output; // @[Main.scala 53:23:@32206.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x529_valid; // @[sm_RootController.scala 61:23:@32324.4]
  assign io_memStreams_stores_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x529_bits_addr; // @[sm_RootController.scala 61:23:@32323.4]
  assign io_memStreams_stores_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x529_bits_size; // @[sm_RootController.scala 61:23:@32322.4]
  assign io_memStreams_stores_0_data_valid = RootController_kernelRootController_concrete1_io_in_x530_valid; // @[sm_RootController.scala 63:23:@32337.4]
  assign io_memStreams_stores_0_data_bits_wdata_0 = RootController_kernelRootController_concrete1_io_in_x530_bits_wdata_0; // @[sm_RootController.scala 63:23:@32336.4]
  assign io_memStreams_stores_0_data_bits_wstrb = RootController_kernelRootController_concrete1_io_in_x530_bits_wstrb; // @[sm_RootController.scala 63:23:@32335.4]
  assign io_memStreams_stores_0_wresp_ready = RootController_kernelRootController_concrete1_io_in_x531_ready; // @[sm_RootController.scala 64:23:@32341.4]
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x348_TREADY; // @[sm_RootController.scala 60:23:@32320.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x349_TVALID; // @[sm_RootController.scala 62:23:@32334.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x349_TDATA; // @[sm_RootController.scala 62:23:@32332.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 62:23:@32331.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 62:23:@32330.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 62:23:@32329.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 62:23:@32328.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 62:23:@32327.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 62:23:@32326.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@32093.4]
  assign SingleCounter_reset = reset; // @[:@32094.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 41:79:@32108.4]
  assign RetimeWrapper_clock = clock; // @[:@32111.4]
  assign RetimeWrapper_reset = reset; // @[:@32112.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@32114.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@32113.4]
  assign SRFF_clock = clock; // @[:@32120.4]
  assign SRFF_reset = reset; // @[:@32121.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 62:29:@32370.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 51:31:@32204.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 52:36:@32205.4]
  assign RootController_sm_clock = clock; // @[:@32159.4]
  assign RootController_sm_reset = reset; // @[:@32160.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 50:33:@32203.4 SpatialBlocks.scala 140:18:@32237.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@32231.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 54:34:@32211.4]
  assign RootController_sm_io_parentAck = 1'h0; // @[Main.scala 49:36:@32199.4 SpatialBlocks.scala 142:21:@32239.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@32228.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32191.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32192.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@32194.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@32193.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@32253.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@32254.4]
  assign RootController_kernelRootController_concrete1_io_in_x348_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 60:23:@32321.4]
  assign RootController_kernelRootController_concrete1_io_in_x348_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 60:23:@32319.4]
  assign RootController_kernelRootController_concrete1_io_in_x348_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 60:23:@32315.4]
  assign RootController_kernelRootController_concrete1_io_in_x348_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 60:23:@32314.4]
  assign RootController_kernelRootController_concrete1_io_in_x529_ready = io_memStreams_stores_0_cmd_ready; // @[sm_RootController.scala 61:23:@32325.4]
  assign RootController_kernelRootController_concrete1_io_in_x349_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 62:23:@32333.4]
  assign RootController_kernelRootController_concrete1_io_in_x530_ready = io_memStreams_stores_0_data_ready; // @[sm_RootController.scala 63:23:@32338.4]
  assign RootController_kernelRootController_concrete1_io_in_x531_valid = io_memStreams_stores_0_wresp_valid; // @[sm_RootController.scala 64:23:@32340.4]
  assign RootController_kernelRootController_concrete1_io_in_x346_outdram_number = io_argIns_1; // @[sm_RootController.scala 65:31:@32342.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 96:22:@32351.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 96:22:@32349.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 95:18:@32343.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module SpatialIP( // @[:@32372.2]
  input         clock, // @[:@32373.4]
  input         reset, // @[:@32374.4]
  input  [31:0] io_raddr, // @[:@32375.4]
  input         io_wen, // @[:@32375.4]
  input  [31:0] io_waddr, // @[:@32375.4]
  input  [63:0] io_wdata, // @[:@32375.4]
  output [63:0] io_rdata // @[:@32375.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@32377.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@32377.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@32377.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@32377.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@32377.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@32377.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@32377.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@32377.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@32377.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@32377.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@32377.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@32377.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  assign io_rdata = 64'h0;
  assign accel_clock = clock; // @[:@32378.4]
  assign accel_reset = reset; // @[:@32379.4]
  assign accel_io_enable = 1'h0;
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_loads_0_data_valid = 1'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0;
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_stores_0_data_ready = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0;
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0;
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0;
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0;
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = 1'h0;
  assign accel_io_heap_0_resp_bits_allocDealloc = 1'h0;
  assign accel_io_heap_0_resp_bits_sizeAddr = 64'h0;
  assign accel_io_argIns_0 = 64'h0;
  assign accel_io_argIns_1 = 64'h0;
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0;
endmodule
