// Latency = 4
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [31:0] I_0,
  output [31:0] O_0
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(clock), // @[:@1296.4]
    .reset(reset), // @[:@1297.4]
    .io_in_x184_TREADY(dontcare), // @[:@1298.4]
    .io_in_x184_TDATA(I_0), // @[:@1298.4]
    .io_in_x184_TID(8'h0),
    .io_in_x184_TDEST(8'h0),
    .io_in_x185_TVALID(valid_down), // @[:@1298.4]
    .io_in_x185_TDATA(O_0), // @[:@1298.4]
    .io_in_x185_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x192_ctrchain cchain ( // @[:@2879.2]
    .clock(clock), // @[:@2880.4]
    .reset(reset), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule


module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule


// End boilerplate
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 321:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 325:12:@24.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : io_wPort_0_data_0; // @[MemPrimitives.scala 325:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        ff <= io_wPort_0_data_0;
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh42); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh42); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_parentAck, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  _T_81; // @[Controllers.scala 86:43:@328.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_93; // @[Controllers.scala 92:52:@342.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_134; // @[Controllers.scala 129:57:@382.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  wire  _T_167; // @[package.scala 100:41:@414.4]
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign _T_81 = io_rst | done_0_io_output; // @[Controllers.scala 86:43:@328.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_93 = synchronize | io_rst; // @[Controllers.scala 92:52:@342.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_134 = _T_133 | io_parentAck; // @[Controllers.scala 129:57:@382.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign _T_167 = done_0_io_output & _T_166; // @[package.scala 100:41:@414.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_134 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = _T_81 | io_parentAck; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = _T_93 | io_parentAck; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = _T_167 | io_parentAck; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module SRAM( // @[:@507.2]
  input         clock, // @[:@508.4]
  input  [20:0] io_raddr, // @[:@510.4]
  output [31:0] io_rdata, // @[:@510.4]
  input         io_backpressure // @[:@510.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@512.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@512.4]
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(2073600), .AWIDTH(21)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@512.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign io_rdata = SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@539.4]
  assign SRAMVerilogAWS_wdata = 32'h0; // @[SRAM.scala 175:20:@526.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@527.4]
  assign SRAMVerilogAWS_wen = 1'h0; // @[SRAM.scala 173:18:@524.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@529.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@528.4]
  assign SRAMVerilogAWS_waddr = 21'h0; // @[SRAM.scala 174:20:@525.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@523.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@522.4]
endmodule
module RetimeWrapper_5( // @[:@553.2]
  input         clock, // @[:@554.4]
  input         reset, // @[:@555.4]
  input         io_flow, // @[:@556.4]
  input  [20:0] io_in, // @[:@556.4]
  output [20:0] io_out // @[:@556.4]
);
  wire [20:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@558.4]
  RetimeShiftRegister #(.WIDTH(21), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@558.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@571.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@570.4]
  assign sr_init = 21'h0; // @[RetimeShiftRegister.scala 19:16:@569.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@568.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@567.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@565.4]
endmodule
module Mem1D( // @[:@573.2]
  input         clock, // @[:@574.4]
  input         reset, // @[:@575.4]
  input  [20:0] io_r_ofs_0, // @[:@576.4]
  input         io_r_backpressure, // @[:@576.4]
  output [31:0] io_output // @[:@576.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@580.4]
  wire [20:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@580.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@580.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@580.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_in; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_out; // @[package.scala 93:22:@583.4]
  SRAM SRAM ( // @[MemPrimitives.scala 715:21:@580.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@583.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@596.4]
  assign SRAM_clock = clock; // @[:@581.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@590.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@595.4]
  assign RetimeWrapper_clock = clock; // @[:@584.4]
  assign RetimeWrapper_reset = reset; // @[:@585.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@587.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@586.4]
endmodule
module StickySelects( // @[:@598.2]
  input   io_ins_0, // @[:@601.4]
  output  io_outs_0 // @[:@601.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 34:26:@603.4]
endmodule
module RetimeWrapper_6( // @[:@617.2]
  input   clock, // @[:@618.4]
  input   reset, // @[:@619.4]
  input   io_flow, // @[:@620.4]
  input   io_in, // @[:@620.4]
  output  io_out // @[:@620.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@622.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@622.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@635.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@634.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@633.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@632.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@631.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@629.4]
endmodule
module x186_outbuf_0( // @[:@637.2]
  input         clock, // @[:@638.4]
  input         reset, // @[:@639.4]
  input  [20:0] io_rPort_0_ofs_0, // @[:@640.4]
  input         io_rPort_0_en_0, // @[:@640.4]
  input         io_rPort_0_backpressure, // @[:@640.4]
  output [31:0] io_rPort_0_output_0 // @[:@640.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@655.4]
  wire [20:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@655.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@655.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@695.4]
  wire  _T_76; // @[MemPrimitives.scala 126:35:@685.4]
  wire [22:0] _T_78; // @[Cat.scala 30:58:@687.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@655.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@681.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@695.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@685.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@687.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@702.4]
  assign Mem1D_clock = clock; // @[:@656.4]
  assign Mem1D_reset = reset; // @[:@657.4]
  assign Mem1D_io_r_ofs_0 = _T_78[20:0]; // @[MemPrimitives.scala 131:28:@691.4]
  assign Mem1D_io_r_backpressure = _T_78[21]; // @[MemPrimitives.scala 132:32:@692.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@684.4]
  assign RetimeWrapper_clock = clock; // @[:@696.4]
  assign RetimeWrapper_reset = reset; // @[:@697.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@699.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@698.4]
endmodule
module x455_sm( // @[:@846.2]
  input   clock, // @[:@847.4]
  input   reset, // @[:@848.4]
  input   io_enable, // @[:@849.4]
  output  io_done, // @[:@849.4]
  input   io_ctrDone, // @[:@849.4]
  output  io_ctrInc, // @[:@849.4]
  input   io_parentAck, // @[:@849.4]
  input   io_doneIn_0, // @[:@849.4]
  input   io_doneIn_1, // @[:@849.4]
  output  io_enableOut_0, // @[:@849.4]
  output  io_enableOut_1, // @[:@849.4]
  output  io_childAck_0, // @[:@849.4]
  output  io_childAck_1 // @[:@849.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@852.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@855.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@858.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@861.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@893.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1011.4]
  wire  allDone; // @[Controllers.scala 80:47:@864.4]
  wire  synchronize; // @[Controllers.scala 146:56:@918.4]
  wire  _T_127; // @[Controllers.scala 150:35:@920.4]
  wire  _T_129; // @[Controllers.scala 150:60:@921.4]
  wire  _T_130; // @[Controllers.scala 150:58:@922.4]
  wire  _T_132; // @[Controllers.scala 150:76:@923.4]
  wire  _T_133; // @[Controllers.scala 150:74:@924.4]
  wire  _T_135; // @[Controllers.scala 150:97:@925.4]
  wire  _T_136; // @[Controllers.scala 150:95:@926.4]
  wire  _T_152; // @[Controllers.scala 150:35:@944.4]
  wire  _T_154; // @[Controllers.scala 150:60:@945.4]
  wire  _T_155; // @[Controllers.scala 150:58:@946.4]
  wire  _T_157; // @[Controllers.scala 150:76:@947.4]
  wire  _T_158; // @[Controllers.scala 150:74:@948.4]
  wire  _T_161; // @[Controllers.scala 150:95:@950.4]
  wire  _T_179; // @[Controllers.scala 213:68:@972.4]
  wire  _T_181; // @[Controllers.scala 213:90:@974.4]
  wire  _T_183; // @[Controllers.scala 213:132:@976.4]
  wire  _T_184; // @[Controllers.scala 213:130:@977.4]
  wire  _T_185; // @[Controllers.scala 213:156:@978.4]
  wire  _T_187; // @[Controllers.scala 213:68:@981.4]
  wire  _T_189; // @[Controllers.scala 213:90:@983.4]
  wire  _T_196; // @[package.scala 100:49:@989.4]
  reg  _T_199; // @[package.scala 48:56:@990.4]
  reg [31:0] _RAND_0;
  wire  _T_200; // @[package.scala 100:41:@992.4]
  reg  _T_213; // @[package.scala 48:56:@1008.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@852.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@855.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@858.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@861.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@890.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@893.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@994.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1011.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@864.4]
  assign synchronize = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 146:56:@918.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 150:35:@920.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 150:60:@921.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 150:58:@922.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 150:76:@923.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 150:74:@924.4]
  assign _T_135 = io_ctrDone == 1'h0; // @[Controllers.scala 150:97:@925.4]
  assign _T_136 = _T_133 & _T_135; // @[Controllers.scala 150:95:@926.4]
  assign _T_152 = ~ iterDone_1_io_output; // @[Controllers.scala 150:35:@944.4]
  assign _T_154 = io_doneIn_1 == 1'h0; // @[Controllers.scala 150:60:@945.4]
  assign _T_155 = _T_152 & _T_154; // @[Controllers.scala 150:58:@946.4]
  assign _T_157 = done_1_io_output == 1'h0; // @[Controllers.scala 150:76:@947.4]
  assign _T_158 = _T_155 & _T_157; // @[Controllers.scala 150:74:@948.4]
  assign _T_161 = _T_158 & _T_135; // @[Controllers.scala 150:95:@950.4]
  assign _T_179 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@972.4]
  assign _T_181 = _T_179 & _T_127; // @[Controllers.scala 213:90:@974.4]
  assign _T_183 = ~ allDone; // @[Controllers.scala 213:132:@976.4]
  assign _T_184 = _T_181 & _T_183; // @[Controllers.scala 213:130:@977.4]
  assign _T_185 = ~ io_ctrDone; // @[Controllers.scala 213:156:@978.4]
  assign _T_187 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@981.4]
  assign _T_189 = _T_187 & _T_152; // @[Controllers.scala 213:90:@983.4]
  assign _T_196 = allDone == 1'h0; // @[package.scala 100:49:@989.4]
  assign _T_200 = allDone & _T_199; // @[package.scala 100:41:@992.4]
  assign io_done = RetimeWrapper_1_io_out; // @[Controllers.scala 245:13:@1018.4]
  assign io_ctrInc = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 143:17:@917.4]
  assign io_enableOut_0 = _T_184 & _T_185; // @[Controllers.scala 213:55:@980.4]
  assign io_enableOut_1 = _T_189 & _T_183; // @[Controllers.scala 213:55:@988.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@969.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@971.4]
  assign active_0_clock = clock; // @[:@853.4]
  assign active_0_reset = reset; // @[:@854.4]
  assign active_0_io_input_set = _T_136 & io_enable; // @[Controllers.scala 150:32:@929.4]
  assign active_0_io_input_reset = io_doneIn_0 | io_parentAck; // @[Controllers.scala 151:34:@933.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@867.4]
  assign active_1_clock = clock; // @[:@856.4]
  assign active_1_reset = reset; // @[:@857.4]
  assign active_1_io_input_set = _T_161 & io_enable; // @[Controllers.scala 150:32:@953.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_parentAck; // @[Controllers.scala 151:34:@957.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@868.4]
  assign done_0_clock = clock; // @[:@859.4]
  assign done_0_reset = reset; // @[:@860.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@943.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@879.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@869.4]
  assign done_1_clock = clock; // @[:@862.4]
  assign done_1_reset = reset; // @[:@863.4]
  assign done_1_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@967.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@888.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@870.4]
  assign iterDone_0_clock = clock; // @[:@891.4]
  assign iterDone_0_reset = reset; // @[:@892.4]
  assign iterDone_0_io_input_set = io_doneIn_0; // @[Controllers.scala 152:34:@939.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@906.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@896.4]
  assign iterDone_1_clock = clock; // @[:@894.4]
  assign iterDone_1_reset = reset; // @[:@895.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 152:34:@963.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@915.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@897.4]
  assign RetimeWrapper_clock = clock; // @[:@995.4]
  assign RetimeWrapper_reset = reset; // @[:@996.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@998.4]
  assign RetimeWrapper_io_in = _T_200 | io_parentAck; // @[package.scala 94:16:@997.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1012.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1013.4]
  assign RetimeWrapper_1_io_flow = io_enable; // @[package.scala 95:18:@1015.4]
  assign RetimeWrapper_1_io_in = allDone & _T_213; // @[package.scala 94:16:@1014.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_199 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_213 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_199 <= 1'h0;
    end else begin
      _T_199 <= _T_196;
    end
    if (reset) begin
      _T_213 <= 1'h0;
    end else begin
      _T_213 <= _T_196;
    end
  end
endmodule
module x321_outr_UnitPipe_sm( // @[:@1435.2]
  input   clock, // @[:@1436.4]
  input   reset, // @[:@1437.4]
  input   io_enable, // @[:@1438.4]
  output  io_done, // @[:@1438.4]
  input   io_parentAck, // @[:@1438.4]
  input   io_doneIn_0, // @[:@1438.4]
  input   io_doneIn_1, // @[:@1438.4]
  output  io_enableOut_0, // @[:@1438.4]
  output  io_enableOut_1, // @[:@1438.4]
  output  io_childAck_0, // @[:@1438.4]
  output  io_childAck_1, // @[:@1438.4]
  input   io_ctrCopyDone_0, // @[:@1438.4]
  input   io_ctrCopyDone_1 // @[:@1438.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@1441.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@1444.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@1447.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1450.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1482.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1688.4]
  wire  allDone; // @[Controllers.scala 80:47:@1453.4]
  wire  _T_127; // @[Controllers.scala 165:35:@1507.4]
  wire  _T_129; // @[Controllers.scala 165:60:@1508.4]
  wire  _T_130; // @[Controllers.scala 165:58:@1509.4]
  wire  _T_132; // @[Controllers.scala 165:76:@1510.4]
  wire  _T_133; // @[Controllers.scala 165:74:@1511.4]
  wire  _T_137; // @[Controllers.scala 165:109:@1514.4]
  wire  _T_140; // @[Controllers.scala 165:141:@1516.4]
  wire  _T_148; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  wire  _T_152; // @[Controllers.scala 167:54:@1531.4]
  wire  _T_153; // @[Controllers.scala 167:52:@1532.4]
  wire  _T_160; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  wire  _T_178; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  wire  _T_182; // @[Controllers.scala 169:67:@1563.4]
  wire  _T_183; // @[Controllers.scala 169:86:@1564.4]
  wire  _T_195; // @[Controllers.scala 165:35:@1576.4]
  wire  _T_197; // @[Controllers.scala 165:60:@1577.4]
  wire  _T_198; // @[Controllers.scala 165:58:@1578.4]
  wire  _T_200; // @[Controllers.scala 165:76:@1579.4]
  wire  _T_201; // @[Controllers.scala 165:74:@1580.4]
  wire  _T_205; // @[Controllers.scala 165:109:@1583.4]
  wire  _T_208; // @[Controllers.scala 165:141:@1585.4]
  wire  _T_216; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  wire  _T_220; // @[Controllers.scala 167:54:@1600.4]
  wire  _T_221; // @[Controllers.scala 167:52:@1601.4]
  wire  _T_228; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  wire  _T_246; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  wire  _T_250; // @[Controllers.scala 169:67:@1632.4]
  wire  _T_251; // @[Controllers.scala 169:86:@1633.4]
  wire  _T_265; // @[Controllers.scala 213:68:@1649.4]
  wire  _T_267; // @[Controllers.scala 213:90:@1651.4]
  wire  _T_269; // @[Controllers.scala 213:132:@1653.4]
  wire  _T_273; // @[Controllers.scala 213:68:@1658.4]
  wire  _T_275; // @[Controllers.scala 213:90:@1660.4]
  wire  _T_282; // @[package.scala 100:49:@1666.4]
  reg  _T_285; // @[package.scala 48:56:@1667.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@1669.4]
  reg  _T_299; // @[package.scala 48:56:@1685.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@1441.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@1444.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@1447.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1450.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1479.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1482.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1523.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1537.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1555.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1592.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1606.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1624.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1671.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1688.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1453.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1507.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1508.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@1509.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1510.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@1511.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@1514.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1516.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@1531.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@1532.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@1563.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@1564.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1576.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1577.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@1578.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1579.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@1580.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@1583.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1585.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@1600.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@1601.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@1632.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@1633.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1649.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@1651.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@1653.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1658.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@1660.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@1666.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@1669.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@1695.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@1657.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@1665.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1646.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1648.4]
  assign active_0_clock = clock; // @[:@1442.4]
  assign active_0_reset = reset; // @[:@1443.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@1518.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1522.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1456.4]
  assign active_1_clock = clock; // @[:@1445.4]
  assign active_1_reset = reset; // @[:@1446.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@1587.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1591.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1457.4]
  assign done_0_clock = clock; // @[:@1448.4]
  assign done_0_reset = reset; // @[:@1449.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@1568.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1468.4 Controllers.scala 170:32:@1575.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1458.4]
  assign done_1_clock = clock; // @[:@1451.4]
  assign done_1_reset = reset; // @[:@1452.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@1637.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1477.4 Controllers.scala 170:32:@1644.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1459.4]
  assign iterDone_0_clock = clock; // @[:@1480.4]
  assign iterDone_0_reset = reset; // @[:@1481.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@1536.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@1495.4 Controllers.scala 168:36:@1552.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1485.4]
  assign iterDone_1_clock = clock; // @[:@1483.4]
  assign iterDone_1_reset = reset; // @[:@1484.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@1605.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@1504.4 Controllers.scala 168:36:@1621.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1486.4]
  assign RetimeWrapper_clock = clock; // @[:@1524.4]
  assign RetimeWrapper_reset = reset; // @[:@1525.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1527.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1526.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1538.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1539.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1541.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1540.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1556.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1557.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1559.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1558.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1593.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1594.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1596.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1595.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1607.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1608.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1610.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1609.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1625.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1626.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1628.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1627.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1672.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1673.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1675.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@1674.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1689.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1690.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@1692.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@1691.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module CompactingIncDincCtr( // @[:@1924.2]
  input   clock, // @[:@1925.4]
  input   reset, // @[:@1926.4]
  input   io_input_inc_en_0, // @[:@1927.4]
  input   io_input_dinc_en_0, // @[:@1927.4]
  output  io_output_full // @[:@1927.4]
);
  reg [31:0] cnt; // @[Counter.scala 170:20:@1929.4]
  reg [31:0] _RAND_0;
  wire [14:0] numPushed; // @[Counter.scala 172:47:@1930.4]
  wire [14:0] numPopped; // @[Counter.scala 173:48:@1931.4]
  wire [31:0] _GEN_0; // @[Counter.scala 174:14:@1932.4]
  wire [32:0] _T_37; // @[Counter.scala 174:14:@1932.4]
  wire [31:0] _T_38; // @[Counter.scala 174:14:@1933.4]
  wire [31:0] _T_39; // @[Counter.scala 174:14:@1934.4]
  wire [31:0] _GEN_1; // @[Counter.scala 174:26:@1935.4]
  wire [32:0] _T_40; // @[Counter.scala 174:26:@1935.4]
  wire [31:0] _T_41; // @[Counter.scala 174:26:@1936.4]
  wire [31:0] _T_42; // @[Counter.scala 174:26:@1937.4]
  assign numPushed = io_input_inc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 172:47:@1930.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 173:48:@1931.4]
  assign _GEN_0 = {{17{numPushed[14]}},numPushed}; // @[Counter.scala 174:14:@1932.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1932.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1933.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 174:14:@1934.4]
  assign _GEN_1 = {{17{numPopped[14]}},numPopped}; // @[Counter.scala 174:26:@1935.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1935.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1936.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 174:26:@1937.4]
  assign io_output_full = $signed(cnt) > $signed(32'sh1dff); // @[Counter.scala 180:18:@1951.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module x187_fifoinraw_0( // @[:@2074.2]
  input   clock, // @[:@2075.4]
  input   reset // @[:@2076.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2121.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2121.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign elements_clock = clock; // @[:@2122.4]
  assign elements_reset = reset; // @[:@2123.4]
  assign elements_io_input_inc_en_0 = 1'h0; // @[MemPrimitives.scala 394:79:@2133.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2134.4]
endmodule
module x188_fifoinpacked_0( // @[:@2497.2]
  input   clock, // @[:@2498.4]
  input   reset, // @[:@2499.4]
  input   io_wPort_0_en_0, // @[:@2500.4]
  output  io_full, // @[:@2500.4]
  input   io_active_0_in, // @[:@2500.4]
  output  io_active_0_out // @[:@2500.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2544.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2544.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 439:39:@2618.4]
  assign io_active_0_out = io_active_0_in; // @[MemPrimitives.scala 437:129:@2616.4]
  assign elements_clock = clock; // @[:@2545.4]
  assign elements_reset = reset; // @[:@2546.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 394:79:@2556.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2557.4]
endmodule
module FF_7( // @[:@3047.2]
  input         clock, // @[:@3048.4]
  input         reset, // @[:@3049.4]
  output [12:0] io_rPort_0_output_0, // @[:@3050.4]
  input  [12:0] io_wPort_0_data_0, // @[:@3050.4]
  input         io_wPort_0_reset, // @[:@3050.4]
  input         io_wPort_0_en_0 // @[:@3050.4]
);
  reg [12:0] ff; // @[MemPrimitives.scala 321:19:@3065.4]
  reg [31:0] _RAND_0;
  wire [12:0] _T_68; // @[MemPrimitives.scala 325:32:@3067.4]
  wire [12:0] _T_69; // @[MemPrimitives.scala 325:12:@3068.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@3067.4]
  assign _T_69 = io_wPort_0_reset ? 13'h0 : _T_68; // @[MemPrimitives.scala 325:12:@3068.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@3070.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 13'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 13'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_1( // @[:@3085.2]
  input         clock, // @[:@3086.4]
  input         reset, // @[:@3087.4]
  input         io_setup_saturate, // @[:@3088.4]
  input         io_input_reset, // @[:@3088.4]
  input         io_input_enable, // @[:@3088.4]
  output [12:0] io_output_count_0, // @[:@3088.4]
  output        io_output_oobs_0, // @[:@3088.4]
  output        io_output_done, // @[:@3088.4]
  output        io_output_saturated // @[:@3088.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3101.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3117.4]
  wire  _T_36; // @[Counter.scala 264:45:@3120.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3145.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3146.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3147.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3148.4]
  wire  _T_57; // @[Counter.scala 293:18:@3150.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3158.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3160.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3161.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3162.4]
  wire  _T_75; // @[Counter.scala 322:102:@3166.4]
  wire  _T_77; // @[Counter.scala 322:130:@3167.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3101.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3117.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3120.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3145.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3146.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3147.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3148.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh438); // @[Counter.scala 293:18:@3150.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3158.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3160.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3161.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3162.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3166.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh438); // @[Counter.scala 322:130:@3167.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3165.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3169.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3171.4]
  assign io_output_saturated = io_setup_saturate & _T_57; // @[Counter.scala 340:25:@3174.4]
  assign bases_0_clock = clock; // @[:@3102.4]
  assign bases_0_reset = reset; // @[:@3103.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3164.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3143.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3144.4]
  assign SRFF_clock = clock; // @[:@3118.4]
  assign SRFF_reset = reset; // @[:@3119.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3122.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3124.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3125.4]
endmodule
module SingleCounter_2( // @[:@3214.2]
  input         clock, // @[:@3215.4]
  input         reset, // @[:@3216.4]
  input         io_setup_saturate, // @[:@3217.4]
  input         io_input_reset, // @[:@3217.4]
  input         io_input_enable, // @[:@3217.4]
  output [12:0] io_output_count_0, // @[:@3217.4]
  output        io_output_oobs_0, // @[:@3217.4]
  output        io_output_done // @[:@3217.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3230.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3246.4]
  wire  _T_36; // @[Counter.scala 264:45:@3249.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3274.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3275.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3276.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3277.4]
  wire  _T_57; // @[Counter.scala 293:18:@3279.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3287.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3289.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3290.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3291.4]
  wire  _T_75; // @[Counter.scala 322:102:@3295.4]
  wire  _T_77; // @[Counter.scala 322:130:@3296.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3230.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3246.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3249.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3274.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3275.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3276.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3277.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh780); // @[Counter.scala 293:18:@3279.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3287.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3289.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3290.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3291.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3295.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh780); // @[Counter.scala 322:130:@3296.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3294.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3298.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3300.4]
  assign bases_0_clock = clock; // @[:@3231.4]
  assign bases_0_reset = reset; // @[:@3232.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3293.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3272.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3273.4]
  assign SRFF_clock = clock; // @[:@3247.4]
  assign SRFF_reset = reset; // @[:@3248.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3251.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3253.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3254.4]
endmodule
module x192_ctrchain( // @[:@3305.2]
  input         clock, // @[:@3306.4]
  input         reset, // @[:@3307.4]
  input         io_input_reset, // @[:@3308.4]
  input         io_input_enable, // @[:@3308.4]
  output [12:0] io_output_counts_1, // @[:@3308.4]
  output [12:0] io_output_counts_0, // @[:@3308.4]
  output        io_output_oobs_0, // @[:@3308.4]
  output        io_output_oobs_1, // @[:@3308.4]
  output        io_output_done // @[:@3308.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@3310.4]
  wire [12:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@3313.4]
  wire [12:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@3313.4]
  wire  isDone; // @[Counter.scala 541:51:@3330.4]
  reg  wasDone; // @[Counter.scala 542:24:@3331.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@3339.4]
  wire  _T_66; // @[Counter.scala 546:80:@3340.4]
  reg  doneLatch; // @[Counter.scala 550:26:@3345.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@3346.4]
  wire  _T_74; // @[Counter.scala 551:19:@3347.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@3310.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@3313.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@3330.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@3339.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@3340.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@3346.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@3347.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@3352.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@3349.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3351.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3354.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@3342.4]
  assign ctrs_0_clock = clock; // @[:@3311.4]
  assign ctrs_0_reset = reset; // @[:@3312.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 530:29:@3327.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3319.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@3326.4]
  assign ctrs_1_clock = clock; // @[:@3314.4]
  assign ctrs_1_reset = reset; // @[:@3315.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@3329.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3323.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@3324.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_21( // @[:@3394.2]
  input   clock, // @[:@3395.4]
  input   reset, // @[:@3396.4]
  input   io_flow, // @[:@3397.4]
  input   io_in, // @[:@3397.4]
  output  io_out // @[:@3397.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@3399.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3412.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3411.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3410.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3409.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3408.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3406.4]
endmodule
module RetimeWrapper_25( // @[:@3522.2]
  input   clock, // @[:@3523.4]
  input   reset, // @[:@3524.4]
  input   io_flow, // @[:@3525.4]
  input   io_in, // @[:@3525.4]
  output  io_out // @[:@3525.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@3527.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3540.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3539.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3538.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3537.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3536.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3534.4]
endmodule
module x206_inr_Foreach_sm( // @[:@3542.2]
  input   clock, // @[:@3543.4]
  input   reset, // @[:@3544.4]
  input   io_enable, // @[:@3545.4]
  output  io_done, // @[:@3545.4]
  output  io_doneLatch, // @[:@3545.4]
  input   io_ctrDone, // @[:@3545.4]
  output  io_datapathEn, // @[:@3545.4]
  output  io_ctrInc, // @[:@3545.4]
  output  io_ctrRst, // @[:@3545.4]
  input   io_parentAck, // @[:@3545.4]
  input   io_backpressure, // @[:@3545.4]
  input   io_break // @[:@3545.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3547.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3547.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3550.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3550.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3642.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3555.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3556.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3557.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3558.4]
  wire  _T_100; // @[package.scala 100:49:@3575.4]
  reg  _T_103; // @[package.scala 48:56:@3576.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  wire  _T_110; // @[package.scala 100:49:@3591.4]
  reg  _T_113; // @[package.scala 48:56:@3592.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3594.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3599.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3600.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3603.4]
  wire  _T_124; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  wire  _T_126; // @[package.scala 100:49:@3613.4]
  reg  _T_129; // @[package.scala 48:56:@3614.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3636.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3638.4]
  reg  _T_153; // @[package.scala 48:56:@3639.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3649.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3650.4]
  SRFF active ( // @[Controllers.scala 261:22:@3547.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3550.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@3584.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3606.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3618.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3626.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@3642.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3555.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3556.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3557.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3558.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3575.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3591.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3594.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3599.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3600.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3603.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3613.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3638.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3649.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3650.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3617.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3652.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3602.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3605.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3597.4]
  assign active_clock = clock; // @[:@3548.4]
  assign active_reset = reset; // @[:@3549.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3560.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3564.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3565.4]
  assign done_clock = clock; // @[:@3551.4]
  assign done_reset = reset; // @[:@3552.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3580.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3573.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3574.4]
  assign RetimeWrapper_clock = clock; // @[:@3585.4]
  assign RetimeWrapper_reset = reset; // @[:@3586.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3588.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3587.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3607.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3608.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3610.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3609.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3619.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3620.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3622.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3621.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3627.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3628.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3630.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3629.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3643.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3644.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3646.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3645.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module fix2fixBox( // @[:@3759.2]
  input  [31:0] io_a, // @[:@3762.4]
  output [31:0] io_b // @[:@3762.4]
);
  assign io_b = io_a; // @[Converter.scala 95:38:@3775.4]
endmodule
module _( // @[:@3777.2]
  input  [31:0] io_b, // @[:@3780.4]
  output [31:0] io_result // @[:@3780.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3785.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3785.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@3785.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3793.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3788.4]
endmodule
module fix2fixBox_2( // @[:@3831.2]
  input  [31:0] io_a, // @[:@3834.4]
  output [32:0] io_b // @[:@3834.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@3844.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@3844.4]
  assign io_b = {_T_20,io_a}; // @[Converter.scala 95:38:@3849.4]
endmodule
module __2( // @[:@3851.2]
  input  [31:0] io_b, // @[:@3854.4]
  output [32:0] io_result // @[:@3854.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3859.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3859.4]
  fix2fixBox_2 fix2fixBox ( // @[BigIPZynq.scala 219:30:@3859.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3867.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3862.4]
endmodule
module RetimeWrapper_29( // @[:@3919.2]
  input         clock, // @[:@3920.4]
  input         reset, // @[:@3921.4]
  input         io_flow, // @[:@3922.4]
  input  [31:0] io_in, // @[:@3922.4]
  output [31:0] io_out // @[:@3922.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3924.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3937.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3936.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3935.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3934.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3933.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3931.4]
endmodule
module fix2fixBox_4( // @[:@3939.2]
  input         clock, // @[:@3940.4]
  input         reset, // @[:@3941.4]
  input  [32:0] io_a, // @[:@3942.4]
  input         io_flow, // @[:@3942.4]
  output [31:0] io_b // @[:@3942.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3955.4]
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@3955.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@3962.4]
  assign RetimeWrapper_clock = clock; // @[:@3956.4]
  assign RetimeWrapper_reset = reset; // @[:@3957.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@3959.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@3958.4]
endmodule
module x370_sub( // @[:@3964.2]
  input         clock, // @[:@3965.4]
  input         reset, // @[:@3966.4]
  input  [31:0] io_a, // @[:@3967.4]
  input  [31:0] io_b, // @[:@3967.4]
  input         io_flow, // @[:@3967.4]
  output [31:0] io_result // @[:@3967.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@3975.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@3975.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@3982.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@3982.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@4001.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@4001.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@4001.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@3989.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@3990.4]
  __2 _ ( // @[Math.scala 720:24:@3975.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@3982.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 182:30:@4001.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@3989.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@3990.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@4009.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@3978.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@3985.4]
  assign fix2fixBox_clock = clock; // @[:@4002.4]
  assign fix2fixBox_reset = reset; // @[:@4003.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@4004.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@4007.4]
endmodule
module x198_sum( // @[:@4176.2]
  input         clock, // @[:@4177.4]
  input         reset, // @[:@4178.4]
  input  [31:0] io_a, // @[:@4179.4]
  input  [31:0] io_b, // @[:@4179.4]
  input         io_flow, // @[:@4179.4]
  output [31:0] io_result // @[:@4179.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4187.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@4187.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@4194.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@4194.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4212.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4212.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4212.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@4201.4]
  __2 _ ( // @[Math.scala 720:24:@4187.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@4194.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@4212.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4201.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4220.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@4190.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@4197.4]
  assign fix2fixBox_clock = clock; // @[:@4213.4]
  assign fix2fixBox_reset = reset; // @[:@4214.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4215.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4218.4]
endmodule
module x206_inr_Foreach_kernelx206_inr_Foreach_concrete1( // @[:@4712.2]
  input         clock, // @[:@4713.4]
  input         reset, // @[:@4714.4]
  output        io_in_x188_fifoinpacked_0_wPort_0_en_0, // @[:@4715.4]
  input         io_in_x188_fifoinpacked_0_full, // @[:@4715.4]
  output        io_in_x188_fifoinpacked_0_active_0_in, // @[:@4715.4]
  input         io_in_x188_fifoinpacked_0_active_0_out, // @[:@4715.4]
  input         io_sigsIn_backpressure, // @[:@4715.4]
  input         io_sigsIn_datapathEn, // @[:@4715.4]
  input         io_sigsIn_break, // @[:@4715.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_1, // @[:@4715.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@4715.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@4715.4]
  input         io_sigsIn_cchainOutputs_0_oobs_1, // @[:@4715.4]
  input         io_rr // @[:@4715.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4749.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@4749.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@4761.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@4761.4]
  wire  x370_sub_1_clock; // @[Math.scala 191:24:@4788.4]
  wire  x370_sub_1_reset; // @[Math.scala 191:24:@4788.4]
  wire [31:0] x370_sub_1_io_a; // @[Math.scala 191:24:@4788.4]
  wire [31:0] x370_sub_1_io_b; // @[Math.scala 191:24:@4788.4]
  wire  x370_sub_1_io_flow; // @[Math.scala 191:24:@4788.4]
  wire [31:0] x370_sub_1_io_result; // @[Math.scala 191:24:@4788.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4798.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4798.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@4798.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@4798.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@4798.4]
  wire  x198_sum_1_clock; // @[Math.scala 150:24:@4807.4]
  wire  x198_sum_1_reset; // @[Math.scala 150:24:@4807.4]
  wire [31:0] x198_sum_1_io_a; // @[Math.scala 150:24:@4807.4]
  wire [31:0] x198_sum_1_io_b; // @[Math.scala 150:24:@4807.4]
  wire  x198_sum_1_io_flow; // @[Math.scala 150:24:@4807.4]
  wire [31:0] x198_sum_1_io_result; // @[Math.scala 150:24:@4807.4]
  wire  x199_sum_1_clock; // @[Math.scala 150:24:@4819.4]
  wire  x199_sum_1_reset; // @[Math.scala 150:24:@4819.4]
  wire [31:0] x199_sum_1_io_a; // @[Math.scala 150:24:@4819.4]
  wire [31:0] x199_sum_1_io_b; // @[Math.scala 150:24:@4819.4]
  wire  x199_sum_1_io_flow; // @[Math.scala 150:24:@4819.4]
  wire [31:0] x199_sum_1_io_result; // @[Math.scala 150:24:@4819.4]
  wire  x372_sum_1_clock; // @[Math.scala 150:24:@4834.4]
  wire  x372_sum_1_reset; // @[Math.scala 150:24:@4834.4]
  wire [31:0] x372_sum_1_io_a; // @[Math.scala 150:24:@4834.4]
  wire [31:0] x372_sum_1_io_b; // @[Math.scala 150:24:@4834.4]
  wire  x372_sum_1_io_flow; // @[Math.scala 150:24:@4834.4]
  wire [31:0] x372_sum_1_io_result; // @[Math.scala 150:24:@4834.4]
  wire [31:0] x202_1_io_b; // @[Math.scala 720:24:@4855.4]
  wire [31:0] x202_1_io_result; // @[Math.scala 720:24:@4855.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@4868.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@4868.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@4868.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@4868.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@4868.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@4877.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@4877.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@4877.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@4877.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@4877.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@4888.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@4888.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@4888.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@4888.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@4888.4]
  wire  _T_327; // @[sm_x206_inr_Foreach.scala 62:18:@4774.4]
  wire  _T_328; // @[sm_x206_inr_Foreach.scala 62:55:@4775.4]
  wire [31:0] b193_number; // @[Math.scala 723:22:@4754.4 Math.scala 724:14:@4755.4]
  wire [42:0] _GEN_0; // @[Math.scala 461:32:@4779.4]
  wire [42:0] _T_331; // @[Math.scala 461:32:@4779.4]
  wire [38:0] _GEN_1; // @[Math.scala 461:32:@4784.4]
  wire [38:0] _T_334; // @[Math.scala 461:32:@4784.4]
  wire [31:0] x199_sum_number; // @[Math.scala 154:22:@4825.4 Math.scala 155:14:@4826.4]
  wire [33:0] _GEN_2; // @[Math.scala 461:32:@4830.4]
  wire [33:0] _T_353; // @[Math.scala 461:32:@4830.4]
  wire [31:0] x372_sum_number; // @[Math.scala 154:22:@4840.4 Math.scala 155:14:@4841.4]
  wire [31:0] _T_364; // @[Math.scala 406:49:@4847.4]
  wire [31:0] _T_366; // @[Math.scala 406:56:@4849.4]
  wire [31:0] _T_367; // @[Math.scala 406:56:@4850.4]
  wire  _T_385; // @[sm_x206_inr_Foreach.scala 93:131:@4885.4]
  wire  _T_389; // @[package.scala 96:25:@4893.4 package.scala 96:25:@4894.4]
  wire  _T_391; // @[implicits.scala 55:10:@4895.4]
  wire  _T_392; // @[sm_x206_inr_Foreach.scala 93:148:@4896.4]
  wire  _T_394; // @[sm_x206_inr_Foreach.scala 93:236:@4898.4]
  wire  _T_395; // @[sm_x206_inr_Foreach.scala 93:255:@4899.4]
  wire  x458_b195_D4; // @[package.scala 96:25:@4873.4 package.scala 96:25:@4874.4]
  wire  _T_398; // @[sm_x206_inr_Foreach.scala 93:291:@4901.4]
  wire  x459_b196_D4; // @[package.scala 96:25:@4882.4 package.scala 96:25:@4883.4]
  _ _ ( // @[Math.scala 720:24:@4749.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@4761.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x370_sub x370_sub_1 ( // @[Math.scala 191:24:@4788.4]
    .clock(x370_sub_1_clock),
    .reset(x370_sub_1_reset),
    .io_a(x370_sub_1_io_a),
    .io_b(x370_sub_1_io_b),
    .io_flow(x370_sub_1_io_flow),
    .io_result(x370_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@4798.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x198_sum x198_sum_1 ( // @[Math.scala 150:24:@4807.4]
    .clock(x198_sum_1_clock),
    .reset(x198_sum_1_reset),
    .io_a(x198_sum_1_io_a),
    .io_b(x198_sum_1_io_b),
    .io_flow(x198_sum_1_io_flow),
    .io_result(x198_sum_1_io_result)
  );
  x198_sum x199_sum_1 ( // @[Math.scala 150:24:@4819.4]
    .clock(x199_sum_1_clock),
    .reset(x199_sum_1_reset),
    .io_a(x199_sum_1_io_a),
    .io_b(x199_sum_1_io_b),
    .io_flow(x199_sum_1_io_flow),
    .io_result(x199_sum_1_io_result)
  );
  x198_sum x372_sum_1 ( // @[Math.scala 150:24:@4834.4]
    .clock(x372_sum_1_clock),
    .reset(x372_sum_1_reset),
    .io_a(x372_sum_1_io_a),
    .io_b(x372_sum_1_io_b),
    .io_flow(x372_sum_1_io_flow),
    .io_result(x372_sum_1_io_result)
  );
  _ x202_1 ( // @[Math.scala 720:24:@4855.4]
    .io_b(x202_1_io_b),
    .io_result(x202_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@4868.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_2 ( // @[package.scala 93:22:@4877.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_3 ( // @[package.scala 93:22:@4888.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_327 = ~ io_in_x188_fifoinpacked_0_full; // @[sm_x206_inr_Foreach.scala 62:18:@4774.4]
  assign _T_328 = ~ io_in_x188_fifoinpacked_0_active_0_out; // @[sm_x206_inr_Foreach.scala 62:55:@4775.4]
  assign b193_number = __io_result; // @[Math.scala 723:22:@4754.4 Math.scala 724:14:@4755.4]
  assign _GEN_0 = {{11'd0}, b193_number}; // @[Math.scala 461:32:@4779.4]
  assign _T_331 = _GEN_0 << 11; // @[Math.scala 461:32:@4779.4]
  assign _GEN_1 = {{7'd0}, b193_number}; // @[Math.scala 461:32:@4784.4]
  assign _T_334 = _GEN_1 << 7; // @[Math.scala 461:32:@4784.4]
  assign x199_sum_number = x199_sum_1_io_result; // @[Math.scala 154:22:@4825.4 Math.scala 155:14:@4826.4]
  assign _GEN_2 = {{2'd0}, x199_sum_number}; // @[Math.scala 461:32:@4830.4]
  assign _T_353 = _GEN_2 << 2; // @[Math.scala 461:32:@4830.4]
  assign x372_sum_number = x372_sum_1_io_result; // @[Math.scala 154:22:@4840.4 Math.scala 155:14:@4841.4]
  assign _T_364 = $signed(x372_sum_number); // @[Math.scala 406:49:@4847.4]
  assign _T_366 = $signed(_T_364) & $signed(32'shff); // @[Math.scala 406:56:@4849.4]
  assign _T_367 = $signed(_T_366); // @[Math.scala 406:56:@4850.4]
  assign _T_385 = ~ io_sigsIn_break; // @[sm_x206_inr_Foreach.scala 93:131:@4885.4]
  assign _T_389 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@4893.4 package.scala 96:25:@4894.4]
  assign _T_391 = io_rr ? _T_389 : 1'h0; // @[implicits.scala 55:10:@4895.4]
  assign _T_392 = _T_385 & _T_391; // @[sm_x206_inr_Foreach.scala 93:148:@4896.4]
  assign _T_394 = _T_392 & _T_385; // @[sm_x206_inr_Foreach.scala 93:236:@4898.4]
  assign _T_395 = _T_394 & io_sigsIn_backpressure; // @[sm_x206_inr_Foreach.scala 93:255:@4899.4]
  assign x458_b195_D4 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@4873.4 package.scala 96:25:@4874.4]
  assign _T_398 = _T_395 & x458_b195_D4; // @[sm_x206_inr_Foreach.scala 93:291:@4901.4]
  assign x459_b196_D4 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@4882.4 package.scala 96:25:@4883.4]
  assign io_in_x188_fifoinpacked_0_wPort_0_en_0 = _T_398 & x459_b196_D4; // @[MemInterfaceType.scala 93:57:@4905.4]
  assign io_in_x188_fifoinpacked_0_active_0_in = x458_b195_D4 & x459_b196_D4; // @[MemInterfaceType.scala 147:18:@4908.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@4752.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@4764.4]
  assign x370_sub_1_clock = clock; // @[:@4789.4]
  assign x370_sub_1_reset = reset; // @[:@4790.4]
  assign x370_sub_1_io_a = _T_331[31:0]; // @[Math.scala 192:17:@4791.4]
  assign x370_sub_1_io_b = _T_334[31:0]; // @[Math.scala 193:17:@4792.4]
  assign x370_sub_1_io_flow = _T_327 | _T_328; // @[Math.scala 194:20:@4793.4]
  assign RetimeWrapper_clock = clock; // @[:@4799.4]
  assign RetimeWrapper_reset = reset; // @[:@4800.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4802.4]
  assign RetimeWrapper_io_in = __1_io_result; // @[package.scala 94:16:@4801.4]
  assign x198_sum_1_clock = clock; // @[:@4808.4]
  assign x198_sum_1_reset = reset; // @[:@4809.4]
  assign x198_sum_1_io_a = x370_sub_1_io_result; // @[Math.scala 151:17:@4810.4]
  assign x198_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@4811.4]
  assign x198_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4812.4]
  assign x199_sum_1_clock = clock; // @[:@4820.4]
  assign x199_sum_1_reset = reset; // @[:@4821.4]
  assign x199_sum_1_io_a = x198_sum_1_io_result; // @[Math.scala 151:17:@4822.4]
  assign x199_sum_1_io_b = 32'h1; // @[Math.scala 152:17:@4823.4]
  assign x199_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4824.4]
  assign x372_sum_1_clock = clock; // @[:@4835.4]
  assign x372_sum_1_reset = reset; // @[:@4836.4]
  assign x372_sum_1_io_a = _T_353[31:0]; // @[Math.scala 151:17:@4837.4]
  assign x372_sum_1_io_b = x199_sum_1_io_result; // @[Math.scala 152:17:@4838.4]
  assign x372_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4839.4]
  assign x202_1_io_b = $unsigned(_T_367); // @[Math.scala 721:17:@4858.4]
  assign RetimeWrapper_1_clock = clock; // @[:@4869.4]
  assign RetimeWrapper_1_reset = reset; // @[:@4870.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4872.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@4871.4]
  assign RetimeWrapper_2_clock = clock; // @[:@4878.4]
  assign RetimeWrapper_2_reset = reset; // @[:@4879.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4881.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@4880.4]
  assign RetimeWrapper_3_clock = clock; // @[:@4889.4]
  assign RetimeWrapper_3_reset = reset; // @[:@4890.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4892.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@4891.4]
endmodule
module RetimeWrapper_42( // @[:@6026.2]
  input   clock, // @[:@6027.4]
  input   reset, // @[:@6028.4]
  input   io_flow, // @[:@6029.4]
  input   io_in, // @[:@6029.4]
  output  io_out // @[:@6029.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6031.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6031.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6031.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6031.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6031.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6031.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(67)) sr ( // @[RetimeShiftRegister.scala 15:20:@6031.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6044.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6043.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6042.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6041.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6040.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6038.4]
endmodule
module RetimeWrapper_46( // @[:@6154.2]
  input   clock, // @[:@6155.4]
  input   reset, // @[:@6156.4]
  input   io_flow, // @[:@6157.4]
  input   io_in, // @[:@6157.4]
  output  io_out // @[:@6157.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6159.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6159.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6159.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6159.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6159.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6159.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(66)) sr ( // @[RetimeShiftRegister.scala 15:20:@6159.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6172.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6171.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6170.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6169.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6168.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6166.4]
endmodule
module x319_inr_Foreach_SAMPLER_BOX_sm( // @[:@6174.2]
  input   clock, // @[:@6175.4]
  input   reset, // @[:@6176.4]
  input   io_enable, // @[:@6177.4]
  output  io_done, // @[:@6177.4]
  output  io_doneLatch, // @[:@6177.4]
  input   io_ctrDone, // @[:@6177.4]
  output  io_datapathEn, // @[:@6177.4]
  output  io_ctrInc, // @[:@6177.4]
  output  io_ctrRst, // @[:@6177.4]
  input   io_parentAck, // @[:@6177.4]
  input   io_backpressure, // @[:@6177.4]
  input   io_break // @[:@6177.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@6179.4]
  wire  active_reset; // @[Controllers.scala 261:22:@6179.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@6179.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@6179.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@6179.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@6179.4]
  wire  done_clock; // @[Controllers.scala 262:20:@6182.4]
  wire  done_reset; // @[Controllers.scala 262:20:@6182.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@6182.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@6182.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@6182.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@6182.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6216.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6216.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6216.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@6216.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@6216.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6238.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6238.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6238.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6238.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6238.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6250.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6250.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6250.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6250.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6250.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6258.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6258.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6258.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6258.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6258.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@6274.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@6274.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@6274.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@6274.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@6274.4]
  wire  _T_80; // @[Controllers.scala 264:48:@6187.4]
  wire  _T_81; // @[Controllers.scala 264:46:@6188.4]
  wire  _T_82; // @[Controllers.scala 264:62:@6189.4]
  wire  _T_83; // @[Controllers.scala 264:60:@6190.4]
  wire  _T_100; // @[package.scala 100:49:@6207.4]
  reg  _T_103; // @[package.scala 48:56:@6208.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@6221.4 package.scala 96:25:@6222.4]
  wire  _T_110; // @[package.scala 100:49:@6223.4]
  reg  _T_113; // @[package.scala 48:56:@6224.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@6226.4]
  wire  _T_118; // @[Controllers.scala 283:41:@6231.4]
  wire  _T_119; // @[Controllers.scala 283:59:@6232.4]
  wire  _T_121; // @[Controllers.scala 284:37:@6235.4]
  wire  _T_124; // @[package.scala 96:25:@6243.4 package.scala 96:25:@6244.4]
  wire  _T_126; // @[package.scala 100:49:@6245.4]
  reg  _T_129; // @[package.scala 48:56:@6246.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@6268.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@6270.4]
  reg  _T_153; // @[package.scala 48:56:@6271.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@6279.4 package.scala 96:25:@6280.4]
  wire  _T_158; // @[Controllers.scala 292:61:@6281.4]
  wire  _T_159; // @[Controllers.scala 292:24:@6282.4]
  SRFF active ( // @[Controllers.scala 261:22:@6179.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@6182.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_42 RetimeWrapper ( // @[package.scala 93:22:@6216.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_42 RetimeWrapper_1 ( // @[package.scala 93:22:@6238.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@6250.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@6258.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_46 RetimeWrapper_4 ( // @[package.scala 93:22:@6274.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@6187.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@6188.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@6189.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@6190.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@6207.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@6221.4 package.scala 96:25:@6222.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@6223.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@6226.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@6231.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@6232.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@6235.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6243.4 package.scala 96:25:@6244.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@6245.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@6270.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@6279.4 package.scala 96:25:@6280.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@6281.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@6282.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@6249.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@6284.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@6234.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@6237.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@6229.4]
  assign active_clock = clock; // @[:@6180.4]
  assign active_reset = reset; // @[:@6181.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@6192.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@6196.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@6197.4]
  assign done_clock = clock; // @[:@6183.4]
  assign done_reset = reset; // @[:@6184.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@6212.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@6205.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@6206.4]
  assign RetimeWrapper_clock = clock; // @[:@6217.4]
  assign RetimeWrapper_reset = reset; // @[:@6218.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@6220.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@6219.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6239.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6240.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@6242.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@6241.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6251.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6252.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@6254.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@6253.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6259.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6260.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@6262.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@6261.4]
  assign RetimeWrapper_4_clock = clock; // @[:@6275.4]
  assign RetimeWrapper_4_reset = reset; // @[:@6276.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@6278.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@6277.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SRAM_1( // @[:@6511.2]
  input         clock, // @[:@6512.4]
  input         reset, // @[:@6513.4]
  input  [9:0]  io_raddr, // @[:@6514.4]
  input         io_wen, // @[:@6514.4]
  input  [9:0]  io_waddr, // @[:@6514.4]
  input  [31:0] io_wdata, // @[:@6514.4]
  output [31:0] io_rdata, // @[:@6514.4]
  input         io_backpressure // @[:@6514.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@6516.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@6516.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@6516.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@6516.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@6516.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@6516.4]
  wire [9:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@6516.4]
  wire [9:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@6516.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@6516.4]
  wire  _T_19; // @[SRAM.scala 182:49:@6534.4]
  wire  _T_20; // @[SRAM.scala 182:37:@6535.4]
  reg  _T_23; // @[SRAM.scala 182:29:@6536.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@6538.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(640), .AWIDTH(10)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@6516.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@6534.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@6535.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@6543.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@6530.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@6531.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@6528.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@6533.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@6532.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@6529.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@6527.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@6526.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module RetimeWrapper_51( // @[:@6557.2]
  input        clock, // @[:@6558.4]
  input        reset, // @[:@6559.4]
  input        io_flow, // @[:@6560.4]
  input  [9:0] io_in, // @[:@6560.4]
  output [9:0] io_out // @[:@6560.4]
);
  wire [9:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@6562.4]
  wire [9:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@6562.4]
  wire [9:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@6562.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6562.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6562.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6562.4]
  RetimeShiftRegister #(.WIDTH(10), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@6562.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6575.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6574.4]
  assign sr_init = 10'h0; // @[RetimeShiftRegister.scala 19:16:@6573.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6572.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6571.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6569.4]
endmodule
module Mem1D_5( // @[:@6577.2]
  input         clock, // @[:@6578.4]
  input         reset, // @[:@6579.4]
  input  [9:0]  io_r_ofs_0, // @[:@6580.4]
  input         io_r_backpressure, // @[:@6580.4]
  input  [9:0]  io_w_ofs_0, // @[:@6580.4]
  input  [31:0] io_w_data_0, // @[:@6580.4]
  input         io_w_en_0, // @[:@6580.4]
  output [31:0] io_output // @[:@6580.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@6584.4]
  wire  SRAM_reset; // @[MemPrimitives.scala 715:21:@6584.4]
  wire [9:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@6584.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 715:21:@6584.4]
  wire [9:0] SRAM_io_waddr; // @[MemPrimitives.scala 715:21:@6584.4]
  wire [31:0] SRAM_io_wdata; // @[MemPrimitives.scala 715:21:@6584.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@6584.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@6584.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6587.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6587.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6587.4]
  wire [9:0] RetimeWrapper_io_in; // @[package.scala 93:22:@6587.4]
  wire [9:0] RetimeWrapper_io_out; // @[package.scala 93:22:@6587.4]
  wire  wInBound; // @[MemPrimitives.scala 702:32:@6582.4]
  SRAM_1 SRAM ( // @[MemPrimitives.scala 715:21:@6584.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_51 RetimeWrapper ( // @[package.scala 93:22:@6587.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 10'h280; // @[MemPrimitives.scala 702:32:@6582.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@6600.4]
  assign SRAM_clock = clock; // @[:@6585.4]
  assign SRAM_reset = reset; // @[:@6586.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@6594.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 719:22:@6597.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 718:22:@6595.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 720:22:@6598.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@6599.4]
  assign RetimeWrapper_clock = clock; // @[:@6588.4]
  assign RetimeWrapper_reset = reset; // @[:@6589.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@6591.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@6590.4]
endmodule
module StickySelects_1( // @[:@7779.2]
  input   clock, // @[:@7780.4]
  input   reset, // @[:@7781.4]
  input   io_ins_0, // @[:@7782.4]
  input   io_ins_1, // @[:@7782.4]
  input   io_ins_2, // @[:@7782.4]
  input   io_ins_3, // @[:@7782.4]
  input   io_ins_4, // @[:@7782.4]
  input   io_ins_5, // @[:@7782.4]
  input   io_ins_6, // @[:@7782.4]
  input   io_ins_7, // @[:@7782.4]
  input   io_ins_8, // @[:@7782.4]
  output  io_outs_0, // @[:@7782.4]
  output  io_outs_1, // @[:@7782.4]
  output  io_outs_2, // @[:@7782.4]
  output  io_outs_3, // @[:@7782.4]
  output  io_outs_4, // @[:@7782.4]
  output  io_outs_5, // @[:@7782.4]
  output  io_outs_6, // @[:@7782.4]
  output  io_outs_7, // @[:@7782.4]
  output  io_outs_8 // @[:@7782.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@7784.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@7785.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@7786.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@7787.4]
  reg [31:0] _RAND_3;
  reg  _T_31; // @[StickySelects.scala 37:46:@7788.4]
  reg [31:0] _RAND_4;
  reg  _T_34; // @[StickySelects.scala 37:46:@7789.4]
  reg [31:0] _RAND_5;
  reg  _T_37; // @[StickySelects.scala 37:46:@7790.4]
  reg [31:0] _RAND_6;
  reg  _T_40; // @[StickySelects.scala 37:46:@7791.4]
  reg [31:0] _RAND_7;
  reg  _T_43; // @[StickySelects.scala 37:46:@7792.4]
  reg [31:0] _RAND_8;
  wire  _T_44; // @[StickySelects.scala 47:46:@7793.4]
  wire  _T_45; // @[StickySelects.scala 47:46:@7794.4]
  wire  _T_46; // @[StickySelects.scala 47:46:@7795.4]
  wire  _T_47; // @[StickySelects.scala 47:46:@7796.4]
  wire  _T_48; // @[StickySelects.scala 47:46:@7797.4]
  wire  _T_49; // @[StickySelects.scala 47:46:@7798.4]
  wire  _T_50; // @[StickySelects.scala 47:46:@7799.4]
  wire  _T_51; // @[StickySelects.scala 49:53:@7800.4]
  wire  _T_52; // @[StickySelects.scala 49:21:@7801.4]
  wire  _T_53; // @[StickySelects.scala 47:46:@7803.4]
  wire  _T_54; // @[StickySelects.scala 47:46:@7804.4]
  wire  _T_55; // @[StickySelects.scala 47:46:@7805.4]
  wire  _T_56; // @[StickySelects.scala 47:46:@7806.4]
  wire  _T_57; // @[StickySelects.scala 47:46:@7807.4]
  wire  _T_58; // @[StickySelects.scala 47:46:@7808.4]
  wire  _T_59; // @[StickySelects.scala 47:46:@7809.4]
  wire  _T_60; // @[StickySelects.scala 49:53:@7810.4]
  wire  _T_61; // @[StickySelects.scala 49:21:@7811.4]
  wire  _T_62; // @[StickySelects.scala 47:46:@7813.4]
  wire  _T_63; // @[StickySelects.scala 47:46:@7814.4]
  wire  _T_64; // @[StickySelects.scala 47:46:@7815.4]
  wire  _T_65; // @[StickySelects.scala 47:46:@7816.4]
  wire  _T_66; // @[StickySelects.scala 47:46:@7817.4]
  wire  _T_67; // @[StickySelects.scala 47:46:@7818.4]
  wire  _T_68; // @[StickySelects.scala 47:46:@7819.4]
  wire  _T_69; // @[StickySelects.scala 49:53:@7820.4]
  wire  _T_70; // @[StickySelects.scala 49:21:@7821.4]
  wire  _T_72; // @[StickySelects.scala 47:46:@7824.4]
  wire  _T_73; // @[StickySelects.scala 47:46:@7825.4]
  wire  _T_74; // @[StickySelects.scala 47:46:@7826.4]
  wire  _T_75; // @[StickySelects.scala 47:46:@7827.4]
  wire  _T_76; // @[StickySelects.scala 47:46:@7828.4]
  wire  _T_77; // @[StickySelects.scala 47:46:@7829.4]
  wire  _T_78; // @[StickySelects.scala 49:53:@7830.4]
  wire  _T_79; // @[StickySelects.scala 49:21:@7831.4]
  wire  _T_82; // @[StickySelects.scala 47:46:@7835.4]
  wire  _T_83; // @[StickySelects.scala 47:46:@7836.4]
  wire  _T_84; // @[StickySelects.scala 47:46:@7837.4]
  wire  _T_85; // @[StickySelects.scala 47:46:@7838.4]
  wire  _T_86; // @[StickySelects.scala 47:46:@7839.4]
  wire  _T_87; // @[StickySelects.scala 49:53:@7840.4]
  wire  _T_88; // @[StickySelects.scala 49:21:@7841.4]
  wire  _T_92; // @[StickySelects.scala 47:46:@7846.4]
  wire  _T_93; // @[StickySelects.scala 47:46:@7847.4]
  wire  _T_94; // @[StickySelects.scala 47:46:@7848.4]
  wire  _T_95; // @[StickySelects.scala 47:46:@7849.4]
  wire  _T_96; // @[StickySelects.scala 49:53:@7850.4]
  wire  _T_97; // @[StickySelects.scala 49:21:@7851.4]
  wire  _T_102; // @[StickySelects.scala 47:46:@7857.4]
  wire  _T_103; // @[StickySelects.scala 47:46:@7858.4]
  wire  _T_104; // @[StickySelects.scala 47:46:@7859.4]
  wire  _T_105; // @[StickySelects.scala 49:53:@7860.4]
  wire  _T_106; // @[StickySelects.scala 49:21:@7861.4]
  wire  _T_112; // @[StickySelects.scala 47:46:@7868.4]
  wire  _T_113; // @[StickySelects.scala 47:46:@7869.4]
  wire  _T_114; // @[StickySelects.scala 49:53:@7870.4]
  wire  _T_115; // @[StickySelects.scala 49:21:@7871.4]
  wire  _T_122; // @[StickySelects.scala 47:46:@7879.4]
  wire  _T_123; // @[StickySelects.scala 49:53:@7880.4]
  wire  _T_124; // @[StickySelects.scala 49:21:@7881.4]
  assign _T_44 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@7793.4]
  assign _T_45 = _T_44 | io_ins_3; // @[StickySelects.scala 47:46:@7794.4]
  assign _T_46 = _T_45 | io_ins_4; // @[StickySelects.scala 47:46:@7795.4]
  assign _T_47 = _T_46 | io_ins_5; // @[StickySelects.scala 47:46:@7796.4]
  assign _T_48 = _T_47 | io_ins_6; // @[StickySelects.scala 47:46:@7797.4]
  assign _T_49 = _T_48 | io_ins_7; // @[StickySelects.scala 47:46:@7798.4]
  assign _T_50 = _T_49 | io_ins_8; // @[StickySelects.scala 47:46:@7799.4]
  assign _T_51 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@7800.4]
  assign _T_52 = _T_50 ? io_ins_0 : _T_51; // @[StickySelects.scala 49:21:@7801.4]
  assign _T_53 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@7803.4]
  assign _T_54 = _T_53 | io_ins_3; // @[StickySelects.scala 47:46:@7804.4]
  assign _T_55 = _T_54 | io_ins_4; // @[StickySelects.scala 47:46:@7805.4]
  assign _T_56 = _T_55 | io_ins_5; // @[StickySelects.scala 47:46:@7806.4]
  assign _T_57 = _T_56 | io_ins_6; // @[StickySelects.scala 47:46:@7807.4]
  assign _T_58 = _T_57 | io_ins_7; // @[StickySelects.scala 47:46:@7808.4]
  assign _T_59 = _T_58 | io_ins_8; // @[StickySelects.scala 47:46:@7809.4]
  assign _T_60 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@7810.4]
  assign _T_61 = _T_59 ? io_ins_1 : _T_60; // @[StickySelects.scala 49:21:@7811.4]
  assign _T_62 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@7813.4]
  assign _T_63 = _T_62 | io_ins_3; // @[StickySelects.scala 47:46:@7814.4]
  assign _T_64 = _T_63 | io_ins_4; // @[StickySelects.scala 47:46:@7815.4]
  assign _T_65 = _T_64 | io_ins_5; // @[StickySelects.scala 47:46:@7816.4]
  assign _T_66 = _T_65 | io_ins_6; // @[StickySelects.scala 47:46:@7817.4]
  assign _T_67 = _T_66 | io_ins_7; // @[StickySelects.scala 47:46:@7818.4]
  assign _T_68 = _T_67 | io_ins_8; // @[StickySelects.scala 47:46:@7819.4]
  assign _T_69 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@7820.4]
  assign _T_70 = _T_68 ? io_ins_2 : _T_69; // @[StickySelects.scala 49:21:@7821.4]
  assign _T_72 = _T_62 | io_ins_2; // @[StickySelects.scala 47:46:@7824.4]
  assign _T_73 = _T_72 | io_ins_4; // @[StickySelects.scala 47:46:@7825.4]
  assign _T_74 = _T_73 | io_ins_5; // @[StickySelects.scala 47:46:@7826.4]
  assign _T_75 = _T_74 | io_ins_6; // @[StickySelects.scala 47:46:@7827.4]
  assign _T_76 = _T_75 | io_ins_7; // @[StickySelects.scala 47:46:@7828.4]
  assign _T_77 = _T_76 | io_ins_8; // @[StickySelects.scala 47:46:@7829.4]
  assign _T_78 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@7830.4]
  assign _T_79 = _T_77 ? io_ins_3 : _T_78; // @[StickySelects.scala 49:21:@7831.4]
  assign _T_82 = _T_72 | io_ins_3; // @[StickySelects.scala 47:46:@7835.4]
  assign _T_83 = _T_82 | io_ins_5; // @[StickySelects.scala 47:46:@7836.4]
  assign _T_84 = _T_83 | io_ins_6; // @[StickySelects.scala 47:46:@7837.4]
  assign _T_85 = _T_84 | io_ins_7; // @[StickySelects.scala 47:46:@7838.4]
  assign _T_86 = _T_85 | io_ins_8; // @[StickySelects.scala 47:46:@7839.4]
  assign _T_87 = io_ins_4 | _T_31; // @[StickySelects.scala 49:53:@7840.4]
  assign _T_88 = _T_86 ? io_ins_4 : _T_87; // @[StickySelects.scala 49:21:@7841.4]
  assign _T_92 = _T_82 | io_ins_4; // @[StickySelects.scala 47:46:@7846.4]
  assign _T_93 = _T_92 | io_ins_6; // @[StickySelects.scala 47:46:@7847.4]
  assign _T_94 = _T_93 | io_ins_7; // @[StickySelects.scala 47:46:@7848.4]
  assign _T_95 = _T_94 | io_ins_8; // @[StickySelects.scala 47:46:@7849.4]
  assign _T_96 = io_ins_5 | _T_34; // @[StickySelects.scala 49:53:@7850.4]
  assign _T_97 = _T_95 ? io_ins_5 : _T_96; // @[StickySelects.scala 49:21:@7851.4]
  assign _T_102 = _T_92 | io_ins_5; // @[StickySelects.scala 47:46:@7857.4]
  assign _T_103 = _T_102 | io_ins_7; // @[StickySelects.scala 47:46:@7858.4]
  assign _T_104 = _T_103 | io_ins_8; // @[StickySelects.scala 47:46:@7859.4]
  assign _T_105 = io_ins_6 | _T_37; // @[StickySelects.scala 49:53:@7860.4]
  assign _T_106 = _T_104 ? io_ins_6 : _T_105; // @[StickySelects.scala 49:21:@7861.4]
  assign _T_112 = _T_102 | io_ins_6; // @[StickySelects.scala 47:46:@7868.4]
  assign _T_113 = _T_112 | io_ins_8; // @[StickySelects.scala 47:46:@7869.4]
  assign _T_114 = io_ins_7 | _T_40; // @[StickySelects.scala 49:53:@7870.4]
  assign _T_115 = _T_113 ? io_ins_7 : _T_114; // @[StickySelects.scala 49:21:@7871.4]
  assign _T_122 = _T_112 | io_ins_7; // @[StickySelects.scala 47:46:@7879.4]
  assign _T_123 = io_ins_8 | _T_43; // @[StickySelects.scala 49:53:@7880.4]
  assign _T_124 = _T_122 ? io_ins_8 : _T_123; // @[StickySelects.scala 49:21:@7881.4]
  assign io_outs_0 = _T_50 ? io_ins_0 : _T_51; // @[StickySelects.scala 53:57:@7883.4]
  assign io_outs_1 = _T_59 ? io_ins_1 : _T_60; // @[StickySelects.scala 53:57:@7884.4]
  assign io_outs_2 = _T_68 ? io_ins_2 : _T_69; // @[StickySelects.scala 53:57:@7885.4]
  assign io_outs_3 = _T_77 ? io_ins_3 : _T_78; // @[StickySelects.scala 53:57:@7886.4]
  assign io_outs_4 = _T_86 ? io_ins_4 : _T_87; // @[StickySelects.scala 53:57:@7887.4]
  assign io_outs_5 = _T_95 ? io_ins_5 : _T_96; // @[StickySelects.scala 53:57:@7888.4]
  assign io_outs_6 = _T_104 ? io_ins_6 : _T_105; // @[StickySelects.scala 53:57:@7889.4]
  assign io_outs_7 = _T_113 ? io_ins_7 : _T_114; // @[StickySelects.scala 53:57:@7890.4]
  assign io_outs_8 = _T_122 ? io_ins_8 : _T_123; // @[StickySelects.scala 53:57:@7891.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_31 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_37 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_40 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_43 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_50) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_51;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_59) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_60;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_68) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_69;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_77) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_78;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_86) begin
        _T_31 <= io_ins_4;
      end else begin
        _T_31 <= _T_87;
      end
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (_T_95) begin
        _T_34 <= io_ins_5;
      end else begin
        _T_34 <= _T_96;
      end
    end
    if (reset) begin
      _T_37 <= 1'h0;
    end else begin
      if (_T_104) begin
        _T_37 <= io_ins_6;
      end else begin
        _T_37 <= _T_105;
      end
    end
    if (reset) begin
      _T_40 <= 1'h0;
    end else begin
      if (_T_113) begin
        _T_40 <= io_ins_7;
      end else begin
        _T_40 <= _T_114;
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_122) begin
        _T_43 <= io_ins_8;
      end else begin
        _T_43 <= _T_123;
      end
    end
  end
endmodule
module x217_lb_0( // @[:@12603.2]
  input         clock, // @[:@12604.4]
  input         reset, // @[:@12605.4]
  input  [1:0]  io_rPort_8_banks_1, // @[:@12606.4]
  input  [2:0]  io_rPort_8_banks_0, // @[:@12606.4]
  input  [9:0]  io_rPort_8_ofs_0, // @[:@12606.4]
  input         io_rPort_8_en_0, // @[:@12606.4]
  input         io_rPort_8_backpressure, // @[:@12606.4]
  output [31:0] io_rPort_8_output_0, // @[:@12606.4]
  input  [1:0]  io_rPort_7_banks_1, // @[:@12606.4]
  input  [2:0]  io_rPort_7_banks_0, // @[:@12606.4]
  input  [9:0]  io_rPort_7_ofs_0, // @[:@12606.4]
  input         io_rPort_7_en_0, // @[:@12606.4]
  input         io_rPort_7_backpressure, // @[:@12606.4]
  output [31:0] io_rPort_7_output_0, // @[:@12606.4]
  input  [1:0]  io_rPort_6_banks_1, // @[:@12606.4]
  input  [2:0]  io_rPort_6_banks_0, // @[:@12606.4]
  input  [9:0]  io_rPort_6_ofs_0, // @[:@12606.4]
  input         io_rPort_6_en_0, // @[:@12606.4]
  input         io_rPort_6_backpressure, // @[:@12606.4]
  output [31:0] io_rPort_6_output_0, // @[:@12606.4]
  input  [1:0]  io_rPort_5_banks_1, // @[:@12606.4]
  input  [2:0]  io_rPort_5_banks_0, // @[:@12606.4]
  input  [9:0]  io_rPort_5_ofs_0, // @[:@12606.4]
  input         io_rPort_5_en_0, // @[:@12606.4]
  input         io_rPort_5_backpressure, // @[:@12606.4]
  output [31:0] io_rPort_5_output_0, // @[:@12606.4]
  input  [1:0]  io_rPort_4_banks_1, // @[:@12606.4]
  input  [2:0]  io_rPort_4_banks_0, // @[:@12606.4]
  input  [9:0]  io_rPort_4_ofs_0, // @[:@12606.4]
  input         io_rPort_4_en_0, // @[:@12606.4]
  input         io_rPort_4_backpressure, // @[:@12606.4]
  output [31:0] io_rPort_4_output_0, // @[:@12606.4]
  input  [1:0]  io_rPort_3_banks_1, // @[:@12606.4]
  input  [2:0]  io_rPort_3_banks_0, // @[:@12606.4]
  input  [9:0]  io_rPort_3_ofs_0, // @[:@12606.4]
  input         io_rPort_3_en_0, // @[:@12606.4]
  input         io_rPort_3_backpressure, // @[:@12606.4]
  output [31:0] io_rPort_3_output_0, // @[:@12606.4]
  input  [1:0]  io_rPort_2_banks_1, // @[:@12606.4]
  input  [2:0]  io_rPort_2_banks_0, // @[:@12606.4]
  input  [9:0]  io_rPort_2_ofs_0, // @[:@12606.4]
  input         io_rPort_2_en_0, // @[:@12606.4]
  input         io_rPort_2_backpressure, // @[:@12606.4]
  output [31:0] io_rPort_2_output_0, // @[:@12606.4]
  input  [1:0]  io_rPort_1_banks_1, // @[:@12606.4]
  input  [2:0]  io_rPort_1_banks_0, // @[:@12606.4]
  input  [9:0]  io_rPort_1_ofs_0, // @[:@12606.4]
  input         io_rPort_1_en_0, // @[:@12606.4]
  input         io_rPort_1_backpressure, // @[:@12606.4]
  output [31:0] io_rPort_1_output_0, // @[:@12606.4]
  input  [1:0]  io_rPort_0_banks_1, // @[:@12606.4]
  input  [2:0]  io_rPort_0_banks_0, // @[:@12606.4]
  input  [9:0]  io_rPort_0_ofs_0, // @[:@12606.4]
  input         io_rPort_0_en_0, // @[:@12606.4]
  input         io_rPort_0_backpressure, // @[:@12606.4]
  output [31:0] io_rPort_0_output_0, // @[:@12606.4]
  input  [1:0]  io_wPort_0_banks_1, // @[:@12606.4]
  input  [2:0]  io_wPort_0_banks_0, // @[:@12606.4]
  input  [9:0]  io_wPort_0_ofs_0, // @[:@12606.4]
  input  [31:0] io_wPort_0_data_0, // @[:@12606.4]
  input         io_wPort_0_en_0 // @[:@12606.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@12671.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@12671.4]
  wire [9:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12671.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12671.4]
  wire [9:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12671.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@12671.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@12671.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@12671.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@12687.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@12687.4]
  wire [9:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12687.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12687.4]
  wire [9:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12687.4]
  wire [31:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@12687.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@12687.4]
  wire [31:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@12687.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@12703.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@12703.4]
  wire [9:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12703.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12703.4]
  wire [9:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12703.4]
  wire [31:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@12703.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@12703.4]
  wire [31:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@12703.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@12719.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@12719.4]
  wire [9:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12719.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12719.4]
  wire [9:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12719.4]
  wire [31:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@12719.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@12719.4]
  wire [31:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@12719.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@12735.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@12735.4]
  wire [9:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12735.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12735.4]
  wire [9:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12735.4]
  wire [31:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@12735.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@12735.4]
  wire [31:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@12735.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@12751.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@12751.4]
  wire [9:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12751.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12751.4]
  wire [9:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12751.4]
  wire [31:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@12751.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@12751.4]
  wire [31:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@12751.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@12767.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@12767.4]
  wire [9:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12767.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12767.4]
  wire [9:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12767.4]
  wire [31:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@12767.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@12767.4]
  wire [31:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@12767.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@12783.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@12783.4]
  wire [9:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12783.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12783.4]
  wire [9:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12783.4]
  wire [31:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@12783.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@12783.4]
  wire [31:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@12783.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@12799.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@12799.4]
  wire [9:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12799.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12799.4]
  wire [9:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12799.4]
  wire [31:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@12799.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@12799.4]
  wire [31:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@12799.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@12815.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@12815.4]
  wire [9:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12815.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12815.4]
  wire [9:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12815.4]
  wire [31:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@12815.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@12815.4]
  wire [31:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@12815.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@12831.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@12831.4]
  wire [9:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12831.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12831.4]
  wire [9:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12831.4]
  wire [31:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@12831.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@12831.4]
  wire [31:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@12831.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@12847.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@12847.4]
  wire [9:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12847.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12847.4]
  wire [9:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12847.4]
  wire [31:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@12847.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@12847.4]
  wire [31:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@12847.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_ins_6; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_ins_7; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_ins_8; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_outs_6; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_outs_7; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_io_outs_8; // @[MemPrimitives.scala 124:33:@13043.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_ins_6; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_ins_7; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_ins_8; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_outs_6; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_outs_7; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_1_io_outs_8; // @[MemPrimitives.scala 124:33:@13132.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_ins_6; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_ins_7; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_ins_8; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_outs_6; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_outs_7; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_2_io_outs_8; // @[MemPrimitives.scala 124:33:@13221.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_ins_6; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_ins_7; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_ins_8; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_outs_6; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_outs_7; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_3_io_outs_8; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_ins_6; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_ins_7; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_ins_8; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_outs_6; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_outs_7; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_4_io_outs_8; // @[MemPrimitives.scala 124:33:@13399.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_ins_6; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_ins_7; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_ins_8; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_outs_6; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_outs_7; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_5_io_outs_8; // @[MemPrimitives.scala 124:33:@13488.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_ins_6; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_ins_7; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_ins_8; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_outs_6; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_outs_7; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_6_io_outs_8; // @[MemPrimitives.scala 124:33:@13577.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_ins_6; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_ins_7; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_ins_8; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_outs_6; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_outs_7; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_7_io_outs_8; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_ins_6; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_ins_7; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_ins_8; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_outs_6; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_outs_7; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_8_io_outs_8; // @[MemPrimitives.scala 124:33:@13755.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_ins_6; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_ins_7; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_ins_8; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_outs_6; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_outs_7; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_9_io_outs_8; // @[MemPrimitives.scala 124:33:@13844.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_ins_6; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_ins_7; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_ins_8; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_outs_6; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_outs_7; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_10_io_outs_8; // @[MemPrimitives.scala 124:33:@13933.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_ins_6; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_ins_7; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_ins_8; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_outs_6; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_outs_7; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  StickySelects_11_io_outs_8; // @[MemPrimitives.scala 124:33:@14022.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@14112.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@14112.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@14112.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@14112.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@14112.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@14120.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@14120.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@14120.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@14120.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@14120.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@14128.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@14128.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@14128.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@14128.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@14128.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@14136.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@14136.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@14136.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@14136.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@14136.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@14144.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@14144.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@14144.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@14144.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@14144.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@14152.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@14152.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@14152.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@14152.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@14152.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@14160.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@14160.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@14160.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@14160.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@14160.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@14168.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@14168.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@14168.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@14168.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@14168.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@14176.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@14176.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@14176.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@14176.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@14176.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@14184.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@14184.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@14184.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@14184.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@14184.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@14192.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@14192.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@14192.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@14192.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@14192.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@14200.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@14200.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@14200.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@14200.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@14200.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@14256.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@14256.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@14256.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@14256.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@14256.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@14264.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@14264.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@14264.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@14264.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@14264.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@14272.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@14272.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@14272.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@14272.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@14272.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@14280.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@14280.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@14280.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@14280.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@14280.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@14288.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@14288.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@14288.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@14288.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@14288.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@14296.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@14296.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@14296.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@14296.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@14296.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@14304.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@14304.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@14304.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@14304.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@14304.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@14312.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@14312.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@14312.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@14312.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@14312.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@14320.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@14320.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@14320.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@14320.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@14320.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@14328.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@14328.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@14328.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@14328.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@14328.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@14336.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@14336.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@14336.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@14336.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@14336.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@14344.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@14344.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@14344.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@14344.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@14344.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@14400.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@14400.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@14400.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@14400.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@14400.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@14408.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@14408.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@14408.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@14408.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@14408.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@14416.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@14416.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@14416.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@14416.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@14416.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@14424.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@14424.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@14424.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@14424.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@14424.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@14432.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@14432.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@14432.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@14432.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@14432.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@14440.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@14440.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@14440.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@14440.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@14440.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@14448.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@14448.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@14448.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@14448.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@14448.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@14456.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@14456.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@14456.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@14456.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@14456.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@14464.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@14464.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@14464.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@14464.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@14464.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@14472.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@14472.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@14472.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@14472.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@14472.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@14480.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@14480.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@14480.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@14480.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@14480.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@14488.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@14488.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@14488.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@14488.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@14488.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@14544.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@14544.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@14544.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@14544.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@14544.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@14552.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@14552.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@14552.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@14552.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@14552.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@14560.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@14560.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@14560.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@14560.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@14560.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@14568.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@14568.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@14568.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@14568.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@14568.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@14576.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@14576.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@14576.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@14576.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@14576.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@14584.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@14584.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@14584.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@14584.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@14584.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@14592.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@14592.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@14592.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@14592.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@14592.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@14600.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@14600.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@14600.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@14600.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@14600.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@14608.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@14608.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@14608.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@14608.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@14608.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@14616.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@14616.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@14616.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@14616.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@14616.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@14624.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@14624.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@14624.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@14624.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@14624.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@14632.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@14632.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@14632.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@14632.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@14632.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@14688.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@14688.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@14688.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@14688.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@14688.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@14696.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@14696.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@14696.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@14696.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@14696.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@14704.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@14704.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@14704.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@14704.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@14704.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@14712.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@14712.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@14712.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@14712.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@14712.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@14720.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@14720.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@14720.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@14720.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@14720.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@14728.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@14728.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@14728.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@14728.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@14728.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@14736.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@14736.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@14736.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@14736.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@14736.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@14744.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@14744.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@14744.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@14744.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@14744.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@14752.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@14752.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@14752.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@14752.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@14752.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@14760.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@14760.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@14760.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@14760.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@14760.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@14768.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@14768.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@14768.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@14768.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@14768.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@14776.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@14776.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@14776.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@14776.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@14776.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@14832.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@14832.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@14832.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@14832.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@14832.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@14840.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@14840.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@14840.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@14840.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@14840.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@14848.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@14848.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@14848.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@14848.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@14848.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@14856.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@14856.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@14856.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@14856.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@14856.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@14864.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@14864.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@14864.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@14864.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@14864.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@14872.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@14872.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@14872.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@14872.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@14872.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@14880.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@14880.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@14880.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@14880.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@14880.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@14888.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@14888.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@14888.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@14888.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@14888.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@14896.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@14896.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@14896.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@14896.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@14896.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@14904.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@14904.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@14904.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@14904.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@14904.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@14912.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@14912.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@14912.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@14912.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@14912.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@14920.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@14920.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@14920.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@14920.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@14920.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@14976.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@14976.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@14976.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@14976.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@14976.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@14984.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@14984.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@14984.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@14984.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@14984.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@14992.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@14992.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@14992.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@14992.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@14992.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@15000.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@15000.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@15000.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@15000.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@15000.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@15008.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@15008.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@15008.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@15008.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@15008.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@15016.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@15016.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@15016.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@15016.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@15016.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@15024.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@15024.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@15024.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@15024.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@15024.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@15032.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@15032.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@15032.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@15032.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@15032.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@15040.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@15040.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@15040.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@15040.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@15040.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@15048.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@15048.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@15048.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@15048.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@15048.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@15056.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@15056.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@15056.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@15056.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@15056.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@15064.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@15064.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@15064.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@15064.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@15064.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@15120.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@15120.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@15120.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@15120.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@15120.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@15128.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@15128.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@15128.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@15128.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@15128.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@15136.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@15136.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@15136.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@15136.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@15136.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@15144.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@15144.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@15144.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@15144.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@15144.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@15152.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@15152.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@15152.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@15152.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@15152.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@15160.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@15160.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@15160.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@15160.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@15160.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@15168.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@15168.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@15168.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@15168.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@15168.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@15176.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@15176.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@15176.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@15176.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@15176.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@15184.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@15184.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@15184.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@15184.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@15184.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@15192.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@15192.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@15192.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@15192.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@15192.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@15200.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@15200.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@15200.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@15200.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@15200.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@15208.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@15208.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@15208.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@15208.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@15208.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@15264.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@15264.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@15264.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@15264.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@15264.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@15272.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@15272.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@15272.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@15272.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@15272.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@15280.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@15280.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@15280.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@15280.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@15280.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@15288.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@15288.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@15288.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@15288.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@15288.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@15296.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@15296.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@15296.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@15296.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@15296.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@15304.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@15304.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@15304.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@15304.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@15304.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@15312.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@15312.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@15312.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@15312.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@15312.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@15320.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@15320.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@15320.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@15320.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@15320.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@15328.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@15328.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@15328.4]
  wire  RetimeWrapper_104_io_in; // @[package.scala 93:22:@15328.4]
  wire  RetimeWrapper_104_io_out; // @[package.scala 93:22:@15328.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@15336.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@15336.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@15336.4]
  wire  RetimeWrapper_105_io_in; // @[package.scala 93:22:@15336.4]
  wire  RetimeWrapper_105_io_out; // @[package.scala 93:22:@15336.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@15344.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@15344.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@15344.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@15344.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@15344.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@15352.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@15352.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@15352.4]
  wire  RetimeWrapper_107_io_in; // @[package.scala 93:22:@15352.4]
  wire  RetimeWrapper_107_io_out; // @[package.scala 93:22:@15352.4]
  wire  _T_316; // @[MemPrimitives.scala 82:210:@12863.4]
  wire  _T_318; // @[MemPrimitives.scala 82:210:@12864.4]
  wire  _T_319; // @[MemPrimitives.scala 82:228:@12865.4]
  wire  _T_320; // @[MemPrimitives.scala 83:102:@12866.4]
  wire [42:0] _T_322; // @[Cat.scala 30:58:@12868.4]
  wire  _T_329; // @[MemPrimitives.scala 82:210:@12876.4]
  wire  _T_330; // @[MemPrimitives.scala 82:228:@12877.4]
  wire  _T_331; // @[MemPrimitives.scala 83:102:@12878.4]
  wire [42:0] _T_333; // @[Cat.scala 30:58:@12880.4]
  wire  _T_340; // @[MemPrimitives.scala 82:210:@12888.4]
  wire  _T_341; // @[MemPrimitives.scala 82:228:@12889.4]
  wire  _T_342; // @[MemPrimitives.scala 83:102:@12890.4]
  wire [42:0] _T_344; // @[Cat.scala 30:58:@12892.4]
  wire  _T_349; // @[MemPrimitives.scala 82:210:@12899.4]
  wire  _T_352; // @[MemPrimitives.scala 82:228:@12901.4]
  wire  _T_353; // @[MemPrimitives.scala 83:102:@12902.4]
  wire [42:0] _T_355; // @[Cat.scala 30:58:@12904.4]
  wire  _T_363; // @[MemPrimitives.scala 82:228:@12913.4]
  wire  _T_364; // @[MemPrimitives.scala 83:102:@12914.4]
  wire [42:0] _T_366; // @[Cat.scala 30:58:@12916.4]
  wire  _T_374; // @[MemPrimitives.scala 82:228:@12925.4]
  wire  _T_375; // @[MemPrimitives.scala 83:102:@12926.4]
  wire [42:0] _T_377; // @[Cat.scala 30:58:@12928.4]
  wire  _T_382; // @[MemPrimitives.scala 82:210:@12935.4]
  wire  _T_385; // @[MemPrimitives.scala 82:228:@12937.4]
  wire  _T_386; // @[MemPrimitives.scala 83:102:@12938.4]
  wire [42:0] _T_388; // @[Cat.scala 30:58:@12940.4]
  wire  _T_396; // @[MemPrimitives.scala 82:228:@12949.4]
  wire  _T_397; // @[MemPrimitives.scala 83:102:@12950.4]
  wire [42:0] _T_399; // @[Cat.scala 30:58:@12952.4]
  wire  _T_407; // @[MemPrimitives.scala 82:228:@12961.4]
  wire  _T_408; // @[MemPrimitives.scala 83:102:@12962.4]
  wire [42:0] _T_410; // @[Cat.scala 30:58:@12964.4]
  wire  _T_415; // @[MemPrimitives.scala 82:210:@12971.4]
  wire  _T_418; // @[MemPrimitives.scala 82:228:@12973.4]
  wire  _T_419; // @[MemPrimitives.scala 83:102:@12974.4]
  wire [42:0] _T_421; // @[Cat.scala 30:58:@12976.4]
  wire  _T_429; // @[MemPrimitives.scala 82:228:@12985.4]
  wire  _T_430; // @[MemPrimitives.scala 83:102:@12986.4]
  wire [42:0] _T_432; // @[Cat.scala 30:58:@12988.4]
  wire  _T_440; // @[MemPrimitives.scala 82:228:@12997.4]
  wire  _T_441; // @[MemPrimitives.scala 83:102:@12998.4]
  wire [42:0] _T_443; // @[Cat.scala 30:58:@13000.4]
  wire  _T_448; // @[MemPrimitives.scala 110:210:@13007.4]
  wire  _T_450; // @[MemPrimitives.scala 110:210:@13008.4]
  wire  _T_451; // @[MemPrimitives.scala 110:228:@13009.4]
  wire  _T_454; // @[MemPrimitives.scala 110:210:@13011.4]
  wire  _T_456; // @[MemPrimitives.scala 110:210:@13012.4]
  wire  _T_457; // @[MemPrimitives.scala 110:228:@13013.4]
  wire  _T_460; // @[MemPrimitives.scala 110:210:@13015.4]
  wire  _T_462; // @[MemPrimitives.scala 110:210:@13016.4]
  wire  _T_463; // @[MemPrimitives.scala 110:228:@13017.4]
  wire  _T_466; // @[MemPrimitives.scala 110:210:@13019.4]
  wire  _T_468; // @[MemPrimitives.scala 110:210:@13020.4]
  wire  _T_469; // @[MemPrimitives.scala 110:228:@13021.4]
  wire  _T_472; // @[MemPrimitives.scala 110:210:@13023.4]
  wire  _T_474; // @[MemPrimitives.scala 110:210:@13024.4]
  wire  _T_475; // @[MemPrimitives.scala 110:228:@13025.4]
  wire  _T_478; // @[MemPrimitives.scala 110:210:@13027.4]
  wire  _T_480; // @[MemPrimitives.scala 110:210:@13028.4]
  wire  _T_481; // @[MemPrimitives.scala 110:228:@13029.4]
  wire  _T_484; // @[MemPrimitives.scala 110:210:@13031.4]
  wire  _T_486; // @[MemPrimitives.scala 110:210:@13032.4]
  wire  _T_487; // @[MemPrimitives.scala 110:228:@13033.4]
  wire  _T_490; // @[MemPrimitives.scala 110:210:@13035.4]
  wire  _T_492; // @[MemPrimitives.scala 110:210:@13036.4]
  wire  _T_493; // @[MemPrimitives.scala 110:228:@13037.4]
  wire  _T_496; // @[MemPrimitives.scala 110:210:@13039.4]
  wire  _T_498; // @[MemPrimitives.scala 110:210:@13040.4]
  wire  _T_499; // @[MemPrimitives.scala 110:228:@13041.4]
  wire  _T_501; // @[MemPrimitives.scala 126:35:@13055.4]
  wire  _T_502; // @[MemPrimitives.scala 126:35:@13056.4]
  wire  _T_503; // @[MemPrimitives.scala 126:35:@13057.4]
  wire  _T_504; // @[MemPrimitives.scala 126:35:@13058.4]
  wire  _T_505; // @[MemPrimitives.scala 126:35:@13059.4]
  wire  _T_506; // @[MemPrimitives.scala 126:35:@13060.4]
  wire  _T_507; // @[MemPrimitives.scala 126:35:@13061.4]
  wire  _T_508; // @[MemPrimitives.scala 126:35:@13062.4]
  wire  _T_509; // @[MemPrimitives.scala 126:35:@13063.4]
  wire [11:0] _T_511; // @[Cat.scala 30:58:@13065.4]
  wire [11:0] _T_513; // @[Cat.scala 30:58:@13067.4]
  wire [11:0] _T_515; // @[Cat.scala 30:58:@13069.4]
  wire [11:0] _T_517; // @[Cat.scala 30:58:@13071.4]
  wire [11:0] _T_519; // @[Cat.scala 30:58:@13073.4]
  wire [11:0] _T_521; // @[Cat.scala 30:58:@13075.4]
  wire [11:0] _T_523; // @[Cat.scala 30:58:@13077.4]
  wire [11:0] _T_525; // @[Cat.scala 30:58:@13079.4]
  wire [11:0] _T_527; // @[Cat.scala 30:58:@13081.4]
  wire [11:0] _T_528; // @[Mux.scala 31:69:@13082.4]
  wire [11:0] _T_529; // @[Mux.scala 31:69:@13083.4]
  wire [11:0] _T_530; // @[Mux.scala 31:69:@13084.4]
  wire [11:0] _T_531; // @[Mux.scala 31:69:@13085.4]
  wire [11:0] _T_532; // @[Mux.scala 31:69:@13086.4]
  wire [11:0] _T_533; // @[Mux.scala 31:69:@13087.4]
  wire [11:0] _T_534; // @[Mux.scala 31:69:@13088.4]
  wire [11:0] _T_535; // @[Mux.scala 31:69:@13089.4]
  wire  _T_542; // @[MemPrimitives.scala 110:210:@13097.4]
  wire  _T_543; // @[MemPrimitives.scala 110:228:@13098.4]
  wire  _T_548; // @[MemPrimitives.scala 110:210:@13101.4]
  wire  _T_549; // @[MemPrimitives.scala 110:228:@13102.4]
  wire  _T_554; // @[MemPrimitives.scala 110:210:@13105.4]
  wire  _T_555; // @[MemPrimitives.scala 110:228:@13106.4]
  wire  _T_560; // @[MemPrimitives.scala 110:210:@13109.4]
  wire  _T_561; // @[MemPrimitives.scala 110:228:@13110.4]
  wire  _T_566; // @[MemPrimitives.scala 110:210:@13113.4]
  wire  _T_567; // @[MemPrimitives.scala 110:228:@13114.4]
  wire  _T_572; // @[MemPrimitives.scala 110:210:@13117.4]
  wire  _T_573; // @[MemPrimitives.scala 110:228:@13118.4]
  wire  _T_578; // @[MemPrimitives.scala 110:210:@13121.4]
  wire  _T_579; // @[MemPrimitives.scala 110:228:@13122.4]
  wire  _T_584; // @[MemPrimitives.scala 110:210:@13125.4]
  wire  _T_585; // @[MemPrimitives.scala 110:228:@13126.4]
  wire  _T_590; // @[MemPrimitives.scala 110:210:@13129.4]
  wire  _T_591; // @[MemPrimitives.scala 110:228:@13130.4]
  wire  _T_593; // @[MemPrimitives.scala 126:35:@13144.4]
  wire  _T_594; // @[MemPrimitives.scala 126:35:@13145.4]
  wire  _T_595; // @[MemPrimitives.scala 126:35:@13146.4]
  wire  _T_596; // @[MemPrimitives.scala 126:35:@13147.4]
  wire  _T_597; // @[MemPrimitives.scala 126:35:@13148.4]
  wire  _T_598; // @[MemPrimitives.scala 126:35:@13149.4]
  wire  _T_599; // @[MemPrimitives.scala 126:35:@13150.4]
  wire  _T_600; // @[MemPrimitives.scala 126:35:@13151.4]
  wire  _T_601; // @[MemPrimitives.scala 126:35:@13152.4]
  wire [11:0] _T_603; // @[Cat.scala 30:58:@13154.4]
  wire [11:0] _T_605; // @[Cat.scala 30:58:@13156.4]
  wire [11:0] _T_607; // @[Cat.scala 30:58:@13158.4]
  wire [11:0] _T_609; // @[Cat.scala 30:58:@13160.4]
  wire [11:0] _T_611; // @[Cat.scala 30:58:@13162.4]
  wire [11:0] _T_613; // @[Cat.scala 30:58:@13164.4]
  wire [11:0] _T_615; // @[Cat.scala 30:58:@13166.4]
  wire [11:0] _T_617; // @[Cat.scala 30:58:@13168.4]
  wire [11:0] _T_619; // @[Cat.scala 30:58:@13170.4]
  wire [11:0] _T_620; // @[Mux.scala 31:69:@13171.4]
  wire [11:0] _T_621; // @[Mux.scala 31:69:@13172.4]
  wire [11:0] _T_622; // @[Mux.scala 31:69:@13173.4]
  wire [11:0] _T_623; // @[Mux.scala 31:69:@13174.4]
  wire [11:0] _T_624; // @[Mux.scala 31:69:@13175.4]
  wire [11:0] _T_625; // @[Mux.scala 31:69:@13176.4]
  wire [11:0] _T_626; // @[Mux.scala 31:69:@13177.4]
  wire [11:0] _T_627; // @[Mux.scala 31:69:@13178.4]
  wire  _T_634; // @[MemPrimitives.scala 110:210:@13186.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@13187.4]
  wire  _T_640; // @[MemPrimitives.scala 110:210:@13190.4]
  wire  _T_641; // @[MemPrimitives.scala 110:228:@13191.4]
  wire  _T_646; // @[MemPrimitives.scala 110:210:@13194.4]
  wire  _T_647; // @[MemPrimitives.scala 110:228:@13195.4]
  wire  _T_652; // @[MemPrimitives.scala 110:210:@13198.4]
  wire  _T_653; // @[MemPrimitives.scala 110:228:@13199.4]
  wire  _T_658; // @[MemPrimitives.scala 110:210:@13202.4]
  wire  _T_659; // @[MemPrimitives.scala 110:228:@13203.4]
  wire  _T_664; // @[MemPrimitives.scala 110:210:@13206.4]
  wire  _T_665; // @[MemPrimitives.scala 110:228:@13207.4]
  wire  _T_670; // @[MemPrimitives.scala 110:210:@13210.4]
  wire  _T_671; // @[MemPrimitives.scala 110:228:@13211.4]
  wire  _T_676; // @[MemPrimitives.scala 110:210:@13214.4]
  wire  _T_677; // @[MemPrimitives.scala 110:228:@13215.4]
  wire  _T_682; // @[MemPrimitives.scala 110:210:@13218.4]
  wire  _T_683; // @[MemPrimitives.scala 110:228:@13219.4]
  wire  _T_685; // @[MemPrimitives.scala 126:35:@13233.4]
  wire  _T_686; // @[MemPrimitives.scala 126:35:@13234.4]
  wire  _T_687; // @[MemPrimitives.scala 126:35:@13235.4]
  wire  _T_688; // @[MemPrimitives.scala 126:35:@13236.4]
  wire  _T_689; // @[MemPrimitives.scala 126:35:@13237.4]
  wire  _T_690; // @[MemPrimitives.scala 126:35:@13238.4]
  wire  _T_691; // @[MemPrimitives.scala 126:35:@13239.4]
  wire  _T_692; // @[MemPrimitives.scala 126:35:@13240.4]
  wire  _T_693; // @[MemPrimitives.scala 126:35:@13241.4]
  wire [11:0] _T_695; // @[Cat.scala 30:58:@13243.4]
  wire [11:0] _T_697; // @[Cat.scala 30:58:@13245.4]
  wire [11:0] _T_699; // @[Cat.scala 30:58:@13247.4]
  wire [11:0] _T_701; // @[Cat.scala 30:58:@13249.4]
  wire [11:0] _T_703; // @[Cat.scala 30:58:@13251.4]
  wire [11:0] _T_705; // @[Cat.scala 30:58:@13253.4]
  wire [11:0] _T_707; // @[Cat.scala 30:58:@13255.4]
  wire [11:0] _T_709; // @[Cat.scala 30:58:@13257.4]
  wire [11:0] _T_711; // @[Cat.scala 30:58:@13259.4]
  wire [11:0] _T_712; // @[Mux.scala 31:69:@13260.4]
  wire [11:0] _T_713; // @[Mux.scala 31:69:@13261.4]
  wire [11:0] _T_714; // @[Mux.scala 31:69:@13262.4]
  wire [11:0] _T_715; // @[Mux.scala 31:69:@13263.4]
  wire [11:0] _T_716; // @[Mux.scala 31:69:@13264.4]
  wire [11:0] _T_717; // @[Mux.scala 31:69:@13265.4]
  wire [11:0] _T_718; // @[Mux.scala 31:69:@13266.4]
  wire [11:0] _T_719; // @[Mux.scala 31:69:@13267.4]
  wire  _T_724; // @[MemPrimitives.scala 110:210:@13274.4]
  wire  _T_727; // @[MemPrimitives.scala 110:228:@13276.4]
  wire  _T_730; // @[MemPrimitives.scala 110:210:@13278.4]
  wire  _T_733; // @[MemPrimitives.scala 110:228:@13280.4]
  wire  _T_736; // @[MemPrimitives.scala 110:210:@13282.4]
  wire  _T_739; // @[MemPrimitives.scala 110:228:@13284.4]
  wire  _T_742; // @[MemPrimitives.scala 110:210:@13286.4]
  wire  _T_745; // @[MemPrimitives.scala 110:228:@13288.4]
  wire  _T_748; // @[MemPrimitives.scala 110:210:@13290.4]
  wire  _T_751; // @[MemPrimitives.scala 110:228:@13292.4]
  wire  _T_754; // @[MemPrimitives.scala 110:210:@13294.4]
  wire  _T_757; // @[MemPrimitives.scala 110:228:@13296.4]
  wire  _T_760; // @[MemPrimitives.scala 110:210:@13298.4]
  wire  _T_763; // @[MemPrimitives.scala 110:228:@13300.4]
  wire  _T_766; // @[MemPrimitives.scala 110:210:@13302.4]
  wire  _T_769; // @[MemPrimitives.scala 110:228:@13304.4]
  wire  _T_772; // @[MemPrimitives.scala 110:210:@13306.4]
  wire  _T_775; // @[MemPrimitives.scala 110:228:@13308.4]
  wire  _T_777; // @[MemPrimitives.scala 126:35:@13322.4]
  wire  _T_778; // @[MemPrimitives.scala 126:35:@13323.4]
  wire  _T_779; // @[MemPrimitives.scala 126:35:@13324.4]
  wire  _T_780; // @[MemPrimitives.scala 126:35:@13325.4]
  wire  _T_781; // @[MemPrimitives.scala 126:35:@13326.4]
  wire  _T_782; // @[MemPrimitives.scala 126:35:@13327.4]
  wire  _T_783; // @[MemPrimitives.scala 126:35:@13328.4]
  wire  _T_784; // @[MemPrimitives.scala 126:35:@13329.4]
  wire  _T_785; // @[MemPrimitives.scala 126:35:@13330.4]
  wire [11:0] _T_787; // @[Cat.scala 30:58:@13332.4]
  wire [11:0] _T_789; // @[Cat.scala 30:58:@13334.4]
  wire [11:0] _T_791; // @[Cat.scala 30:58:@13336.4]
  wire [11:0] _T_793; // @[Cat.scala 30:58:@13338.4]
  wire [11:0] _T_795; // @[Cat.scala 30:58:@13340.4]
  wire [11:0] _T_797; // @[Cat.scala 30:58:@13342.4]
  wire [11:0] _T_799; // @[Cat.scala 30:58:@13344.4]
  wire [11:0] _T_801; // @[Cat.scala 30:58:@13346.4]
  wire [11:0] _T_803; // @[Cat.scala 30:58:@13348.4]
  wire [11:0] _T_804; // @[Mux.scala 31:69:@13349.4]
  wire [11:0] _T_805; // @[Mux.scala 31:69:@13350.4]
  wire [11:0] _T_806; // @[Mux.scala 31:69:@13351.4]
  wire [11:0] _T_807; // @[Mux.scala 31:69:@13352.4]
  wire [11:0] _T_808; // @[Mux.scala 31:69:@13353.4]
  wire [11:0] _T_809; // @[Mux.scala 31:69:@13354.4]
  wire [11:0] _T_810; // @[Mux.scala 31:69:@13355.4]
  wire [11:0] _T_811; // @[Mux.scala 31:69:@13356.4]
  wire  _T_819; // @[MemPrimitives.scala 110:228:@13365.4]
  wire  _T_825; // @[MemPrimitives.scala 110:228:@13369.4]
  wire  _T_831; // @[MemPrimitives.scala 110:228:@13373.4]
  wire  _T_837; // @[MemPrimitives.scala 110:228:@13377.4]
  wire  _T_843; // @[MemPrimitives.scala 110:228:@13381.4]
  wire  _T_849; // @[MemPrimitives.scala 110:228:@13385.4]
  wire  _T_855; // @[MemPrimitives.scala 110:228:@13389.4]
  wire  _T_861; // @[MemPrimitives.scala 110:228:@13393.4]
  wire  _T_867; // @[MemPrimitives.scala 110:228:@13397.4]
  wire  _T_869; // @[MemPrimitives.scala 126:35:@13411.4]
  wire  _T_870; // @[MemPrimitives.scala 126:35:@13412.4]
  wire  _T_871; // @[MemPrimitives.scala 126:35:@13413.4]
  wire  _T_872; // @[MemPrimitives.scala 126:35:@13414.4]
  wire  _T_873; // @[MemPrimitives.scala 126:35:@13415.4]
  wire  _T_874; // @[MemPrimitives.scala 126:35:@13416.4]
  wire  _T_875; // @[MemPrimitives.scala 126:35:@13417.4]
  wire  _T_876; // @[MemPrimitives.scala 126:35:@13418.4]
  wire  _T_877; // @[MemPrimitives.scala 126:35:@13419.4]
  wire [11:0] _T_879; // @[Cat.scala 30:58:@13421.4]
  wire [11:0] _T_881; // @[Cat.scala 30:58:@13423.4]
  wire [11:0] _T_883; // @[Cat.scala 30:58:@13425.4]
  wire [11:0] _T_885; // @[Cat.scala 30:58:@13427.4]
  wire [11:0] _T_887; // @[Cat.scala 30:58:@13429.4]
  wire [11:0] _T_889; // @[Cat.scala 30:58:@13431.4]
  wire [11:0] _T_891; // @[Cat.scala 30:58:@13433.4]
  wire [11:0] _T_893; // @[Cat.scala 30:58:@13435.4]
  wire [11:0] _T_895; // @[Cat.scala 30:58:@13437.4]
  wire [11:0] _T_896; // @[Mux.scala 31:69:@13438.4]
  wire [11:0] _T_897; // @[Mux.scala 31:69:@13439.4]
  wire [11:0] _T_898; // @[Mux.scala 31:69:@13440.4]
  wire [11:0] _T_899; // @[Mux.scala 31:69:@13441.4]
  wire [11:0] _T_900; // @[Mux.scala 31:69:@13442.4]
  wire [11:0] _T_901; // @[Mux.scala 31:69:@13443.4]
  wire [11:0] _T_902; // @[Mux.scala 31:69:@13444.4]
  wire [11:0] _T_903; // @[Mux.scala 31:69:@13445.4]
  wire  _T_911; // @[MemPrimitives.scala 110:228:@13454.4]
  wire  _T_917; // @[MemPrimitives.scala 110:228:@13458.4]
  wire  _T_923; // @[MemPrimitives.scala 110:228:@13462.4]
  wire  _T_929; // @[MemPrimitives.scala 110:228:@13466.4]
  wire  _T_935; // @[MemPrimitives.scala 110:228:@13470.4]
  wire  _T_941; // @[MemPrimitives.scala 110:228:@13474.4]
  wire  _T_947; // @[MemPrimitives.scala 110:228:@13478.4]
  wire  _T_953; // @[MemPrimitives.scala 110:228:@13482.4]
  wire  _T_959; // @[MemPrimitives.scala 110:228:@13486.4]
  wire  _T_961; // @[MemPrimitives.scala 126:35:@13500.4]
  wire  _T_962; // @[MemPrimitives.scala 126:35:@13501.4]
  wire  _T_963; // @[MemPrimitives.scala 126:35:@13502.4]
  wire  _T_964; // @[MemPrimitives.scala 126:35:@13503.4]
  wire  _T_965; // @[MemPrimitives.scala 126:35:@13504.4]
  wire  _T_966; // @[MemPrimitives.scala 126:35:@13505.4]
  wire  _T_967; // @[MemPrimitives.scala 126:35:@13506.4]
  wire  _T_968; // @[MemPrimitives.scala 126:35:@13507.4]
  wire  _T_969; // @[MemPrimitives.scala 126:35:@13508.4]
  wire [11:0] _T_971; // @[Cat.scala 30:58:@13510.4]
  wire [11:0] _T_973; // @[Cat.scala 30:58:@13512.4]
  wire [11:0] _T_975; // @[Cat.scala 30:58:@13514.4]
  wire [11:0] _T_977; // @[Cat.scala 30:58:@13516.4]
  wire [11:0] _T_979; // @[Cat.scala 30:58:@13518.4]
  wire [11:0] _T_981; // @[Cat.scala 30:58:@13520.4]
  wire [11:0] _T_983; // @[Cat.scala 30:58:@13522.4]
  wire [11:0] _T_985; // @[Cat.scala 30:58:@13524.4]
  wire [11:0] _T_987; // @[Cat.scala 30:58:@13526.4]
  wire [11:0] _T_988; // @[Mux.scala 31:69:@13527.4]
  wire [11:0] _T_989; // @[Mux.scala 31:69:@13528.4]
  wire [11:0] _T_990; // @[Mux.scala 31:69:@13529.4]
  wire [11:0] _T_991; // @[Mux.scala 31:69:@13530.4]
  wire [11:0] _T_992; // @[Mux.scala 31:69:@13531.4]
  wire [11:0] _T_993; // @[Mux.scala 31:69:@13532.4]
  wire [11:0] _T_994; // @[Mux.scala 31:69:@13533.4]
  wire [11:0] _T_995; // @[Mux.scala 31:69:@13534.4]
  wire  _T_1000; // @[MemPrimitives.scala 110:210:@13541.4]
  wire  _T_1003; // @[MemPrimitives.scala 110:228:@13543.4]
  wire  _T_1006; // @[MemPrimitives.scala 110:210:@13545.4]
  wire  _T_1009; // @[MemPrimitives.scala 110:228:@13547.4]
  wire  _T_1012; // @[MemPrimitives.scala 110:210:@13549.4]
  wire  _T_1015; // @[MemPrimitives.scala 110:228:@13551.4]
  wire  _T_1018; // @[MemPrimitives.scala 110:210:@13553.4]
  wire  _T_1021; // @[MemPrimitives.scala 110:228:@13555.4]
  wire  _T_1024; // @[MemPrimitives.scala 110:210:@13557.4]
  wire  _T_1027; // @[MemPrimitives.scala 110:228:@13559.4]
  wire  _T_1030; // @[MemPrimitives.scala 110:210:@13561.4]
  wire  _T_1033; // @[MemPrimitives.scala 110:228:@13563.4]
  wire  _T_1036; // @[MemPrimitives.scala 110:210:@13565.4]
  wire  _T_1039; // @[MemPrimitives.scala 110:228:@13567.4]
  wire  _T_1042; // @[MemPrimitives.scala 110:210:@13569.4]
  wire  _T_1045; // @[MemPrimitives.scala 110:228:@13571.4]
  wire  _T_1048; // @[MemPrimitives.scala 110:210:@13573.4]
  wire  _T_1051; // @[MemPrimitives.scala 110:228:@13575.4]
  wire  _T_1053; // @[MemPrimitives.scala 126:35:@13589.4]
  wire  _T_1054; // @[MemPrimitives.scala 126:35:@13590.4]
  wire  _T_1055; // @[MemPrimitives.scala 126:35:@13591.4]
  wire  _T_1056; // @[MemPrimitives.scala 126:35:@13592.4]
  wire  _T_1057; // @[MemPrimitives.scala 126:35:@13593.4]
  wire  _T_1058; // @[MemPrimitives.scala 126:35:@13594.4]
  wire  _T_1059; // @[MemPrimitives.scala 126:35:@13595.4]
  wire  _T_1060; // @[MemPrimitives.scala 126:35:@13596.4]
  wire  _T_1061; // @[MemPrimitives.scala 126:35:@13597.4]
  wire [11:0] _T_1063; // @[Cat.scala 30:58:@13599.4]
  wire [11:0] _T_1065; // @[Cat.scala 30:58:@13601.4]
  wire [11:0] _T_1067; // @[Cat.scala 30:58:@13603.4]
  wire [11:0] _T_1069; // @[Cat.scala 30:58:@13605.4]
  wire [11:0] _T_1071; // @[Cat.scala 30:58:@13607.4]
  wire [11:0] _T_1073; // @[Cat.scala 30:58:@13609.4]
  wire [11:0] _T_1075; // @[Cat.scala 30:58:@13611.4]
  wire [11:0] _T_1077; // @[Cat.scala 30:58:@13613.4]
  wire [11:0] _T_1079; // @[Cat.scala 30:58:@13615.4]
  wire [11:0] _T_1080; // @[Mux.scala 31:69:@13616.4]
  wire [11:0] _T_1081; // @[Mux.scala 31:69:@13617.4]
  wire [11:0] _T_1082; // @[Mux.scala 31:69:@13618.4]
  wire [11:0] _T_1083; // @[Mux.scala 31:69:@13619.4]
  wire [11:0] _T_1084; // @[Mux.scala 31:69:@13620.4]
  wire [11:0] _T_1085; // @[Mux.scala 31:69:@13621.4]
  wire [11:0] _T_1086; // @[Mux.scala 31:69:@13622.4]
  wire [11:0] _T_1087; // @[Mux.scala 31:69:@13623.4]
  wire  _T_1095; // @[MemPrimitives.scala 110:228:@13632.4]
  wire  _T_1101; // @[MemPrimitives.scala 110:228:@13636.4]
  wire  _T_1107; // @[MemPrimitives.scala 110:228:@13640.4]
  wire  _T_1113; // @[MemPrimitives.scala 110:228:@13644.4]
  wire  _T_1119; // @[MemPrimitives.scala 110:228:@13648.4]
  wire  _T_1125; // @[MemPrimitives.scala 110:228:@13652.4]
  wire  _T_1131; // @[MemPrimitives.scala 110:228:@13656.4]
  wire  _T_1137; // @[MemPrimitives.scala 110:228:@13660.4]
  wire  _T_1143; // @[MemPrimitives.scala 110:228:@13664.4]
  wire  _T_1145; // @[MemPrimitives.scala 126:35:@13678.4]
  wire  _T_1146; // @[MemPrimitives.scala 126:35:@13679.4]
  wire  _T_1147; // @[MemPrimitives.scala 126:35:@13680.4]
  wire  _T_1148; // @[MemPrimitives.scala 126:35:@13681.4]
  wire  _T_1149; // @[MemPrimitives.scala 126:35:@13682.4]
  wire  _T_1150; // @[MemPrimitives.scala 126:35:@13683.4]
  wire  _T_1151; // @[MemPrimitives.scala 126:35:@13684.4]
  wire  _T_1152; // @[MemPrimitives.scala 126:35:@13685.4]
  wire  _T_1153; // @[MemPrimitives.scala 126:35:@13686.4]
  wire [11:0] _T_1155; // @[Cat.scala 30:58:@13688.4]
  wire [11:0] _T_1157; // @[Cat.scala 30:58:@13690.4]
  wire [11:0] _T_1159; // @[Cat.scala 30:58:@13692.4]
  wire [11:0] _T_1161; // @[Cat.scala 30:58:@13694.4]
  wire [11:0] _T_1163; // @[Cat.scala 30:58:@13696.4]
  wire [11:0] _T_1165; // @[Cat.scala 30:58:@13698.4]
  wire [11:0] _T_1167; // @[Cat.scala 30:58:@13700.4]
  wire [11:0] _T_1169; // @[Cat.scala 30:58:@13702.4]
  wire [11:0] _T_1171; // @[Cat.scala 30:58:@13704.4]
  wire [11:0] _T_1172; // @[Mux.scala 31:69:@13705.4]
  wire [11:0] _T_1173; // @[Mux.scala 31:69:@13706.4]
  wire [11:0] _T_1174; // @[Mux.scala 31:69:@13707.4]
  wire [11:0] _T_1175; // @[Mux.scala 31:69:@13708.4]
  wire [11:0] _T_1176; // @[Mux.scala 31:69:@13709.4]
  wire [11:0] _T_1177; // @[Mux.scala 31:69:@13710.4]
  wire [11:0] _T_1178; // @[Mux.scala 31:69:@13711.4]
  wire [11:0] _T_1179; // @[Mux.scala 31:69:@13712.4]
  wire  _T_1187; // @[MemPrimitives.scala 110:228:@13721.4]
  wire  _T_1193; // @[MemPrimitives.scala 110:228:@13725.4]
  wire  _T_1199; // @[MemPrimitives.scala 110:228:@13729.4]
  wire  _T_1205; // @[MemPrimitives.scala 110:228:@13733.4]
  wire  _T_1211; // @[MemPrimitives.scala 110:228:@13737.4]
  wire  _T_1217; // @[MemPrimitives.scala 110:228:@13741.4]
  wire  _T_1223; // @[MemPrimitives.scala 110:228:@13745.4]
  wire  _T_1229; // @[MemPrimitives.scala 110:228:@13749.4]
  wire  _T_1235; // @[MemPrimitives.scala 110:228:@13753.4]
  wire  _T_1237; // @[MemPrimitives.scala 126:35:@13767.4]
  wire  _T_1238; // @[MemPrimitives.scala 126:35:@13768.4]
  wire  _T_1239; // @[MemPrimitives.scala 126:35:@13769.4]
  wire  _T_1240; // @[MemPrimitives.scala 126:35:@13770.4]
  wire  _T_1241; // @[MemPrimitives.scala 126:35:@13771.4]
  wire  _T_1242; // @[MemPrimitives.scala 126:35:@13772.4]
  wire  _T_1243; // @[MemPrimitives.scala 126:35:@13773.4]
  wire  _T_1244; // @[MemPrimitives.scala 126:35:@13774.4]
  wire  _T_1245; // @[MemPrimitives.scala 126:35:@13775.4]
  wire [11:0] _T_1247; // @[Cat.scala 30:58:@13777.4]
  wire [11:0] _T_1249; // @[Cat.scala 30:58:@13779.4]
  wire [11:0] _T_1251; // @[Cat.scala 30:58:@13781.4]
  wire [11:0] _T_1253; // @[Cat.scala 30:58:@13783.4]
  wire [11:0] _T_1255; // @[Cat.scala 30:58:@13785.4]
  wire [11:0] _T_1257; // @[Cat.scala 30:58:@13787.4]
  wire [11:0] _T_1259; // @[Cat.scala 30:58:@13789.4]
  wire [11:0] _T_1261; // @[Cat.scala 30:58:@13791.4]
  wire [11:0] _T_1263; // @[Cat.scala 30:58:@13793.4]
  wire [11:0] _T_1264; // @[Mux.scala 31:69:@13794.4]
  wire [11:0] _T_1265; // @[Mux.scala 31:69:@13795.4]
  wire [11:0] _T_1266; // @[Mux.scala 31:69:@13796.4]
  wire [11:0] _T_1267; // @[Mux.scala 31:69:@13797.4]
  wire [11:0] _T_1268; // @[Mux.scala 31:69:@13798.4]
  wire [11:0] _T_1269; // @[Mux.scala 31:69:@13799.4]
  wire [11:0] _T_1270; // @[Mux.scala 31:69:@13800.4]
  wire [11:0] _T_1271; // @[Mux.scala 31:69:@13801.4]
  wire  _T_1276; // @[MemPrimitives.scala 110:210:@13808.4]
  wire  _T_1279; // @[MemPrimitives.scala 110:228:@13810.4]
  wire  _T_1282; // @[MemPrimitives.scala 110:210:@13812.4]
  wire  _T_1285; // @[MemPrimitives.scala 110:228:@13814.4]
  wire  _T_1288; // @[MemPrimitives.scala 110:210:@13816.4]
  wire  _T_1291; // @[MemPrimitives.scala 110:228:@13818.4]
  wire  _T_1294; // @[MemPrimitives.scala 110:210:@13820.4]
  wire  _T_1297; // @[MemPrimitives.scala 110:228:@13822.4]
  wire  _T_1300; // @[MemPrimitives.scala 110:210:@13824.4]
  wire  _T_1303; // @[MemPrimitives.scala 110:228:@13826.4]
  wire  _T_1306; // @[MemPrimitives.scala 110:210:@13828.4]
  wire  _T_1309; // @[MemPrimitives.scala 110:228:@13830.4]
  wire  _T_1312; // @[MemPrimitives.scala 110:210:@13832.4]
  wire  _T_1315; // @[MemPrimitives.scala 110:228:@13834.4]
  wire  _T_1318; // @[MemPrimitives.scala 110:210:@13836.4]
  wire  _T_1321; // @[MemPrimitives.scala 110:228:@13838.4]
  wire  _T_1324; // @[MemPrimitives.scala 110:210:@13840.4]
  wire  _T_1327; // @[MemPrimitives.scala 110:228:@13842.4]
  wire  _T_1329; // @[MemPrimitives.scala 126:35:@13856.4]
  wire  _T_1330; // @[MemPrimitives.scala 126:35:@13857.4]
  wire  _T_1331; // @[MemPrimitives.scala 126:35:@13858.4]
  wire  _T_1332; // @[MemPrimitives.scala 126:35:@13859.4]
  wire  _T_1333; // @[MemPrimitives.scala 126:35:@13860.4]
  wire  _T_1334; // @[MemPrimitives.scala 126:35:@13861.4]
  wire  _T_1335; // @[MemPrimitives.scala 126:35:@13862.4]
  wire  _T_1336; // @[MemPrimitives.scala 126:35:@13863.4]
  wire  _T_1337; // @[MemPrimitives.scala 126:35:@13864.4]
  wire [11:0] _T_1339; // @[Cat.scala 30:58:@13866.4]
  wire [11:0] _T_1341; // @[Cat.scala 30:58:@13868.4]
  wire [11:0] _T_1343; // @[Cat.scala 30:58:@13870.4]
  wire [11:0] _T_1345; // @[Cat.scala 30:58:@13872.4]
  wire [11:0] _T_1347; // @[Cat.scala 30:58:@13874.4]
  wire [11:0] _T_1349; // @[Cat.scala 30:58:@13876.4]
  wire [11:0] _T_1351; // @[Cat.scala 30:58:@13878.4]
  wire [11:0] _T_1353; // @[Cat.scala 30:58:@13880.4]
  wire [11:0] _T_1355; // @[Cat.scala 30:58:@13882.4]
  wire [11:0] _T_1356; // @[Mux.scala 31:69:@13883.4]
  wire [11:0] _T_1357; // @[Mux.scala 31:69:@13884.4]
  wire [11:0] _T_1358; // @[Mux.scala 31:69:@13885.4]
  wire [11:0] _T_1359; // @[Mux.scala 31:69:@13886.4]
  wire [11:0] _T_1360; // @[Mux.scala 31:69:@13887.4]
  wire [11:0] _T_1361; // @[Mux.scala 31:69:@13888.4]
  wire [11:0] _T_1362; // @[Mux.scala 31:69:@13889.4]
  wire [11:0] _T_1363; // @[Mux.scala 31:69:@13890.4]
  wire  _T_1371; // @[MemPrimitives.scala 110:228:@13899.4]
  wire  _T_1377; // @[MemPrimitives.scala 110:228:@13903.4]
  wire  _T_1383; // @[MemPrimitives.scala 110:228:@13907.4]
  wire  _T_1389; // @[MemPrimitives.scala 110:228:@13911.4]
  wire  _T_1395; // @[MemPrimitives.scala 110:228:@13915.4]
  wire  _T_1401; // @[MemPrimitives.scala 110:228:@13919.4]
  wire  _T_1407; // @[MemPrimitives.scala 110:228:@13923.4]
  wire  _T_1413; // @[MemPrimitives.scala 110:228:@13927.4]
  wire  _T_1419; // @[MemPrimitives.scala 110:228:@13931.4]
  wire  _T_1421; // @[MemPrimitives.scala 126:35:@13945.4]
  wire  _T_1422; // @[MemPrimitives.scala 126:35:@13946.4]
  wire  _T_1423; // @[MemPrimitives.scala 126:35:@13947.4]
  wire  _T_1424; // @[MemPrimitives.scala 126:35:@13948.4]
  wire  _T_1425; // @[MemPrimitives.scala 126:35:@13949.4]
  wire  _T_1426; // @[MemPrimitives.scala 126:35:@13950.4]
  wire  _T_1427; // @[MemPrimitives.scala 126:35:@13951.4]
  wire  _T_1428; // @[MemPrimitives.scala 126:35:@13952.4]
  wire  _T_1429; // @[MemPrimitives.scala 126:35:@13953.4]
  wire [11:0] _T_1431; // @[Cat.scala 30:58:@13955.4]
  wire [11:0] _T_1433; // @[Cat.scala 30:58:@13957.4]
  wire [11:0] _T_1435; // @[Cat.scala 30:58:@13959.4]
  wire [11:0] _T_1437; // @[Cat.scala 30:58:@13961.4]
  wire [11:0] _T_1439; // @[Cat.scala 30:58:@13963.4]
  wire [11:0] _T_1441; // @[Cat.scala 30:58:@13965.4]
  wire [11:0] _T_1443; // @[Cat.scala 30:58:@13967.4]
  wire [11:0] _T_1445; // @[Cat.scala 30:58:@13969.4]
  wire [11:0] _T_1447; // @[Cat.scala 30:58:@13971.4]
  wire [11:0] _T_1448; // @[Mux.scala 31:69:@13972.4]
  wire [11:0] _T_1449; // @[Mux.scala 31:69:@13973.4]
  wire [11:0] _T_1450; // @[Mux.scala 31:69:@13974.4]
  wire [11:0] _T_1451; // @[Mux.scala 31:69:@13975.4]
  wire [11:0] _T_1452; // @[Mux.scala 31:69:@13976.4]
  wire [11:0] _T_1453; // @[Mux.scala 31:69:@13977.4]
  wire [11:0] _T_1454; // @[Mux.scala 31:69:@13978.4]
  wire [11:0] _T_1455; // @[Mux.scala 31:69:@13979.4]
  wire  _T_1463; // @[MemPrimitives.scala 110:228:@13988.4]
  wire  _T_1469; // @[MemPrimitives.scala 110:228:@13992.4]
  wire  _T_1475; // @[MemPrimitives.scala 110:228:@13996.4]
  wire  _T_1481; // @[MemPrimitives.scala 110:228:@14000.4]
  wire  _T_1487; // @[MemPrimitives.scala 110:228:@14004.4]
  wire  _T_1493; // @[MemPrimitives.scala 110:228:@14008.4]
  wire  _T_1499; // @[MemPrimitives.scala 110:228:@14012.4]
  wire  _T_1505; // @[MemPrimitives.scala 110:228:@14016.4]
  wire  _T_1511; // @[MemPrimitives.scala 110:228:@14020.4]
  wire  _T_1513; // @[MemPrimitives.scala 126:35:@14034.4]
  wire  _T_1514; // @[MemPrimitives.scala 126:35:@14035.4]
  wire  _T_1515; // @[MemPrimitives.scala 126:35:@14036.4]
  wire  _T_1516; // @[MemPrimitives.scala 126:35:@14037.4]
  wire  _T_1517; // @[MemPrimitives.scala 126:35:@14038.4]
  wire  _T_1518; // @[MemPrimitives.scala 126:35:@14039.4]
  wire  _T_1519; // @[MemPrimitives.scala 126:35:@14040.4]
  wire  _T_1520; // @[MemPrimitives.scala 126:35:@14041.4]
  wire  _T_1521; // @[MemPrimitives.scala 126:35:@14042.4]
  wire [11:0] _T_1523; // @[Cat.scala 30:58:@14044.4]
  wire [11:0] _T_1525; // @[Cat.scala 30:58:@14046.4]
  wire [11:0] _T_1527; // @[Cat.scala 30:58:@14048.4]
  wire [11:0] _T_1529; // @[Cat.scala 30:58:@14050.4]
  wire [11:0] _T_1531; // @[Cat.scala 30:58:@14052.4]
  wire [11:0] _T_1533; // @[Cat.scala 30:58:@14054.4]
  wire [11:0] _T_1535; // @[Cat.scala 30:58:@14056.4]
  wire [11:0] _T_1537; // @[Cat.scala 30:58:@14058.4]
  wire [11:0] _T_1539; // @[Cat.scala 30:58:@14060.4]
  wire [11:0] _T_1540; // @[Mux.scala 31:69:@14061.4]
  wire [11:0] _T_1541; // @[Mux.scala 31:69:@14062.4]
  wire [11:0] _T_1542; // @[Mux.scala 31:69:@14063.4]
  wire [11:0] _T_1543; // @[Mux.scala 31:69:@14064.4]
  wire [11:0] _T_1544; // @[Mux.scala 31:69:@14065.4]
  wire [11:0] _T_1545; // @[Mux.scala 31:69:@14066.4]
  wire [11:0] _T_1546; // @[Mux.scala 31:69:@14067.4]
  wire [11:0] _T_1547; // @[Mux.scala 31:69:@14068.4]
  wire  _T_1643; // @[package.scala 96:25:@14197.4 package.scala 96:25:@14198.4]
  wire [31:0] _T_1647; // @[Mux.scala 31:69:@14207.4]
  wire  _T_1640; // @[package.scala 96:25:@14189.4 package.scala 96:25:@14190.4]
  wire [31:0] _T_1648; // @[Mux.scala 31:69:@14208.4]
  wire  _T_1637; // @[package.scala 96:25:@14181.4 package.scala 96:25:@14182.4]
  wire [31:0] _T_1649; // @[Mux.scala 31:69:@14209.4]
  wire  _T_1634; // @[package.scala 96:25:@14173.4 package.scala 96:25:@14174.4]
  wire [31:0] _T_1650; // @[Mux.scala 31:69:@14210.4]
  wire  _T_1631; // @[package.scala 96:25:@14165.4 package.scala 96:25:@14166.4]
  wire [31:0] _T_1651; // @[Mux.scala 31:69:@14211.4]
  wire  _T_1628; // @[package.scala 96:25:@14157.4 package.scala 96:25:@14158.4]
  wire [31:0] _T_1652; // @[Mux.scala 31:69:@14212.4]
  wire  _T_1625; // @[package.scala 96:25:@14149.4 package.scala 96:25:@14150.4]
  wire [31:0] _T_1653; // @[Mux.scala 31:69:@14213.4]
  wire  _T_1622; // @[package.scala 96:25:@14141.4 package.scala 96:25:@14142.4]
  wire [31:0] _T_1654; // @[Mux.scala 31:69:@14214.4]
  wire  _T_1619; // @[package.scala 96:25:@14133.4 package.scala 96:25:@14134.4]
  wire [31:0] _T_1655; // @[Mux.scala 31:69:@14215.4]
  wire  _T_1616; // @[package.scala 96:25:@14125.4 package.scala 96:25:@14126.4]
  wire [31:0] _T_1656; // @[Mux.scala 31:69:@14216.4]
  wire  _T_1613; // @[package.scala 96:25:@14117.4 package.scala 96:25:@14118.4]
  wire  _T_1750; // @[package.scala 96:25:@14341.4 package.scala 96:25:@14342.4]
  wire [31:0] _T_1754; // @[Mux.scala 31:69:@14351.4]
  wire  _T_1747; // @[package.scala 96:25:@14333.4 package.scala 96:25:@14334.4]
  wire [31:0] _T_1755; // @[Mux.scala 31:69:@14352.4]
  wire  _T_1744; // @[package.scala 96:25:@14325.4 package.scala 96:25:@14326.4]
  wire [31:0] _T_1756; // @[Mux.scala 31:69:@14353.4]
  wire  _T_1741; // @[package.scala 96:25:@14317.4 package.scala 96:25:@14318.4]
  wire [31:0] _T_1757; // @[Mux.scala 31:69:@14354.4]
  wire  _T_1738; // @[package.scala 96:25:@14309.4 package.scala 96:25:@14310.4]
  wire [31:0] _T_1758; // @[Mux.scala 31:69:@14355.4]
  wire  _T_1735; // @[package.scala 96:25:@14301.4 package.scala 96:25:@14302.4]
  wire [31:0] _T_1759; // @[Mux.scala 31:69:@14356.4]
  wire  _T_1732; // @[package.scala 96:25:@14293.4 package.scala 96:25:@14294.4]
  wire [31:0] _T_1760; // @[Mux.scala 31:69:@14357.4]
  wire  _T_1729; // @[package.scala 96:25:@14285.4 package.scala 96:25:@14286.4]
  wire [31:0] _T_1761; // @[Mux.scala 31:69:@14358.4]
  wire  _T_1726; // @[package.scala 96:25:@14277.4 package.scala 96:25:@14278.4]
  wire [31:0] _T_1762; // @[Mux.scala 31:69:@14359.4]
  wire  _T_1723; // @[package.scala 96:25:@14269.4 package.scala 96:25:@14270.4]
  wire [31:0] _T_1763; // @[Mux.scala 31:69:@14360.4]
  wire  _T_1720; // @[package.scala 96:25:@14261.4 package.scala 96:25:@14262.4]
  wire  _T_1857; // @[package.scala 96:25:@14485.4 package.scala 96:25:@14486.4]
  wire [31:0] _T_1861; // @[Mux.scala 31:69:@14495.4]
  wire  _T_1854; // @[package.scala 96:25:@14477.4 package.scala 96:25:@14478.4]
  wire [31:0] _T_1862; // @[Mux.scala 31:69:@14496.4]
  wire  _T_1851; // @[package.scala 96:25:@14469.4 package.scala 96:25:@14470.4]
  wire [31:0] _T_1863; // @[Mux.scala 31:69:@14497.4]
  wire  _T_1848; // @[package.scala 96:25:@14461.4 package.scala 96:25:@14462.4]
  wire [31:0] _T_1864; // @[Mux.scala 31:69:@14498.4]
  wire  _T_1845; // @[package.scala 96:25:@14453.4 package.scala 96:25:@14454.4]
  wire [31:0] _T_1865; // @[Mux.scala 31:69:@14499.4]
  wire  _T_1842; // @[package.scala 96:25:@14445.4 package.scala 96:25:@14446.4]
  wire [31:0] _T_1866; // @[Mux.scala 31:69:@14500.4]
  wire  _T_1839; // @[package.scala 96:25:@14437.4 package.scala 96:25:@14438.4]
  wire [31:0] _T_1867; // @[Mux.scala 31:69:@14501.4]
  wire  _T_1836; // @[package.scala 96:25:@14429.4 package.scala 96:25:@14430.4]
  wire [31:0] _T_1868; // @[Mux.scala 31:69:@14502.4]
  wire  _T_1833; // @[package.scala 96:25:@14421.4 package.scala 96:25:@14422.4]
  wire [31:0] _T_1869; // @[Mux.scala 31:69:@14503.4]
  wire  _T_1830; // @[package.scala 96:25:@14413.4 package.scala 96:25:@14414.4]
  wire [31:0] _T_1870; // @[Mux.scala 31:69:@14504.4]
  wire  _T_1827; // @[package.scala 96:25:@14405.4 package.scala 96:25:@14406.4]
  wire  _T_1964; // @[package.scala 96:25:@14629.4 package.scala 96:25:@14630.4]
  wire [31:0] _T_1968; // @[Mux.scala 31:69:@14639.4]
  wire  _T_1961; // @[package.scala 96:25:@14621.4 package.scala 96:25:@14622.4]
  wire [31:0] _T_1969; // @[Mux.scala 31:69:@14640.4]
  wire  _T_1958; // @[package.scala 96:25:@14613.4 package.scala 96:25:@14614.4]
  wire [31:0] _T_1970; // @[Mux.scala 31:69:@14641.4]
  wire  _T_1955; // @[package.scala 96:25:@14605.4 package.scala 96:25:@14606.4]
  wire [31:0] _T_1971; // @[Mux.scala 31:69:@14642.4]
  wire  _T_1952; // @[package.scala 96:25:@14597.4 package.scala 96:25:@14598.4]
  wire [31:0] _T_1972; // @[Mux.scala 31:69:@14643.4]
  wire  _T_1949; // @[package.scala 96:25:@14589.4 package.scala 96:25:@14590.4]
  wire [31:0] _T_1973; // @[Mux.scala 31:69:@14644.4]
  wire  _T_1946; // @[package.scala 96:25:@14581.4 package.scala 96:25:@14582.4]
  wire [31:0] _T_1974; // @[Mux.scala 31:69:@14645.4]
  wire  _T_1943; // @[package.scala 96:25:@14573.4 package.scala 96:25:@14574.4]
  wire [31:0] _T_1975; // @[Mux.scala 31:69:@14646.4]
  wire  _T_1940; // @[package.scala 96:25:@14565.4 package.scala 96:25:@14566.4]
  wire [31:0] _T_1976; // @[Mux.scala 31:69:@14647.4]
  wire  _T_1937; // @[package.scala 96:25:@14557.4 package.scala 96:25:@14558.4]
  wire [31:0] _T_1977; // @[Mux.scala 31:69:@14648.4]
  wire  _T_1934; // @[package.scala 96:25:@14549.4 package.scala 96:25:@14550.4]
  wire  _T_2071; // @[package.scala 96:25:@14773.4 package.scala 96:25:@14774.4]
  wire [31:0] _T_2075; // @[Mux.scala 31:69:@14783.4]
  wire  _T_2068; // @[package.scala 96:25:@14765.4 package.scala 96:25:@14766.4]
  wire [31:0] _T_2076; // @[Mux.scala 31:69:@14784.4]
  wire  _T_2065; // @[package.scala 96:25:@14757.4 package.scala 96:25:@14758.4]
  wire [31:0] _T_2077; // @[Mux.scala 31:69:@14785.4]
  wire  _T_2062; // @[package.scala 96:25:@14749.4 package.scala 96:25:@14750.4]
  wire [31:0] _T_2078; // @[Mux.scala 31:69:@14786.4]
  wire  _T_2059; // @[package.scala 96:25:@14741.4 package.scala 96:25:@14742.4]
  wire [31:0] _T_2079; // @[Mux.scala 31:69:@14787.4]
  wire  _T_2056; // @[package.scala 96:25:@14733.4 package.scala 96:25:@14734.4]
  wire [31:0] _T_2080; // @[Mux.scala 31:69:@14788.4]
  wire  _T_2053; // @[package.scala 96:25:@14725.4 package.scala 96:25:@14726.4]
  wire [31:0] _T_2081; // @[Mux.scala 31:69:@14789.4]
  wire  _T_2050; // @[package.scala 96:25:@14717.4 package.scala 96:25:@14718.4]
  wire [31:0] _T_2082; // @[Mux.scala 31:69:@14790.4]
  wire  _T_2047; // @[package.scala 96:25:@14709.4 package.scala 96:25:@14710.4]
  wire [31:0] _T_2083; // @[Mux.scala 31:69:@14791.4]
  wire  _T_2044; // @[package.scala 96:25:@14701.4 package.scala 96:25:@14702.4]
  wire [31:0] _T_2084; // @[Mux.scala 31:69:@14792.4]
  wire  _T_2041; // @[package.scala 96:25:@14693.4 package.scala 96:25:@14694.4]
  wire  _T_2178; // @[package.scala 96:25:@14917.4 package.scala 96:25:@14918.4]
  wire [31:0] _T_2182; // @[Mux.scala 31:69:@14927.4]
  wire  _T_2175; // @[package.scala 96:25:@14909.4 package.scala 96:25:@14910.4]
  wire [31:0] _T_2183; // @[Mux.scala 31:69:@14928.4]
  wire  _T_2172; // @[package.scala 96:25:@14901.4 package.scala 96:25:@14902.4]
  wire [31:0] _T_2184; // @[Mux.scala 31:69:@14929.4]
  wire  _T_2169; // @[package.scala 96:25:@14893.4 package.scala 96:25:@14894.4]
  wire [31:0] _T_2185; // @[Mux.scala 31:69:@14930.4]
  wire  _T_2166; // @[package.scala 96:25:@14885.4 package.scala 96:25:@14886.4]
  wire [31:0] _T_2186; // @[Mux.scala 31:69:@14931.4]
  wire  _T_2163; // @[package.scala 96:25:@14877.4 package.scala 96:25:@14878.4]
  wire [31:0] _T_2187; // @[Mux.scala 31:69:@14932.4]
  wire  _T_2160; // @[package.scala 96:25:@14869.4 package.scala 96:25:@14870.4]
  wire [31:0] _T_2188; // @[Mux.scala 31:69:@14933.4]
  wire  _T_2157; // @[package.scala 96:25:@14861.4 package.scala 96:25:@14862.4]
  wire [31:0] _T_2189; // @[Mux.scala 31:69:@14934.4]
  wire  _T_2154; // @[package.scala 96:25:@14853.4 package.scala 96:25:@14854.4]
  wire [31:0] _T_2190; // @[Mux.scala 31:69:@14935.4]
  wire  _T_2151; // @[package.scala 96:25:@14845.4 package.scala 96:25:@14846.4]
  wire [31:0] _T_2191; // @[Mux.scala 31:69:@14936.4]
  wire  _T_2148; // @[package.scala 96:25:@14837.4 package.scala 96:25:@14838.4]
  wire  _T_2285; // @[package.scala 96:25:@15061.4 package.scala 96:25:@15062.4]
  wire [31:0] _T_2289; // @[Mux.scala 31:69:@15071.4]
  wire  _T_2282; // @[package.scala 96:25:@15053.4 package.scala 96:25:@15054.4]
  wire [31:0] _T_2290; // @[Mux.scala 31:69:@15072.4]
  wire  _T_2279; // @[package.scala 96:25:@15045.4 package.scala 96:25:@15046.4]
  wire [31:0] _T_2291; // @[Mux.scala 31:69:@15073.4]
  wire  _T_2276; // @[package.scala 96:25:@15037.4 package.scala 96:25:@15038.4]
  wire [31:0] _T_2292; // @[Mux.scala 31:69:@15074.4]
  wire  _T_2273; // @[package.scala 96:25:@15029.4 package.scala 96:25:@15030.4]
  wire [31:0] _T_2293; // @[Mux.scala 31:69:@15075.4]
  wire  _T_2270; // @[package.scala 96:25:@15021.4 package.scala 96:25:@15022.4]
  wire [31:0] _T_2294; // @[Mux.scala 31:69:@15076.4]
  wire  _T_2267; // @[package.scala 96:25:@15013.4 package.scala 96:25:@15014.4]
  wire [31:0] _T_2295; // @[Mux.scala 31:69:@15077.4]
  wire  _T_2264; // @[package.scala 96:25:@15005.4 package.scala 96:25:@15006.4]
  wire [31:0] _T_2296; // @[Mux.scala 31:69:@15078.4]
  wire  _T_2261; // @[package.scala 96:25:@14997.4 package.scala 96:25:@14998.4]
  wire [31:0] _T_2297; // @[Mux.scala 31:69:@15079.4]
  wire  _T_2258; // @[package.scala 96:25:@14989.4 package.scala 96:25:@14990.4]
  wire [31:0] _T_2298; // @[Mux.scala 31:69:@15080.4]
  wire  _T_2255; // @[package.scala 96:25:@14981.4 package.scala 96:25:@14982.4]
  wire  _T_2392; // @[package.scala 96:25:@15205.4 package.scala 96:25:@15206.4]
  wire [31:0] _T_2396; // @[Mux.scala 31:69:@15215.4]
  wire  _T_2389; // @[package.scala 96:25:@15197.4 package.scala 96:25:@15198.4]
  wire [31:0] _T_2397; // @[Mux.scala 31:69:@15216.4]
  wire  _T_2386; // @[package.scala 96:25:@15189.4 package.scala 96:25:@15190.4]
  wire [31:0] _T_2398; // @[Mux.scala 31:69:@15217.4]
  wire  _T_2383; // @[package.scala 96:25:@15181.4 package.scala 96:25:@15182.4]
  wire [31:0] _T_2399; // @[Mux.scala 31:69:@15218.4]
  wire  _T_2380; // @[package.scala 96:25:@15173.4 package.scala 96:25:@15174.4]
  wire [31:0] _T_2400; // @[Mux.scala 31:69:@15219.4]
  wire  _T_2377; // @[package.scala 96:25:@15165.4 package.scala 96:25:@15166.4]
  wire [31:0] _T_2401; // @[Mux.scala 31:69:@15220.4]
  wire  _T_2374; // @[package.scala 96:25:@15157.4 package.scala 96:25:@15158.4]
  wire [31:0] _T_2402; // @[Mux.scala 31:69:@15221.4]
  wire  _T_2371; // @[package.scala 96:25:@15149.4 package.scala 96:25:@15150.4]
  wire [31:0] _T_2403; // @[Mux.scala 31:69:@15222.4]
  wire  _T_2368; // @[package.scala 96:25:@15141.4 package.scala 96:25:@15142.4]
  wire [31:0] _T_2404; // @[Mux.scala 31:69:@15223.4]
  wire  _T_2365; // @[package.scala 96:25:@15133.4 package.scala 96:25:@15134.4]
  wire [31:0] _T_2405; // @[Mux.scala 31:69:@15224.4]
  wire  _T_2362; // @[package.scala 96:25:@15125.4 package.scala 96:25:@15126.4]
  wire  _T_2499; // @[package.scala 96:25:@15349.4 package.scala 96:25:@15350.4]
  wire [31:0] _T_2503; // @[Mux.scala 31:69:@15359.4]
  wire  _T_2496; // @[package.scala 96:25:@15341.4 package.scala 96:25:@15342.4]
  wire [31:0] _T_2504; // @[Mux.scala 31:69:@15360.4]
  wire  _T_2493; // @[package.scala 96:25:@15333.4 package.scala 96:25:@15334.4]
  wire [31:0] _T_2505; // @[Mux.scala 31:69:@15361.4]
  wire  _T_2490; // @[package.scala 96:25:@15325.4 package.scala 96:25:@15326.4]
  wire [31:0] _T_2506; // @[Mux.scala 31:69:@15362.4]
  wire  _T_2487; // @[package.scala 96:25:@15317.4 package.scala 96:25:@15318.4]
  wire [31:0] _T_2507; // @[Mux.scala 31:69:@15363.4]
  wire  _T_2484; // @[package.scala 96:25:@15309.4 package.scala 96:25:@15310.4]
  wire [31:0] _T_2508; // @[Mux.scala 31:69:@15364.4]
  wire  _T_2481; // @[package.scala 96:25:@15301.4 package.scala 96:25:@15302.4]
  wire [31:0] _T_2509; // @[Mux.scala 31:69:@15365.4]
  wire  _T_2478; // @[package.scala 96:25:@15293.4 package.scala 96:25:@15294.4]
  wire [31:0] _T_2510; // @[Mux.scala 31:69:@15366.4]
  wire  _T_2475; // @[package.scala 96:25:@15285.4 package.scala 96:25:@15286.4]
  wire [31:0] _T_2511; // @[Mux.scala 31:69:@15367.4]
  wire  _T_2472; // @[package.scala 96:25:@15277.4 package.scala 96:25:@15278.4]
  wire [31:0] _T_2512; // @[Mux.scala 31:69:@15368.4]
  wire  _T_2469; // @[package.scala 96:25:@15269.4 package.scala 96:25:@15270.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@12671.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@12687.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@12703.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@12719.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@12735.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@12751.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@12767.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@12783.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@12799.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@12815.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@12831.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@12847.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  StickySelects_1 StickySelects ( // @[MemPrimitives.scala 124:33:@13043.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_ins_6(StickySelects_io_ins_6),
    .io_ins_7(StickySelects_io_ins_7),
    .io_ins_8(StickySelects_io_ins_8),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5),
    .io_outs_6(StickySelects_io_outs_6),
    .io_outs_7(StickySelects_io_outs_7),
    .io_outs_8(StickySelects_io_outs_8)
  );
  StickySelects_1 StickySelects_1 ( // @[MemPrimitives.scala 124:33:@13132.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_ins_6(StickySelects_1_io_ins_6),
    .io_ins_7(StickySelects_1_io_ins_7),
    .io_ins_8(StickySelects_1_io_ins_8),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5),
    .io_outs_6(StickySelects_1_io_outs_6),
    .io_outs_7(StickySelects_1_io_outs_7),
    .io_outs_8(StickySelects_1_io_outs_8)
  );
  StickySelects_1 StickySelects_2 ( // @[MemPrimitives.scala 124:33:@13221.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_ins_6(StickySelects_2_io_ins_6),
    .io_ins_7(StickySelects_2_io_ins_7),
    .io_ins_8(StickySelects_2_io_ins_8),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5),
    .io_outs_6(StickySelects_2_io_outs_6),
    .io_outs_7(StickySelects_2_io_outs_7),
    .io_outs_8(StickySelects_2_io_outs_8)
  );
  StickySelects_1 StickySelects_3 ( // @[MemPrimitives.scala 124:33:@13310.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_ins_6(StickySelects_3_io_ins_6),
    .io_ins_7(StickySelects_3_io_ins_7),
    .io_ins_8(StickySelects_3_io_ins_8),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5),
    .io_outs_6(StickySelects_3_io_outs_6),
    .io_outs_7(StickySelects_3_io_outs_7),
    .io_outs_8(StickySelects_3_io_outs_8)
  );
  StickySelects_1 StickySelects_4 ( // @[MemPrimitives.scala 124:33:@13399.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_ins_6(StickySelects_4_io_ins_6),
    .io_ins_7(StickySelects_4_io_ins_7),
    .io_ins_8(StickySelects_4_io_ins_8),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5),
    .io_outs_6(StickySelects_4_io_outs_6),
    .io_outs_7(StickySelects_4_io_outs_7),
    .io_outs_8(StickySelects_4_io_outs_8)
  );
  StickySelects_1 StickySelects_5 ( // @[MemPrimitives.scala 124:33:@13488.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_ins_6(StickySelects_5_io_ins_6),
    .io_ins_7(StickySelects_5_io_ins_7),
    .io_ins_8(StickySelects_5_io_ins_8),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5),
    .io_outs_6(StickySelects_5_io_outs_6),
    .io_outs_7(StickySelects_5_io_outs_7),
    .io_outs_8(StickySelects_5_io_outs_8)
  );
  StickySelects_1 StickySelects_6 ( // @[MemPrimitives.scala 124:33:@13577.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_ins_6(StickySelects_6_io_ins_6),
    .io_ins_7(StickySelects_6_io_ins_7),
    .io_ins_8(StickySelects_6_io_ins_8),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5),
    .io_outs_6(StickySelects_6_io_outs_6),
    .io_outs_7(StickySelects_6_io_outs_7),
    .io_outs_8(StickySelects_6_io_outs_8)
  );
  StickySelects_1 StickySelects_7 ( // @[MemPrimitives.scala 124:33:@13666.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_ins_6(StickySelects_7_io_ins_6),
    .io_ins_7(StickySelects_7_io_ins_7),
    .io_ins_8(StickySelects_7_io_ins_8),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5),
    .io_outs_6(StickySelects_7_io_outs_6),
    .io_outs_7(StickySelects_7_io_outs_7),
    .io_outs_8(StickySelects_7_io_outs_8)
  );
  StickySelects_1 StickySelects_8 ( // @[MemPrimitives.scala 124:33:@13755.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_ins_6(StickySelects_8_io_ins_6),
    .io_ins_7(StickySelects_8_io_ins_7),
    .io_ins_8(StickySelects_8_io_ins_8),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5),
    .io_outs_6(StickySelects_8_io_outs_6),
    .io_outs_7(StickySelects_8_io_outs_7),
    .io_outs_8(StickySelects_8_io_outs_8)
  );
  StickySelects_1 StickySelects_9 ( // @[MemPrimitives.scala 124:33:@13844.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_ins_6(StickySelects_9_io_ins_6),
    .io_ins_7(StickySelects_9_io_ins_7),
    .io_ins_8(StickySelects_9_io_ins_8),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5),
    .io_outs_6(StickySelects_9_io_outs_6),
    .io_outs_7(StickySelects_9_io_outs_7),
    .io_outs_8(StickySelects_9_io_outs_8)
  );
  StickySelects_1 StickySelects_10 ( // @[MemPrimitives.scala 124:33:@13933.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_ins_6(StickySelects_10_io_ins_6),
    .io_ins_7(StickySelects_10_io_ins_7),
    .io_ins_8(StickySelects_10_io_ins_8),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5),
    .io_outs_6(StickySelects_10_io_outs_6),
    .io_outs_7(StickySelects_10_io_outs_7),
    .io_outs_8(StickySelects_10_io_outs_8)
  );
  StickySelects_1 StickySelects_11 ( // @[MemPrimitives.scala 124:33:@14022.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_ins_6(StickySelects_11_io_ins_6),
    .io_ins_7(StickySelects_11_io_ins_7),
    .io_ins_8(StickySelects_11_io_ins_8),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5),
    .io_outs_6(StickySelects_11_io_outs_6),
    .io_outs_7(StickySelects_11_io_outs_7),
    .io_outs_8(StickySelects_11_io_outs_8)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@14112.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@14120.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@14128.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@14136.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@14144.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@14152.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@14160.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@14168.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@14176.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@14184.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@14192.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@14200.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@14256.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@14264.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@14272.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@14280.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@14288.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@14296.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@14304.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@14312.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@14320.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@14328.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@14336.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@14344.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@14400.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@14408.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@14416.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@14424.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@14432.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@14440.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@14448.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@14456.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@14464.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@14472.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@14480.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@14488.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@14544.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@14552.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@14560.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@14568.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@14576.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@14584.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@14592.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@14600.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@14608.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@14616.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@14624.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@14632.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_48 ( // @[package.scala 93:22:@14688.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@14696.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_50 ( // @[package.scala 93:22:@14704.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@14712.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@14720.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_53 ( // @[package.scala 93:22:@14728.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@14736.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_55 ( // @[package.scala 93:22:@14744.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@14752.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_57 ( // @[package.scala 93:22:@14760.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@14768.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_59 ( // @[package.scala 93:22:@14776.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_60 ( // @[package.scala 93:22:@14832.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_61 ( // @[package.scala 93:22:@14840.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_62 ( // @[package.scala 93:22:@14848.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_63 ( // @[package.scala 93:22:@14856.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_64 ( // @[package.scala 93:22:@14864.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_65 ( // @[package.scala 93:22:@14872.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_66 ( // @[package.scala 93:22:@14880.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_67 ( // @[package.scala 93:22:@14888.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_68 ( // @[package.scala 93:22:@14896.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_69 ( // @[package.scala 93:22:@14904.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_70 ( // @[package.scala 93:22:@14912.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_71 ( // @[package.scala 93:22:@14920.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_72 ( // @[package.scala 93:22:@14976.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_73 ( // @[package.scala 93:22:@14984.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_74 ( // @[package.scala 93:22:@14992.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_75 ( // @[package.scala 93:22:@15000.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_76 ( // @[package.scala 93:22:@15008.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_77 ( // @[package.scala 93:22:@15016.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_78 ( // @[package.scala 93:22:@15024.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_79 ( // @[package.scala 93:22:@15032.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_80 ( // @[package.scala 93:22:@15040.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_81 ( // @[package.scala 93:22:@15048.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_82 ( // @[package.scala 93:22:@15056.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_83 ( // @[package.scala 93:22:@15064.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_84 ( // @[package.scala 93:22:@15120.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_85 ( // @[package.scala 93:22:@15128.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_86 ( // @[package.scala 93:22:@15136.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_87 ( // @[package.scala 93:22:@15144.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_88 ( // @[package.scala 93:22:@15152.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_89 ( // @[package.scala 93:22:@15160.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_90 ( // @[package.scala 93:22:@15168.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_91 ( // @[package.scala 93:22:@15176.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_92 ( // @[package.scala 93:22:@15184.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_93 ( // @[package.scala 93:22:@15192.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_94 ( // @[package.scala 93:22:@15200.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_95 ( // @[package.scala 93:22:@15208.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_96 ( // @[package.scala 93:22:@15264.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_97 ( // @[package.scala 93:22:@15272.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_98 ( // @[package.scala 93:22:@15280.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_99 ( // @[package.scala 93:22:@15288.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_100 ( // @[package.scala 93:22:@15296.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_101 ( // @[package.scala 93:22:@15304.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_102 ( // @[package.scala 93:22:@15312.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_103 ( // @[package.scala 93:22:@15320.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_104 ( // @[package.scala 93:22:@15328.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_105 ( // @[package.scala 93:22:@15336.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_106 ( // @[package.scala 93:22:@15344.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_107 ( // @[package.scala 93:22:@15352.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  assign _T_316 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@12863.4]
  assign _T_318 = io_wPort_0_banks_1 == 2'h0; // @[MemPrimitives.scala 82:210:@12864.4]
  assign _T_319 = _T_316 & _T_318; // @[MemPrimitives.scala 82:228:@12865.4]
  assign _T_320 = io_wPort_0_en_0 & _T_319; // @[MemPrimitives.scala 83:102:@12866.4]
  assign _T_322 = {_T_320,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12868.4]
  assign _T_329 = io_wPort_0_banks_1 == 2'h1; // @[MemPrimitives.scala 82:210:@12876.4]
  assign _T_330 = _T_316 & _T_329; // @[MemPrimitives.scala 82:228:@12877.4]
  assign _T_331 = io_wPort_0_en_0 & _T_330; // @[MemPrimitives.scala 83:102:@12878.4]
  assign _T_333 = {_T_331,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12880.4]
  assign _T_340 = io_wPort_0_banks_1 == 2'h2; // @[MemPrimitives.scala 82:210:@12888.4]
  assign _T_341 = _T_316 & _T_340; // @[MemPrimitives.scala 82:228:@12889.4]
  assign _T_342 = io_wPort_0_en_0 & _T_341; // @[MemPrimitives.scala 83:102:@12890.4]
  assign _T_344 = {_T_342,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12892.4]
  assign _T_349 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@12899.4]
  assign _T_352 = _T_349 & _T_318; // @[MemPrimitives.scala 82:228:@12901.4]
  assign _T_353 = io_wPort_0_en_0 & _T_352; // @[MemPrimitives.scala 83:102:@12902.4]
  assign _T_355 = {_T_353,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12904.4]
  assign _T_363 = _T_349 & _T_329; // @[MemPrimitives.scala 82:228:@12913.4]
  assign _T_364 = io_wPort_0_en_0 & _T_363; // @[MemPrimitives.scala 83:102:@12914.4]
  assign _T_366 = {_T_364,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12916.4]
  assign _T_374 = _T_349 & _T_340; // @[MemPrimitives.scala 82:228:@12925.4]
  assign _T_375 = io_wPort_0_en_0 & _T_374; // @[MemPrimitives.scala 83:102:@12926.4]
  assign _T_377 = {_T_375,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12928.4]
  assign _T_382 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@12935.4]
  assign _T_385 = _T_382 & _T_318; // @[MemPrimitives.scala 82:228:@12937.4]
  assign _T_386 = io_wPort_0_en_0 & _T_385; // @[MemPrimitives.scala 83:102:@12938.4]
  assign _T_388 = {_T_386,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12940.4]
  assign _T_396 = _T_382 & _T_329; // @[MemPrimitives.scala 82:228:@12949.4]
  assign _T_397 = io_wPort_0_en_0 & _T_396; // @[MemPrimitives.scala 83:102:@12950.4]
  assign _T_399 = {_T_397,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12952.4]
  assign _T_407 = _T_382 & _T_340; // @[MemPrimitives.scala 82:228:@12961.4]
  assign _T_408 = io_wPort_0_en_0 & _T_407; // @[MemPrimitives.scala 83:102:@12962.4]
  assign _T_410 = {_T_408,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12964.4]
  assign _T_415 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@12971.4]
  assign _T_418 = _T_415 & _T_318; // @[MemPrimitives.scala 82:228:@12973.4]
  assign _T_419 = io_wPort_0_en_0 & _T_418; // @[MemPrimitives.scala 83:102:@12974.4]
  assign _T_421 = {_T_419,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12976.4]
  assign _T_429 = _T_415 & _T_329; // @[MemPrimitives.scala 82:228:@12985.4]
  assign _T_430 = io_wPort_0_en_0 & _T_429; // @[MemPrimitives.scala 83:102:@12986.4]
  assign _T_432 = {_T_430,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12988.4]
  assign _T_440 = _T_415 & _T_340; // @[MemPrimitives.scala 82:228:@12997.4]
  assign _T_441 = io_wPort_0_en_0 & _T_440; // @[MemPrimitives.scala 83:102:@12998.4]
  assign _T_443 = {_T_441,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13000.4]
  assign _T_448 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13007.4]
  assign _T_450 = io_rPort_0_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13008.4]
  assign _T_451 = _T_448 & _T_450; // @[MemPrimitives.scala 110:228:@13009.4]
  assign _T_454 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13011.4]
  assign _T_456 = io_rPort_1_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13012.4]
  assign _T_457 = _T_454 & _T_456; // @[MemPrimitives.scala 110:228:@13013.4]
  assign _T_460 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13015.4]
  assign _T_462 = io_rPort_2_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13016.4]
  assign _T_463 = _T_460 & _T_462; // @[MemPrimitives.scala 110:228:@13017.4]
  assign _T_466 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13019.4]
  assign _T_468 = io_rPort_3_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13020.4]
  assign _T_469 = _T_466 & _T_468; // @[MemPrimitives.scala 110:228:@13021.4]
  assign _T_472 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13023.4]
  assign _T_474 = io_rPort_4_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13024.4]
  assign _T_475 = _T_472 & _T_474; // @[MemPrimitives.scala 110:228:@13025.4]
  assign _T_478 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13027.4]
  assign _T_480 = io_rPort_5_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13028.4]
  assign _T_481 = _T_478 & _T_480; // @[MemPrimitives.scala 110:228:@13029.4]
  assign _T_484 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13031.4]
  assign _T_486 = io_rPort_6_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13032.4]
  assign _T_487 = _T_484 & _T_486; // @[MemPrimitives.scala 110:228:@13033.4]
  assign _T_490 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13035.4]
  assign _T_492 = io_rPort_7_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13036.4]
  assign _T_493 = _T_490 & _T_492; // @[MemPrimitives.scala 110:228:@13037.4]
  assign _T_496 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13039.4]
  assign _T_498 = io_rPort_8_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13040.4]
  assign _T_499 = _T_496 & _T_498; // @[MemPrimitives.scala 110:228:@13041.4]
  assign _T_501 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@13055.4]
  assign _T_502 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@13056.4]
  assign _T_503 = StickySelects_io_outs_2; // @[MemPrimitives.scala 126:35:@13057.4]
  assign _T_504 = StickySelects_io_outs_3; // @[MemPrimitives.scala 126:35:@13058.4]
  assign _T_505 = StickySelects_io_outs_4; // @[MemPrimitives.scala 126:35:@13059.4]
  assign _T_506 = StickySelects_io_outs_5; // @[MemPrimitives.scala 126:35:@13060.4]
  assign _T_507 = StickySelects_io_outs_6; // @[MemPrimitives.scala 126:35:@13061.4]
  assign _T_508 = StickySelects_io_outs_7; // @[MemPrimitives.scala 126:35:@13062.4]
  assign _T_509 = StickySelects_io_outs_8; // @[MemPrimitives.scala 126:35:@13063.4]
  assign _T_511 = {_T_501,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13065.4]
  assign _T_513 = {_T_502,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13067.4]
  assign _T_515 = {_T_503,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13069.4]
  assign _T_517 = {_T_504,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13071.4]
  assign _T_519 = {_T_505,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13073.4]
  assign _T_521 = {_T_506,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13075.4]
  assign _T_523 = {_T_507,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13077.4]
  assign _T_525 = {_T_508,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13079.4]
  assign _T_527 = {_T_509,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13081.4]
  assign _T_528 = _T_508 ? _T_525 : _T_527; // @[Mux.scala 31:69:@13082.4]
  assign _T_529 = _T_507 ? _T_523 : _T_528; // @[Mux.scala 31:69:@13083.4]
  assign _T_530 = _T_506 ? _T_521 : _T_529; // @[Mux.scala 31:69:@13084.4]
  assign _T_531 = _T_505 ? _T_519 : _T_530; // @[Mux.scala 31:69:@13085.4]
  assign _T_532 = _T_504 ? _T_517 : _T_531; // @[Mux.scala 31:69:@13086.4]
  assign _T_533 = _T_503 ? _T_515 : _T_532; // @[Mux.scala 31:69:@13087.4]
  assign _T_534 = _T_502 ? _T_513 : _T_533; // @[Mux.scala 31:69:@13088.4]
  assign _T_535 = _T_501 ? _T_511 : _T_534; // @[Mux.scala 31:69:@13089.4]
  assign _T_542 = io_rPort_0_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13097.4]
  assign _T_543 = _T_448 & _T_542; // @[MemPrimitives.scala 110:228:@13098.4]
  assign _T_548 = io_rPort_1_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13101.4]
  assign _T_549 = _T_454 & _T_548; // @[MemPrimitives.scala 110:228:@13102.4]
  assign _T_554 = io_rPort_2_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13105.4]
  assign _T_555 = _T_460 & _T_554; // @[MemPrimitives.scala 110:228:@13106.4]
  assign _T_560 = io_rPort_3_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13109.4]
  assign _T_561 = _T_466 & _T_560; // @[MemPrimitives.scala 110:228:@13110.4]
  assign _T_566 = io_rPort_4_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13113.4]
  assign _T_567 = _T_472 & _T_566; // @[MemPrimitives.scala 110:228:@13114.4]
  assign _T_572 = io_rPort_5_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13117.4]
  assign _T_573 = _T_478 & _T_572; // @[MemPrimitives.scala 110:228:@13118.4]
  assign _T_578 = io_rPort_6_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13121.4]
  assign _T_579 = _T_484 & _T_578; // @[MemPrimitives.scala 110:228:@13122.4]
  assign _T_584 = io_rPort_7_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13125.4]
  assign _T_585 = _T_490 & _T_584; // @[MemPrimitives.scala 110:228:@13126.4]
  assign _T_590 = io_rPort_8_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13129.4]
  assign _T_591 = _T_496 & _T_590; // @[MemPrimitives.scala 110:228:@13130.4]
  assign _T_593 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 126:35:@13144.4]
  assign _T_594 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 126:35:@13145.4]
  assign _T_595 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 126:35:@13146.4]
  assign _T_596 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 126:35:@13147.4]
  assign _T_597 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 126:35:@13148.4]
  assign _T_598 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 126:35:@13149.4]
  assign _T_599 = StickySelects_1_io_outs_6; // @[MemPrimitives.scala 126:35:@13150.4]
  assign _T_600 = StickySelects_1_io_outs_7; // @[MemPrimitives.scala 126:35:@13151.4]
  assign _T_601 = StickySelects_1_io_outs_8; // @[MemPrimitives.scala 126:35:@13152.4]
  assign _T_603 = {_T_593,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13154.4]
  assign _T_605 = {_T_594,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13156.4]
  assign _T_607 = {_T_595,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13158.4]
  assign _T_609 = {_T_596,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13160.4]
  assign _T_611 = {_T_597,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13162.4]
  assign _T_613 = {_T_598,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13164.4]
  assign _T_615 = {_T_599,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13166.4]
  assign _T_617 = {_T_600,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13168.4]
  assign _T_619 = {_T_601,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13170.4]
  assign _T_620 = _T_600 ? _T_617 : _T_619; // @[Mux.scala 31:69:@13171.4]
  assign _T_621 = _T_599 ? _T_615 : _T_620; // @[Mux.scala 31:69:@13172.4]
  assign _T_622 = _T_598 ? _T_613 : _T_621; // @[Mux.scala 31:69:@13173.4]
  assign _T_623 = _T_597 ? _T_611 : _T_622; // @[Mux.scala 31:69:@13174.4]
  assign _T_624 = _T_596 ? _T_609 : _T_623; // @[Mux.scala 31:69:@13175.4]
  assign _T_625 = _T_595 ? _T_607 : _T_624; // @[Mux.scala 31:69:@13176.4]
  assign _T_626 = _T_594 ? _T_605 : _T_625; // @[Mux.scala 31:69:@13177.4]
  assign _T_627 = _T_593 ? _T_603 : _T_626; // @[Mux.scala 31:69:@13178.4]
  assign _T_634 = io_rPort_0_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13186.4]
  assign _T_635 = _T_448 & _T_634; // @[MemPrimitives.scala 110:228:@13187.4]
  assign _T_640 = io_rPort_1_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13190.4]
  assign _T_641 = _T_454 & _T_640; // @[MemPrimitives.scala 110:228:@13191.4]
  assign _T_646 = io_rPort_2_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13194.4]
  assign _T_647 = _T_460 & _T_646; // @[MemPrimitives.scala 110:228:@13195.4]
  assign _T_652 = io_rPort_3_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13198.4]
  assign _T_653 = _T_466 & _T_652; // @[MemPrimitives.scala 110:228:@13199.4]
  assign _T_658 = io_rPort_4_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13202.4]
  assign _T_659 = _T_472 & _T_658; // @[MemPrimitives.scala 110:228:@13203.4]
  assign _T_664 = io_rPort_5_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13206.4]
  assign _T_665 = _T_478 & _T_664; // @[MemPrimitives.scala 110:228:@13207.4]
  assign _T_670 = io_rPort_6_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13210.4]
  assign _T_671 = _T_484 & _T_670; // @[MemPrimitives.scala 110:228:@13211.4]
  assign _T_676 = io_rPort_7_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13214.4]
  assign _T_677 = _T_490 & _T_676; // @[MemPrimitives.scala 110:228:@13215.4]
  assign _T_682 = io_rPort_8_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13218.4]
  assign _T_683 = _T_496 & _T_682; // @[MemPrimitives.scala 110:228:@13219.4]
  assign _T_685 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 126:35:@13233.4]
  assign _T_686 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 126:35:@13234.4]
  assign _T_687 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 126:35:@13235.4]
  assign _T_688 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 126:35:@13236.4]
  assign _T_689 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 126:35:@13237.4]
  assign _T_690 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 126:35:@13238.4]
  assign _T_691 = StickySelects_2_io_outs_6; // @[MemPrimitives.scala 126:35:@13239.4]
  assign _T_692 = StickySelects_2_io_outs_7; // @[MemPrimitives.scala 126:35:@13240.4]
  assign _T_693 = StickySelects_2_io_outs_8; // @[MemPrimitives.scala 126:35:@13241.4]
  assign _T_695 = {_T_685,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13243.4]
  assign _T_697 = {_T_686,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13245.4]
  assign _T_699 = {_T_687,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13247.4]
  assign _T_701 = {_T_688,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13249.4]
  assign _T_703 = {_T_689,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13251.4]
  assign _T_705 = {_T_690,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13253.4]
  assign _T_707 = {_T_691,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13255.4]
  assign _T_709 = {_T_692,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13257.4]
  assign _T_711 = {_T_693,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13259.4]
  assign _T_712 = _T_692 ? _T_709 : _T_711; // @[Mux.scala 31:69:@13260.4]
  assign _T_713 = _T_691 ? _T_707 : _T_712; // @[Mux.scala 31:69:@13261.4]
  assign _T_714 = _T_690 ? _T_705 : _T_713; // @[Mux.scala 31:69:@13262.4]
  assign _T_715 = _T_689 ? _T_703 : _T_714; // @[Mux.scala 31:69:@13263.4]
  assign _T_716 = _T_688 ? _T_701 : _T_715; // @[Mux.scala 31:69:@13264.4]
  assign _T_717 = _T_687 ? _T_699 : _T_716; // @[Mux.scala 31:69:@13265.4]
  assign _T_718 = _T_686 ? _T_697 : _T_717; // @[Mux.scala 31:69:@13266.4]
  assign _T_719 = _T_685 ? _T_695 : _T_718; // @[Mux.scala 31:69:@13267.4]
  assign _T_724 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13274.4]
  assign _T_727 = _T_724 & _T_450; // @[MemPrimitives.scala 110:228:@13276.4]
  assign _T_730 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13278.4]
  assign _T_733 = _T_730 & _T_456; // @[MemPrimitives.scala 110:228:@13280.4]
  assign _T_736 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13282.4]
  assign _T_739 = _T_736 & _T_462; // @[MemPrimitives.scala 110:228:@13284.4]
  assign _T_742 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13286.4]
  assign _T_745 = _T_742 & _T_468; // @[MemPrimitives.scala 110:228:@13288.4]
  assign _T_748 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13290.4]
  assign _T_751 = _T_748 & _T_474; // @[MemPrimitives.scala 110:228:@13292.4]
  assign _T_754 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13294.4]
  assign _T_757 = _T_754 & _T_480; // @[MemPrimitives.scala 110:228:@13296.4]
  assign _T_760 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13298.4]
  assign _T_763 = _T_760 & _T_486; // @[MemPrimitives.scala 110:228:@13300.4]
  assign _T_766 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13302.4]
  assign _T_769 = _T_766 & _T_492; // @[MemPrimitives.scala 110:228:@13304.4]
  assign _T_772 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13306.4]
  assign _T_775 = _T_772 & _T_498; // @[MemPrimitives.scala 110:228:@13308.4]
  assign _T_777 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 126:35:@13322.4]
  assign _T_778 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 126:35:@13323.4]
  assign _T_779 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 126:35:@13324.4]
  assign _T_780 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 126:35:@13325.4]
  assign _T_781 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 126:35:@13326.4]
  assign _T_782 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 126:35:@13327.4]
  assign _T_783 = StickySelects_3_io_outs_6; // @[MemPrimitives.scala 126:35:@13328.4]
  assign _T_784 = StickySelects_3_io_outs_7; // @[MemPrimitives.scala 126:35:@13329.4]
  assign _T_785 = StickySelects_3_io_outs_8; // @[MemPrimitives.scala 126:35:@13330.4]
  assign _T_787 = {_T_777,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13332.4]
  assign _T_789 = {_T_778,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13334.4]
  assign _T_791 = {_T_779,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13336.4]
  assign _T_793 = {_T_780,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13338.4]
  assign _T_795 = {_T_781,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13340.4]
  assign _T_797 = {_T_782,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13342.4]
  assign _T_799 = {_T_783,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13344.4]
  assign _T_801 = {_T_784,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13346.4]
  assign _T_803 = {_T_785,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13348.4]
  assign _T_804 = _T_784 ? _T_801 : _T_803; // @[Mux.scala 31:69:@13349.4]
  assign _T_805 = _T_783 ? _T_799 : _T_804; // @[Mux.scala 31:69:@13350.4]
  assign _T_806 = _T_782 ? _T_797 : _T_805; // @[Mux.scala 31:69:@13351.4]
  assign _T_807 = _T_781 ? _T_795 : _T_806; // @[Mux.scala 31:69:@13352.4]
  assign _T_808 = _T_780 ? _T_793 : _T_807; // @[Mux.scala 31:69:@13353.4]
  assign _T_809 = _T_779 ? _T_791 : _T_808; // @[Mux.scala 31:69:@13354.4]
  assign _T_810 = _T_778 ? _T_789 : _T_809; // @[Mux.scala 31:69:@13355.4]
  assign _T_811 = _T_777 ? _T_787 : _T_810; // @[Mux.scala 31:69:@13356.4]
  assign _T_819 = _T_724 & _T_542; // @[MemPrimitives.scala 110:228:@13365.4]
  assign _T_825 = _T_730 & _T_548; // @[MemPrimitives.scala 110:228:@13369.4]
  assign _T_831 = _T_736 & _T_554; // @[MemPrimitives.scala 110:228:@13373.4]
  assign _T_837 = _T_742 & _T_560; // @[MemPrimitives.scala 110:228:@13377.4]
  assign _T_843 = _T_748 & _T_566; // @[MemPrimitives.scala 110:228:@13381.4]
  assign _T_849 = _T_754 & _T_572; // @[MemPrimitives.scala 110:228:@13385.4]
  assign _T_855 = _T_760 & _T_578; // @[MemPrimitives.scala 110:228:@13389.4]
  assign _T_861 = _T_766 & _T_584; // @[MemPrimitives.scala 110:228:@13393.4]
  assign _T_867 = _T_772 & _T_590; // @[MemPrimitives.scala 110:228:@13397.4]
  assign _T_869 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 126:35:@13411.4]
  assign _T_870 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 126:35:@13412.4]
  assign _T_871 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 126:35:@13413.4]
  assign _T_872 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 126:35:@13414.4]
  assign _T_873 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 126:35:@13415.4]
  assign _T_874 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 126:35:@13416.4]
  assign _T_875 = StickySelects_4_io_outs_6; // @[MemPrimitives.scala 126:35:@13417.4]
  assign _T_876 = StickySelects_4_io_outs_7; // @[MemPrimitives.scala 126:35:@13418.4]
  assign _T_877 = StickySelects_4_io_outs_8; // @[MemPrimitives.scala 126:35:@13419.4]
  assign _T_879 = {_T_869,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13421.4]
  assign _T_881 = {_T_870,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13423.4]
  assign _T_883 = {_T_871,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13425.4]
  assign _T_885 = {_T_872,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13427.4]
  assign _T_887 = {_T_873,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13429.4]
  assign _T_889 = {_T_874,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13431.4]
  assign _T_891 = {_T_875,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13433.4]
  assign _T_893 = {_T_876,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13435.4]
  assign _T_895 = {_T_877,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13437.4]
  assign _T_896 = _T_876 ? _T_893 : _T_895; // @[Mux.scala 31:69:@13438.4]
  assign _T_897 = _T_875 ? _T_891 : _T_896; // @[Mux.scala 31:69:@13439.4]
  assign _T_898 = _T_874 ? _T_889 : _T_897; // @[Mux.scala 31:69:@13440.4]
  assign _T_899 = _T_873 ? _T_887 : _T_898; // @[Mux.scala 31:69:@13441.4]
  assign _T_900 = _T_872 ? _T_885 : _T_899; // @[Mux.scala 31:69:@13442.4]
  assign _T_901 = _T_871 ? _T_883 : _T_900; // @[Mux.scala 31:69:@13443.4]
  assign _T_902 = _T_870 ? _T_881 : _T_901; // @[Mux.scala 31:69:@13444.4]
  assign _T_903 = _T_869 ? _T_879 : _T_902; // @[Mux.scala 31:69:@13445.4]
  assign _T_911 = _T_724 & _T_634; // @[MemPrimitives.scala 110:228:@13454.4]
  assign _T_917 = _T_730 & _T_640; // @[MemPrimitives.scala 110:228:@13458.4]
  assign _T_923 = _T_736 & _T_646; // @[MemPrimitives.scala 110:228:@13462.4]
  assign _T_929 = _T_742 & _T_652; // @[MemPrimitives.scala 110:228:@13466.4]
  assign _T_935 = _T_748 & _T_658; // @[MemPrimitives.scala 110:228:@13470.4]
  assign _T_941 = _T_754 & _T_664; // @[MemPrimitives.scala 110:228:@13474.4]
  assign _T_947 = _T_760 & _T_670; // @[MemPrimitives.scala 110:228:@13478.4]
  assign _T_953 = _T_766 & _T_676; // @[MemPrimitives.scala 110:228:@13482.4]
  assign _T_959 = _T_772 & _T_682; // @[MemPrimitives.scala 110:228:@13486.4]
  assign _T_961 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 126:35:@13500.4]
  assign _T_962 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 126:35:@13501.4]
  assign _T_963 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 126:35:@13502.4]
  assign _T_964 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 126:35:@13503.4]
  assign _T_965 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 126:35:@13504.4]
  assign _T_966 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 126:35:@13505.4]
  assign _T_967 = StickySelects_5_io_outs_6; // @[MemPrimitives.scala 126:35:@13506.4]
  assign _T_968 = StickySelects_5_io_outs_7; // @[MemPrimitives.scala 126:35:@13507.4]
  assign _T_969 = StickySelects_5_io_outs_8; // @[MemPrimitives.scala 126:35:@13508.4]
  assign _T_971 = {_T_961,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13510.4]
  assign _T_973 = {_T_962,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13512.4]
  assign _T_975 = {_T_963,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13514.4]
  assign _T_977 = {_T_964,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13516.4]
  assign _T_979 = {_T_965,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13518.4]
  assign _T_981 = {_T_966,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13520.4]
  assign _T_983 = {_T_967,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13522.4]
  assign _T_985 = {_T_968,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13524.4]
  assign _T_987 = {_T_969,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13526.4]
  assign _T_988 = _T_968 ? _T_985 : _T_987; // @[Mux.scala 31:69:@13527.4]
  assign _T_989 = _T_967 ? _T_983 : _T_988; // @[Mux.scala 31:69:@13528.4]
  assign _T_990 = _T_966 ? _T_981 : _T_989; // @[Mux.scala 31:69:@13529.4]
  assign _T_991 = _T_965 ? _T_979 : _T_990; // @[Mux.scala 31:69:@13530.4]
  assign _T_992 = _T_964 ? _T_977 : _T_991; // @[Mux.scala 31:69:@13531.4]
  assign _T_993 = _T_963 ? _T_975 : _T_992; // @[Mux.scala 31:69:@13532.4]
  assign _T_994 = _T_962 ? _T_973 : _T_993; // @[Mux.scala 31:69:@13533.4]
  assign _T_995 = _T_961 ? _T_971 : _T_994; // @[Mux.scala 31:69:@13534.4]
  assign _T_1000 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13541.4]
  assign _T_1003 = _T_1000 & _T_450; // @[MemPrimitives.scala 110:228:@13543.4]
  assign _T_1006 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13545.4]
  assign _T_1009 = _T_1006 & _T_456; // @[MemPrimitives.scala 110:228:@13547.4]
  assign _T_1012 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13549.4]
  assign _T_1015 = _T_1012 & _T_462; // @[MemPrimitives.scala 110:228:@13551.4]
  assign _T_1018 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13553.4]
  assign _T_1021 = _T_1018 & _T_468; // @[MemPrimitives.scala 110:228:@13555.4]
  assign _T_1024 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13557.4]
  assign _T_1027 = _T_1024 & _T_474; // @[MemPrimitives.scala 110:228:@13559.4]
  assign _T_1030 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13561.4]
  assign _T_1033 = _T_1030 & _T_480; // @[MemPrimitives.scala 110:228:@13563.4]
  assign _T_1036 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13565.4]
  assign _T_1039 = _T_1036 & _T_486; // @[MemPrimitives.scala 110:228:@13567.4]
  assign _T_1042 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13569.4]
  assign _T_1045 = _T_1042 & _T_492; // @[MemPrimitives.scala 110:228:@13571.4]
  assign _T_1048 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13573.4]
  assign _T_1051 = _T_1048 & _T_498; // @[MemPrimitives.scala 110:228:@13575.4]
  assign _T_1053 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 126:35:@13589.4]
  assign _T_1054 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 126:35:@13590.4]
  assign _T_1055 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 126:35:@13591.4]
  assign _T_1056 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 126:35:@13592.4]
  assign _T_1057 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 126:35:@13593.4]
  assign _T_1058 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 126:35:@13594.4]
  assign _T_1059 = StickySelects_6_io_outs_6; // @[MemPrimitives.scala 126:35:@13595.4]
  assign _T_1060 = StickySelects_6_io_outs_7; // @[MemPrimitives.scala 126:35:@13596.4]
  assign _T_1061 = StickySelects_6_io_outs_8; // @[MemPrimitives.scala 126:35:@13597.4]
  assign _T_1063 = {_T_1053,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13599.4]
  assign _T_1065 = {_T_1054,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13601.4]
  assign _T_1067 = {_T_1055,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13603.4]
  assign _T_1069 = {_T_1056,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13605.4]
  assign _T_1071 = {_T_1057,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13607.4]
  assign _T_1073 = {_T_1058,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13609.4]
  assign _T_1075 = {_T_1059,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13611.4]
  assign _T_1077 = {_T_1060,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13613.4]
  assign _T_1079 = {_T_1061,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13615.4]
  assign _T_1080 = _T_1060 ? _T_1077 : _T_1079; // @[Mux.scala 31:69:@13616.4]
  assign _T_1081 = _T_1059 ? _T_1075 : _T_1080; // @[Mux.scala 31:69:@13617.4]
  assign _T_1082 = _T_1058 ? _T_1073 : _T_1081; // @[Mux.scala 31:69:@13618.4]
  assign _T_1083 = _T_1057 ? _T_1071 : _T_1082; // @[Mux.scala 31:69:@13619.4]
  assign _T_1084 = _T_1056 ? _T_1069 : _T_1083; // @[Mux.scala 31:69:@13620.4]
  assign _T_1085 = _T_1055 ? _T_1067 : _T_1084; // @[Mux.scala 31:69:@13621.4]
  assign _T_1086 = _T_1054 ? _T_1065 : _T_1085; // @[Mux.scala 31:69:@13622.4]
  assign _T_1087 = _T_1053 ? _T_1063 : _T_1086; // @[Mux.scala 31:69:@13623.4]
  assign _T_1095 = _T_1000 & _T_542; // @[MemPrimitives.scala 110:228:@13632.4]
  assign _T_1101 = _T_1006 & _T_548; // @[MemPrimitives.scala 110:228:@13636.4]
  assign _T_1107 = _T_1012 & _T_554; // @[MemPrimitives.scala 110:228:@13640.4]
  assign _T_1113 = _T_1018 & _T_560; // @[MemPrimitives.scala 110:228:@13644.4]
  assign _T_1119 = _T_1024 & _T_566; // @[MemPrimitives.scala 110:228:@13648.4]
  assign _T_1125 = _T_1030 & _T_572; // @[MemPrimitives.scala 110:228:@13652.4]
  assign _T_1131 = _T_1036 & _T_578; // @[MemPrimitives.scala 110:228:@13656.4]
  assign _T_1137 = _T_1042 & _T_584; // @[MemPrimitives.scala 110:228:@13660.4]
  assign _T_1143 = _T_1048 & _T_590; // @[MemPrimitives.scala 110:228:@13664.4]
  assign _T_1145 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 126:35:@13678.4]
  assign _T_1146 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 126:35:@13679.4]
  assign _T_1147 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 126:35:@13680.4]
  assign _T_1148 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 126:35:@13681.4]
  assign _T_1149 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 126:35:@13682.4]
  assign _T_1150 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 126:35:@13683.4]
  assign _T_1151 = StickySelects_7_io_outs_6; // @[MemPrimitives.scala 126:35:@13684.4]
  assign _T_1152 = StickySelects_7_io_outs_7; // @[MemPrimitives.scala 126:35:@13685.4]
  assign _T_1153 = StickySelects_7_io_outs_8; // @[MemPrimitives.scala 126:35:@13686.4]
  assign _T_1155 = {_T_1145,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13688.4]
  assign _T_1157 = {_T_1146,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13690.4]
  assign _T_1159 = {_T_1147,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13692.4]
  assign _T_1161 = {_T_1148,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13694.4]
  assign _T_1163 = {_T_1149,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13696.4]
  assign _T_1165 = {_T_1150,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13698.4]
  assign _T_1167 = {_T_1151,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13700.4]
  assign _T_1169 = {_T_1152,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13702.4]
  assign _T_1171 = {_T_1153,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13704.4]
  assign _T_1172 = _T_1152 ? _T_1169 : _T_1171; // @[Mux.scala 31:69:@13705.4]
  assign _T_1173 = _T_1151 ? _T_1167 : _T_1172; // @[Mux.scala 31:69:@13706.4]
  assign _T_1174 = _T_1150 ? _T_1165 : _T_1173; // @[Mux.scala 31:69:@13707.4]
  assign _T_1175 = _T_1149 ? _T_1163 : _T_1174; // @[Mux.scala 31:69:@13708.4]
  assign _T_1176 = _T_1148 ? _T_1161 : _T_1175; // @[Mux.scala 31:69:@13709.4]
  assign _T_1177 = _T_1147 ? _T_1159 : _T_1176; // @[Mux.scala 31:69:@13710.4]
  assign _T_1178 = _T_1146 ? _T_1157 : _T_1177; // @[Mux.scala 31:69:@13711.4]
  assign _T_1179 = _T_1145 ? _T_1155 : _T_1178; // @[Mux.scala 31:69:@13712.4]
  assign _T_1187 = _T_1000 & _T_634; // @[MemPrimitives.scala 110:228:@13721.4]
  assign _T_1193 = _T_1006 & _T_640; // @[MemPrimitives.scala 110:228:@13725.4]
  assign _T_1199 = _T_1012 & _T_646; // @[MemPrimitives.scala 110:228:@13729.4]
  assign _T_1205 = _T_1018 & _T_652; // @[MemPrimitives.scala 110:228:@13733.4]
  assign _T_1211 = _T_1024 & _T_658; // @[MemPrimitives.scala 110:228:@13737.4]
  assign _T_1217 = _T_1030 & _T_664; // @[MemPrimitives.scala 110:228:@13741.4]
  assign _T_1223 = _T_1036 & _T_670; // @[MemPrimitives.scala 110:228:@13745.4]
  assign _T_1229 = _T_1042 & _T_676; // @[MemPrimitives.scala 110:228:@13749.4]
  assign _T_1235 = _T_1048 & _T_682; // @[MemPrimitives.scala 110:228:@13753.4]
  assign _T_1237 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 126:35:@13767.4]
  assign _T_1238 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 126:35:@13768.4]
  assign _T_1239 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 126:35:@13769.4]
  assign _T_1240 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 126:35:@13770.4]
  assign _T_1241 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 126:35:@13771.4]
  assign _T_1242 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 126:35:@13772.4]
  assign _T_1243 = StickySelects_8_io_outs_6; // @[MemPrimitives.scala 126:35:@13773.4]
  assign _T_1244 = StickySelects_8_io_outs_7; // @[MemPrimitives.scala 126:35:@13774.4]
  assign _T_1245 = StickySelects_8_io_outs_8; // @[MemPrimitives.scala 126:35:@13775.4]
  assign _T_1247 = {_T_1237,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13777.4]
  assign _T_1249 = {_T_1238,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13779.4]
  assign _T_1251 = {_T_1239,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13781.4]
  assign _T_1253 = {_T_1240,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13783.4]
  assign _T_1255 = {_T_1241,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13785.4]
  assign _T_1257 = {_T_1242,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13787.4]
  assign _T_1259 = {_T_1243,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13789.4]
  assign _T_1261 = {_T_1244,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13791.4]
  assign _T_1263 = {_T_1245,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13793.4]
  assign _T_1264 = _T_1244 ? _T_1261 : _T_1263; // @[Mux.scala 31:69:@13794.4]
  assign _T_1265 = _T_1243 ? _T_1259 : _T_1264; // @[Mux.scala 31:69:@13795.4]
  assign _T_1266 = _T_1242 ? _T_1257 : _T_1265; // @[Mux.scala 31:69:@13796.4]
  assign _T_1267 = _T_1241 ? _T_1255 : _T_1266; // @[Mux.scala 31:69:@13797.4]
  assign _T_1268 = _T_1240 ? _T_1253 : _T_1267; // @[Mux.scala 31:69:@13798.4]
  assign _T_1269 = _T_1239 ? _T_1251 : _T_1268; // @[Mux.scala 31:69:@13799.4]
  assign _T_1270 = _T_1238 ? _T_1249 : _T_1269; // @[Mux.scala 31:69:@13800.4]
  assign _T_1271 = _T_1237 ? _T_1247 : _T_1270; // @[Mux.scala 31:69:@13801.4]
  assign _T_1276 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13808.4]
  assign _T_1279 = _T_1276 & _T_450; // @[MemPrimitives.scala 110:228:@13810.4]
  assign _T_1282 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13812.4]
  assign _T_1285 = _T_1282 & _T_456; // @[MemPrimitives.scala 110:228:@13814.4]
  assign _T_1288 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13816.4]
  assign _T_1291 = _T_1288 & _T_462; // @[MemPrimitives.scala 110:228:@13818.4]
  assign _T_1294 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13820.4]
  assign _T_1297 = _T_1294 & _T_468; // @[MemPrimitives.scala 110:228:@13822.4]
  assign _T_1300 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13824.4]
  assign _T_1303 = _T_1300 & _T_474; // @[MemPrimitives.scala 110:228:@13826.4]
  assign _T_1306 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13828.4]
  assign _T_1309 = _T_1306 & _T_480; // @[MemPrimitives.scala 110:228:@13830.4]
  assign _T_1312 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13832.4]
  assign _T_1315 = _T_1312 & _T_486; // @[MemPrimitives.scala 110:228:@13834.4]
  assign _T_1318 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13836.4]
  assign _T_1321 = _T_1318 & _T_492; // @[MemPrimitives.scala 110:228:@13838.4]
  assign _T_1324 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13840.4]
  assign _T_1327 = _T_1324 & _T_498; // @[MemPrimitives.scala 110:228:@13842.4]
  assign _T_1329 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 126:35:@13856.4]
  assign _T_1330 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 126:35:@13857.4]
  assign _T_1331 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 126:35:@13858.4]
  assign _T_1332 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 126:35:@13859.4]
  assign _T_1333 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 126:35:@13860.4]
  assign _T_1334 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 126:35:@13861.4]
  assign _T_1335 = StickySelects_9_io_outs_6; // @[MemPrimitives.scala 126:35:@13862.4]
  assign _T_1336 = StickySelects_9_io_outs_7; // @[MemPrimitives.scala 126:35:@13863.4]
  assign _T_1337 = StickySelects_9_io_outs_8; // @[MemPrimitives.scala 126:35:@13864.4]
  assign _T_1339 = {_T_1329,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13866.4]
  assign _T_1341 = {_T_1330,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13868.4]
  assign _T_1343 = {_T_1331,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13870.4]
  assign _T_1345 = {_T_1332,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13872.4]
  assign _T_1347 = {_T_1333,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13874.4]
  assign _T_1349 = {_T_1334,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13876.4]
  assign _T_1351 = {_T_1335,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13878.4]
  assign _T_1353 = {_T_1336,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13880.4]
  assign _T_1355 = {_T_1337,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13882.4]
  assign _T_1356 = _T_1336 ? _T_1353 : _T_1355; // @[Mux.scala 31:69:@13883.4]
  assign _T_1357 = _T_1335 ? _T_1351 : _T_1356; // @[Mux.scala 31:69:@13884.4]
  assign _T_1358 = _T_1334 ? _T_1349 : _T_1357; // @[Mux.scala 31:69:@13885.4]
  assign _T_1359 = _T_1333 ? _T_1347 : _T_1358; // @[Mux.scala 31:69:@13886.4]
  assign _T_1360 = _T_1332 ? _T_1345 : _T_1359; // @[Mux.scala 31:69:@13887.4]
  assign _T_1361 = _T_1331 ? _T_1343 : _T_1360; // @[Mux.scala 31:69:@13888.4]
  assign _T_1362 = _T_1330 ? _T_1341 : _T_1361; // @[Mux.scala 31:69:@13889.4]
  assign _T_1363 = _T_1329 ? _T_1339 : _T_1362; // @[Mux.scala 31:69:@13890.4]
  assign _T_1371 = _T_1276 & _T_542; // @[MemPrimitives.scala 110:228:@13899.4]
  assign _T_1377 = _T_1282 & _T_548; // @[MemPrimitives.scala 110:228:@13903.4]
  assign _T_1383 = _T_1288 & _T_554; // @[MemPrimitives.scala 110:228:@13907.4]
  assign _T_1389 = _T_1294 & _T_560; // @[MemPrimitives.scala 110:228:@13911.4]
  assign _T_1395 = _T_1300 & _T_566; // @[MemPrimitives.scala 110:228:@13915.4]
  assign _T_1401 = _T_1306 & _T_572; // @[MemPrimitives.scala 110:228:@13919.4]
  assign _T_1407 = _T_1312 & _T_578; // @[MemPrimitives.scala 110:228:@13923.4]
  assign _T_1413 = _T_1318 & _T_584; // @[MemPrimitives.scala 110:228:@13927.4]
  assign _T_1419 = _T_1324 & _T_590; // @[MemPrimitives.scala 110:228:@13931.4]
  assign _T_1421 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 126:35:@13945.4]
  assign _T_1422 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 126:35:@13946.4]
  assign _T_1423 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 126:35:@13947.4]
  assign _T_1424 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 126:35:@13948.4]
  assign _T_1425 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 126:35:@13949.4]
  assign _T_1426 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 126:35:@13950.4]
  assign _T_1427 = StickySelects_10_io_outs_6; // @[MemPrimitives.scala 126:35:@13951.4]
  assign _T_1428 = StickySelects_10_io_outs_7; // @[MemPrimitives.scala 126:35:@13952.4]
  assign _T_1429 = StickySelects_10_io_outs_8; // @[MemPrimitives.scala 126:35:@13953.4]
  assign _T_1431 = {_T_1421,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13955.4]
  assign _T_1433 = {_T_1422,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13957.4]
  assign _T_1435 = {_T_1423,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13959.4]
  assign _T_1437 = {_T_1424,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13961.4]
  assign _T_1439 = {_T_1425,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13963.4]
  assign _T_1441 = {_T_1426,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13965.4]
  assign _T_1443 = {_T_1427,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13967.4]
  assign _T_1445 = {_T_1428,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13969.4]
  assign _T_1447 = {_T_1429,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13971.4]
  assign _T_1448 = _T_1428 ? _T_1445 : _T_1447; // @[Mux.scala 31:69:@13972.4]
  assign _T_1449 = _T_1427 ? _T_1443 : _T_1448; // @[Mux.scala 31:69:@13973.4]
  assign _T_1450 = _T_1426 ? _T_1441 : _T_1449; // @[Mux.scala 31:69:@13974.4]
  assign _T_1451 = _T_1425 ? _T_1439 : _T_1450; // @[Mux.scala 31:69:@13975.4]
  assign _T_1452 = _T_1424 ? _T_1437 : _T_1451; // @[Mux.scala 31:69:@13976.4]
  assign _T_1453 = _T_1423 ? _T_1435 : _T_1452; // @[Mux.scala 31:69:@13977.4]
  assign _T_1454 = _T_1422 ? _T_1433 : _T_1453; // @[Mux.scala 31:69:@13978.4]
  assign _T_1455 = _T_1421 ? _T_1431 : _T_1454; // @[Mux.scala 31:69:@13979.4]
  assign _T_1463 = _T_1276 & _T_634; // @[MemPrimitives.scala 110:228:@13988.4]
  assign _T_1469 = _T_1282 & _T_640; // @[MemPrimitives.scala 110:228:@13992.4]
  assign _T_1475 = _T_1288 & _T_646; // @[MemPrimitives.scala 110:228:@13996.4]
  assign _T_1481 = _T_1294 & _T_652; // @[MemPrimitives.scala 110:228:@14000.4]
  assign _T_1487 = _T_1300 & _T_658; // @[MemPrimitives.scala 110:228:@14004.4]
  assign _T_1493 = _T_1306 & _T_664; // @[MemPrimitives.scala 110:228:@14008.4]
  assign _T_1499 = _T_1312 & _T_670; // @[MemPrimitives.scala 110:228:@14012.4]
  assign _T_1505 = _T_1318 & _T_676; // @[MemPrimitives.scala 110:228:@14016.4]
  assign _T_1511 = _T_1324 & _T_682; // @[MemPrimitives.scala 110:228:@14020.4]
  assign _T_1513 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 126:35:@14034.4]
  assign _T_1514 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 126:35:@14035.4]
  assign _T_1515 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 126:35:@14036.4]
  assign _T_1516 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 126:35:@14037.4]
  assign _T_1517 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 126:35:@14038.4]
  assign _T_1518 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 126:35:@14039.4]
  assign _T_1519 = StickySelects_11_io_outs_6; // @[MemPrimitives.scala 126:35:@14040.4]
  assign _T_1520 = StickySelects_11_io_outs_7; // @[MemPrimitives.scala 126:35:@14041.4]
  assign _T_1521 = StickySelects_11_io_outs_8; // @[MemPrimitives.scala 126:35:@14042.4]
  assign _T_1523 = {_T_1513,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@14044.4]
  assign _T_1525 = {_T_1514,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@14046.4]
  assign _T_1527 = {_T_1515,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@14048.4]
  assign _T_1529 = {_T_1516,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@14050.4]
  assign _T_1531 = {_T_1517,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@14052.4]
  assign _T_1533 = {_T_1518,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@14054.4]
  assign _T_1535 = {_T_1519,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@14056.4]
  assign _T_1537 = {_T_1520,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@14058.4]
  assign _T_1539 = {_T_1521,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@14060.4]
  assign _T_1540 = _T_1520 ? _T_1537 : _T_1539; // @[Mux.scala 31:69:@14061.4]
  assign _T_1541 = _T_1519 ? _T_1535 : _T_1540; // @[Mux.scala 31:69:@14062.4]
  assign _T_1542 = _T_1518 ? _T_1533 : _T_1541; // @[Mux.scala 31:69:@14063.4]
  assign _T_1543 = _T_1517 ? _T_1531 : _T_1542; // @[Mux.scala 31:69:@14064.4]
  assign _T_1544 = _T_1516 ? _T_1529 : _T_1543; // @[Mux.scala 31:69:@14065.4]
  assign _T_1545 = _T_1515 ? _T_1527 : _T_1544; // @[Mux.scala 31:69:@14066.4]
  assign _T_1546 = _T_1514 ? _T_1525 : _T_1545; // @[Mux.scala 31:69:@14067.4]
  assign _T_1547 = _T_1513 ? _T_1523 : _T_1546; // @[Mux.scala 31:69:@14068.4]
  assign _T_1643 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@14197.4 package.scala 96:25:@14198.4]
  assign _T_1647 = _T_1643 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14207.4]
  assign _T_1640 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@14189.4 package.scala 96:25:@14190.4]
  assign _T_1648 = _T_1640 ? Mem1D_9_io_output : _T_1647; // @[Mux.scala 31:69:@14208.4]
  assign _T_1637 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@14181.4 package.scala 96:25:@14182.4]
  assign _T_1649 = _T_1637 ? Mem1D_8_io_output : _T_1648; // @[Mux.scala 31:69:@14209.4]
  assign _T_1634 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@14173.4 package.scala 96:25:@14174.4]
  assign _T_1650 = _T_1634 ? Mem1D_7_io_output : _T_1649; // @[Mux.scala 31:69:@14210.4]
  assign _T_1631 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@14165.4 package.scala 96:25:@14166.4]
  assign _T_1651 = _T_1631 ? Mem1D_6_io_output : _T_1650; // @[Mux.scala 31:69:@14211.4]
  assign _T_1628 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@14157.4 package.scala 96:25:@14158.4]
  assign _T_1652 = _T_1628 ? Mem1D_5_io_output : _T_1651; // @[Mux.scala 31:69:@14212.4]
  assign _T_1625 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@14149.4 package.scala 96:25:@14150.4]
  assign _T_1653 = _T_1625 ? Mem1D_4_io_output : _T_1652; // @[Mux.scala 31:69:@14213.4]
  assign _T_1622 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@14141.4 package.scala 96:25:@14142.4]
  assign _T_1654 = _T_1622 ? Mem1D_3_io_output : _T_1653; // @[Mux.scala 31:69:@14214.4]
  assign _T_1619 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@14133.4 package.scala 96:25:@14134.4]
  assign _T_1655 = _T_1619 ? Mem1D_2_io_output : _T_1654; // @[Mux.scala 31:69:@14215.4]
  assign _T_1616 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@14125.4 package.scala 96:25:@14126.4]
  assign _T_1656 = _T_1616 ? Mem1D_1_io_output : _T_1655; // @[Mux.scala 31:69:@14216.4]
  assign _T_1613 = RetimeWrapper_io_out; // @[package.scala 96:25:@14117.4 package.scala 96:25:@14118.4]
  assign _T_1750 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@14341.4 package.scala 96:25:@14342.4]
  assign _T_1754 = _T_1750 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14351.4]
  assign _T_1747 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@14333.4 package.scala 96:25:@14334.4]
  assign _T_1755 = _T_1747 ? Mem1D_9_io_output : _T_1754; // @[Mux.scala 31:69:@14352.4]
  assign _T_1744 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@14325.4 package.scala 96:25:@14326.4]
  assign _T_1756 = _T_1744 ? Mem1D_8_io_output : _T_1755; // @[Mux.scala 31:69:@14353.4]
  assign _T_1741 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@14317.4 package.scala 96:25:@14318.4]
  assign _T_1757 = _T_1741 ? Mem1D_7_io_output : _T_1756; // @[Mux.scala 31:69:@14354.4]
  assign _T_1738 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@14309.4 package.scala 96:25:@14310.4]
  assign _T_1758 = _T_1738 ? Mem1D_6_io_output : _T_1757; // @[Mux.scala 31:69:@14355.4]
  assign _T_1735 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@14301.4 package.scala 96:25:@14302.4]
  assign _T_1759 = _T_1735 ? Mem1D_5_io_output : _T_1758; // @[Mux.scala 31:69:@14356.4]
  assign _T_1732 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@14293.4 package.scala 96:25:@14294.4]
  assign _T_1760 = _T_1732 ? Mem1D_4_io_output : _T_1759; // @[Mux.scala 31:69:@14357.4]
  assign _T_1729 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@14285.4 package.scala 96:25:@14286.4]
  assign _T_1761 = _T_1729 ? Mem1D_3_io_output : _T_1760; // @[Mux.scala 31:69:@14358.4]
  assign _T_1726 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@14277.4 package.scala 96:25:@14278.4]
  assign _T_1762 = _T_1726 ? Mem1D_2_io_output : _T_1761; // @[Mux.scala 31:69:@14359.4]
  assign _T_1723 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@14269.4 package.scala 96:25:@14270.4]
  assign _T_1763 = _T_1723 ? Mem1D_1_io_output : _T_1762; // @[Mux.scala 31:69:@14360.4]
  assign _T_1720 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@14261.4 package.scala 96:25:@14262.4]
  assign _T_1857 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@14485.4 package.scala 96:25:@14486.4]
  assign _T_1861 = _T_1857 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14495.4]
  assign _T_1854 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@14477.4 package.scala 96:25:@14478.4]
  assign _T_1862 = _T_1854 ? Mem1D_9_io_output : _T_1861; // @[Mux.scala 31:69:@14496.4]
  assign _T_1851 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@14469.4 package.scala 96:25:@14470.4]
  assign _T_1863 = _T_1851 ? Mem1D_8_io_output : _T_1862; // @[Mux.scala 31:69:@14497.4]
  assign _T_1848 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@14461.4 package.scala 96:25:@14462.4]
  assign _T_1864 = _T_1848 ? Mem1D_7_io_output : _T_1863; // @[Mux.scala 31:69:@14498.4]
  assign _T_1845 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@14453.4 package.scala 96:25:@14454.4]
  assign _T_1865 = _T_1845 ? Mem1D_6_io_output : _T_1864; // @[Mux.scala 31:69:@14499.4]
  assign _T_1842 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@14445.4 package.scala 96:25:@14446.4]
  assign _T_1866 = _T_1842 ? Mem1D_5_io_output : _T_1865; // @[Mux.scala 31:69:@14500.4]
  assign _T_1839 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@14437.4 package.scala 96:25:@14438.4]
  assign _T_1867 = _T_1839 ? Mem1D_4_io_output : _T_1866; // @[Mux.scala 31:69:@14501.4]
  assign _T_1836 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@14429.4 package.scala 96:25:@14430.4]
  assign _T_1868 = _T_1836 ? Mem1D_3_io_output : _T_1867; // @[Mux.scala 31:69:@14502.4]
  assign _T_1833 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@14421.4 package.scala 96:25:@14422.4]
  assign _T_1869 = _T_1833 ? Mem1D_2_io_output : _T_1868; // @[Mux.scala 31:69:@14503.4]
  assign _T_1830 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@14413.4 package.scala 96:25:@14414.4]
  assign _T_1870 = _T_1830 ? Mem1D_1_io_output : _T_1869; // @[Mux.scala 31:69:@14504.4]
  assign _T_1827 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@14405.4 package.scala 96:25:@14406.4]
  assign _T_1964 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@14629.4 package.scala 96:25:@14630.4]
  assign _T_1968 = _T_1964 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14639.4]
  assign _T_1961 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@14621.4 package.scala 96:25:@14622.4]
  assign _T_1969 = _T_1961 ? Mem1D_9_io_output : _T_1968; // @[Mux.scala 31:69:@14640.4]
  assign _T_1958 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@14613.4 package.scala 96:25:@14614.4]
  assign _T_1970 = _T_1958 ? Mem1D_8_io_output : _T_1969; // @[Mux.scala 31:69:@14641.4]
  assign _T_1955 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@14605.4 package.scala 96:25:@14606.4]
  assign _T_1971 = _T_1955 ? Mem1D_7_io_output : _T_1970; // @[Mux.scala 31:69:@14642.4]
  assign _T_1952 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@14597.4 package.scala 96:25:@14598.4]
  assign _T_1972 = _T_1952 ? Mem1D_6_io_output : _T_1971; // @[Mux.scala 31:69:@14643.4]
  assign _T_1949 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@14589.4 package.scala 96:25:@14590.4]
  assign _T_1973 = _T_1949 ? Mem1D_5_io_output : _T_1972; // @[Mux.scala 31:69:@14644.4]
  assign _T_1946 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@14581.4 package.scala 96:25:@14582.4]
  assign _T_1974 = _T_1946 ? Mem1D_4_io_output : _T_1973; // @[Mux.scala 31:69:@14645.4]
  assign _T_1943 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@14573.4 package.scala 96:25:@14574.4]
  assign _T_1975 = _T_1943 ? Mem1D_3_io_output : _T_1974; // @[Mux.scala 31:69:@14646.4]
  assign _T_1940 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@14565.4 package.scala 96:25:@14566.4]
  assign _T_1976 = _T_1940 ? Mem1D_2_io_output : _T_1975; // @[Mux.scala 31:69:@14647.4]
  assign _T_1937 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@14557.4 package.scala 96:25:@14558.4]
  assign _T_1977 = _T_1937 ? Mem1D_1_io_output : _T_1976; // @[Mux.scala 31:69:@14648.4]
  assign _T_1934 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@14549.4 package.scala 96:25:@14550.4]
  assign _T_2071 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@14773.4 package.scala 96:25:@14774.4]
  assign _T_2075 = _T_2071 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14783.4]
  assign _T_2068 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@14765.4 package.scala 96:25:@14766.4]
  assign _T_2076 = _T_2068 ? Mem1D_9_io_output : _T_2075; // @[Mux.scala 31:69:@14784.4]
  assign _T_2065 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@14757.4 package.scala 96:25:@14758.4]
  assign _T_2077 = _T_2065 ? Mem1D_8_io_output : _T_2076; // @[Mux.scala 31:69:@14785.4]
  assign _T_2062 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@14749.4 package.scala 96:25:@14750.4]
  assign _T_2078 = _T_2062 ? Mem1D_7_io_output : _T_2077; // @[Mux.scala 31:69:@14786.4]
  assign _T_2059 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@14741.4 package.scala 96:25:@14742.4]
  assign _T_2079 = _T_2059 ? Mem1D_6_io_output : _T_2078; // @[Mux.scala 31:69:@14787.4]
  assign _T_2056 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@14733.4 package.scala 96:25:@14734.4]
  assign _T_2080 = _T_2056 ? Mem1D_5_io_output : _T_2079; // @[Mux.scala 31:69:@14788.4]
  assign _T_2053 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@14725.4 package.scala 96:25:@14726.4]
  assign _T_2081 = _T_2053 ? Mem1D_4_io_output : _T_2080; // @[Mux.scala 31:69:@14789.4]
  assign _T_2050 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@14717.4 package.scala 96:25:@14718.4]
  assign _T_2082 = _T_2050 ? Mem1D_3_io_output : _T_2081; // @[Mux.scala 31:69:@14790.4]
  assign _T_2047 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@14709.4 package.scala 96:25:@14710.4]
  assign _T_2083 = _T_2047 ? Mem1D_2_io_output : _T_2082; // @[Mux.scala 31:69:@14791.4]
  assign _T_2044 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@14701.4 package.scala 96:25:@14702.4]
  assign _T_2084 = _T_2044 ? Mem1D_1_io_output : _T_2083; // @[Mux.scala 31:69:@14792.4]
  assign _T_2041 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@14693.4 package.scala 96:25:@14694.4]
  assign _T_2178 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@14917.4 package.scala 96:25:@14918.4]
  assign _T_2182 = _T_2178 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14927.4]
  assign _T_2175 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@14909.4 package.scala 96:25:@14910.4]
  assign _T_2183 = _T_2175 ? Mem1D_9_io_output : _T_2182; // @[Mux.scala 31:69:@14928.4]
  assign _T_2172 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@14901.4 package.scala 96:25:@14902.4]
  assign _T_2184 = _T_2172 ? Mem1D_8_io_output : _T_2183; // @[Mux.scala 31:69:@14929.4]
  assign _T_2169 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@14893.4 package.scala 96:25:@14894.4]
  assign _T_2185 = _T_2169 ? Mem1D_7_io_output : _T_2184; // @[Mux.scala 31:69:@14930.4]
  assign _T_2166 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@14885.4 package.scala 96:25:@14886.4]
  assign _T_2186 = _T_2166 ? Mem1D_6_io_output : _T_2185; // @[Mux.scala 31:69:@14931.4]
  assign _T_2163 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@14877.4 package.scala 96:25:@14878.4]
  assign _T_2187 = _T_2163 ? Mem1D_5_io_output : _T_2186; // @[Mux.scala 31:69:@14932.4]
  assign _T_2160 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@14869.4 package.scala 96:25:@14870.4]
  assign _T_2188 = _T_2160 ? Mem1D_4_io_output : _T_2187; // @[Mux.scala 31:69:@14933.4]
  assign _T_2157 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@14861.4 package.scala 96:25:@14862.4]
  assign _T_2189 = _T_2157 ? Mem1D_3_io_output : _T_2188; // @[Mux.scala 31:69:@14934.4]
  assign _T_2154 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@14853.4 package.scala 96:25:@14854.4]
  assign _T_2190 = _T_2154 ? Mem1D_2_io_output : _T_2189; // @[Mux.scala 31:69:@14935.4]
  assign _T_2151 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@14845.4 package.scala 96:25:@14846.4]
  assign _T_2191 = _T_2151 ? Mem1D_1_io_output : _T_2190; // @[Mux.scala 31:69:@14936.4]
  assign _T_2148 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@14837.4 package.scala 96:25:@14838.4]
  assign _T_2285 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@15061.4 package.scala 96:25:@15062.4]
  assign _T_2289 = _T_2285 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@15071.4]
  assign _T_2282 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@15053.4 package.scala 96:25:@15054.4]
  assign _T_2290 = _T_2282 ? Mem1D_9_io_output : _T_2289; // @[Mux.scala 31:69:@15072.4]
  assign _T_2279 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@15045.4 package.scala 96:25:@15046.4]
  assign _T_2291 = _T_2279 ? Mem1D_8_io_output : _T_2290; // @[Mux.scala 31:69:@15073.4]
  assign _T_2276 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@15037.4 package.scala 96:25:@15038.4]
  assign _T_2292 = _T_2276 ? Mem1D_7_io_output : _T_2291; // @[Mux.scala 31:69:@15074.4]
  assign _T_2273 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@15029.4 package.scala 96:25:@15030.4]
  assign _T_2293 = _T_2273 ? Mem1D_6_io_output : _T_2292; // @[Mux.scala 31:69:@15075.4]
  assign _T_2270 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@15021.4 package.scala 96:25:@15022.4]
  assign _T_2294 = _T_2270 ? Mem1D_5_io_output : _T_2293; // @[Mux.scala 31:69:@15076.4]
  assign _T_2267 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@15013.4 package.scala 96:25:@15014.4]
  assign _T_2295 = _T_2267 ? Mem1D_4_io_output : _T_2294; // @[Mux.scala 31:69:@15077.4]
  assign _T_2264 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@15005.4 package.scala 96:25:@15006.4]
  assign _T_2296 = _T_2264 ? Mem1D_3_io_output : _T_2295; // @[Mux.scala 31:69:@15078.4]
  assign _T_2261 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@14997.4 package.scala 96:25:@14998.4]
  assign _T_2297 = _T_2261 ? Mem1D_2_io_output : _T_2296; // @[Mux.scala 31:69:@15079.4]
  assign _T_2258 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@14989.4 package.scala 96:25:@14990.4]
  assign _T_2298 = _T_2258 ? Mem1D_1_io_output : _T_2297; // @[Mux.scala 31:69:@15080.4]
  assign _T_2255 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@14981.4 package.scala 96:25:@14982.4]
  assign _T_2392 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@15205.4 package.scala 96:25:@15206.4]
  assign _T_2396 = _T_2392 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@15215.4]
  assign _T_2389 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@15197.4 package.scala 96:25:@15198.4]
  assign _T_2397 = _T_2389 ? Mem1D_9_io_output : _T_2396; // @[Mux.scala 31:69:@15216.4]
  assign _T_2386 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@15189.4 package.scala 96:25:@15190.4]
  assign _T_2398 = _T_2386 ? Mem1D_8_io_output : _T_2397; // @[Mux.scala 31:69:@15217.4]
  assign _T_2383 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@15181.4 package.scala 96:25:@15182.4]
  assign _T_2399 = _T_2383 ? Mem1D_7_io_output : _T_2398; // @[Mux.scala 31:69:@15218.4]
  assign _T_2380 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@15173.4 package.scala 96:25:@15174.4]
  assign _T_2400 = _T_2380 ? Mem1D_6_io_output : _T_2399; // @[Mux.scala 31:69:@15219.4]
  assign _T_2377 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@15165.4 package.scala 96:25:@15166.4]
  assign _T_2401 = _T_2377 ? Mem1D_5_io_output : _T_2400; // @[Mux.scala 31:69:@15220.4]
  assign _T_2374 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@15157.4 package.scala 96:25:@15158.4]
  assign _T_2402 = _T_2374 ? Mem1D_4_io_output : _T_2401; // @[Mux.scala 31:69:@15221.4]
  assign _T_2371 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@15149.4 package.scala 96:25:@15150.4]
  assign _T_2403 = _T_2371 ? Mem1D_3_io_output : _T_2402; // @[Mux.scala 31:69:@15222.4]
  assign _T_2368 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@15141.4 package.scala 96:25:@15142.4]
  assign _T_2404 = _T_2368 ? Mem1D_2_io_output : _T_2403; // @[Mux.scala 31:69:@15223.4]
  assign _T_2365 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@15133.4 package.scala 96:25:@15134.4]
  assign _T_2405 = _T_2365 ? Mem1D_1_io_output : _T_2404; // @[Mux.scala 31:69:@15224.4]
  assign _T_2362 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@15125.4 package.scala 96:25:@15126.4]
  assign _T_2499 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@15349.4 package.scala 96:25:@15350.4]
  assign _T_2503 = _T_2499 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@15359.4]
  assign _T_2496 = RetimeWrapper_105_io_out; // @[package.scala 96:25:@15341.4 package.scala 96:25:@15342.4]
  assign _T_2504 = _T_2496 ? Mem1D_9_io_output : _T_2503; // @[Mux.scala 31:69:@15360.4]
  assign _T_2493 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@15333.4 package.scala 96:25:@15334.4]
  assign _T_2505 = _T_2493 ? Mem1D_8_io_output : _T_2504; // @[Mux.scala 31:69:@15361.4]
  assign _T_2490 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@15325.4 package.scala 96:25:@15326.4]
  assign _T_2506 = _T_2490 ? Mem1D_7_io_output : _T_2505; // @[Mux.scala 31:69:@15362.4]
  assign _T_2487 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@15317.4 package.scala 96:25:@15318.4]
  assign _T_2507 = _T_2487 ? Mem1D_6_io_output : _T_2506; // @[Mux.scala 31:69:@15363.4]
  assign _T_2484 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@15309.4 package.scala 96:25:@15310.4]
  assign _T_2508 = _T_2484 ? Mem1D_5_io_output : _T_2507; // @[Mux.scala 31:69:@15364.4]
  assign _T_2481 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@15301.4 package.scala 96:25:@15302.4]
  assign _T_2509 = _T_2481 ? Mem1D_4_io_output : _T_2508; // @[Mux.scala 31:69:@15365.4]
  assign _T_2478 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@15293.4 package.scala 96:25:@15294.4]
  assign _T_2510 = _T_2478 ? Mem1D_3_io_output : _T_2509; // @[Mux.scala 31:69:@15366.4]
  assign _T_2475 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@15285.4 package.scala 96:25:@15286.4]
  assign _T_2511 = _T_2475 ? Mem1D_2_io_output : _T_2510; // @[Mux.scala 31:69:@15367.4]
  assign _T_2472 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@15277.4 package.scala 96:25:@15278.4]
  assign _T_2512 = _T_2472 ? Mem1D_1_io_output : _T_2511; // @[Mux.scala 31:69:@15368.4]
  assign _T_2469 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@15269.4 package.scala 96:25:@15270.4]
  assign io_rPort_8_output_0 = _T_2469 ? Mem1D_io_output : _T_2512; // @[MemPrimitives.scala 152:13:@15370.4]
  assign io_rPort_7_output_0 = _T_2362 ? Mem1D_io_output : _T_2405; // @[MemPrimitives.scala 152:13:@15226.4]
  assign io_rPort_6_output_0 = _T_2255 ? Mem1D_io_output : _T_2298; // @[MemPrimitives.scala 152:13:@15082.4]
  assign io_rPort_5_output_0 = _T_2148 ? Mem1D_io_output : _T_2191; // @[MemPrimitives.scala 152:13:@14938.4]
  assign io_rPort_4_output_0 = _T_2041 ? Mem1D_io_output : _T_2084; // @[MemPrimitives.scala 152:13:@14794.4]
  assign io_rPort_3_output_0 = _T_1934 ? Mem1D_io_output : _T_1977; // @[MemPrimitives.scala 152:13:@14650.4]
  assign io_rPort_2_output_0 = _T_1827 ? Mem1D_io_output : _T_1870; // @[MemPrimitives.scala 152:13:@14506.4]
  assign io_rPort_1_output_0 = _T_1720 ? Mem1D_io_output : _T_1763; // @[MemPrimitives.scala 152:13:@14362.4]
  assign io_rPort_0_output_0 = _T_1613 ? Mem1D_io_output : _T_1656; // @[MemPrimitives.scala 152:13:@14218.4]
  assign Mem1D_clock = clock; // @[:@12672.4]
  assign Mem1D_reset = reset; // @[:@12673.4]
  assign Mem1D_io_r_ofs_0 = _T_535[9:0]; // @[MemPrimitives.scala 131:28:@13093.4]
  assign Mem1D_io_r_backpressure = _T_535[10]; // @[MemPrimitives.scala 132:32:@13094.4]
  assign Mem1D_io_w_ofs_0 = _T_322[9:0]; // @[MemPrimitives.scala 94:28:@12872.4]
  assign Mem1D_io_w_data_0 = _T_322[41:10]; // @[MemPrimitives.scala 95:29:@12873.4]
  assign Mem1D_io_w_en_0 = _T_322[42]; // @[MemPrimitives.scala 96:27:@12874.4]
  assign Mem1D_1_clock = clock; // @[:@12688.4]
  assign Mem1D_1_reset = reset; // @[:@12689.4]
  assign Mem1D_1_io_r_ofs_0 = _T_627[9:0]; // @[MemPrimitives.scala 131:28:@13182.4]
  assign Mem1D_1_io_r_backpressure = _T_627[10]; // @[MemPrimitives.scala 132:32:@13183.4]
  assign Mem1D_1_io_w_ofs_0 = _T_333[9:0]; // @[MemPrimitives.scala 94:28:@12884.4]
  assign Mem1D_1_io_w_data_0 = _T_333[41:10]; // @[MemPrimitives.scala 95:29:@12885.4]
  assign Mem1D_1_io_w_en_0 = _T_333[42]; // @[MemPrimitives.scala 96:27:@12886.4]
  assign Mem1D_2_clock = clock; // @[:@12704.4]
  assign Mem1D_2_reset = reset; // @[:@12705.4]
  assign Mem1D_2_io_r_ofs_0 = _T_719[9:0]; // @[MemPrimitives.scala 131:28:@13271.4]
  assign Mem1D_2_io_r_backpressure = _T_719[10]; // @[MemPrimitives.scala 132:32:@13272.4]
  assign Mem1D_2_io_w_ofs_0 = _T_344[9:0]; // @[MemPrimitives.scala 94:28:@12896.4]
  assign Mem1D_2_io_w_data_0 = _T_344[41:10]; // @[MemPrimitives.scala 95:29:@12897.4]
  assign Mem1D_2_io_w_en_0 = _T_344[42]; // @[MemPrimitives.scala 96:27:@12898.4]
  assign Mem1D_3_clock = clock; // @[:@12720.4]
  assign Mem1D_3_reset = reset; // @[:@12721.4]
  assign Mem1D_3_io_r_ofs_0 = _T_811[9:0]; // @[MemPrimitives.scala 131:28:@13360.4]
  assign Mem1D_3_io_r_backpressure = _T_811[10]; // @[MemPrimitives.scala 132:32:@13361.4]
  assign Mem1D_3_io_w_ofs_0 = _T_355[9:0]; // @[MemPrimitives.scala 94:28:@12908.4]
  assign Mem1D_3_io_w_data_0 = _T_355[41:10]; // @[MemPrimitives.scala 95:29:@12909.4]
  assign Mem1D_3_io_w_en_0 = _T_355[42]; // @[MemPrimitives.scala 96:27:@12910.4]
  assign Mem1D_4_clock = clock; // @[:@12736.4]
  assign Mem1D_4_reset = reset; // @[:@12737.4]
  assign Mem1D_4_io_r_ofs_0 = _T_903[9:0]; // @[MemPrimitives.scala 131:28:@13449.4]
  assign Mem1D_4_io_r_backpressure = _T_903[10]; // @[MemPrimitives.scala 132:32:@13450.4]
  assign Mem1D_4_io_w_ofs_0 = _T_366[9:0]; // @[MemPrimitives.scala 94:28:@12920.4]
  assign Mem1D_4_io_w_data_0 = _T_366[41:10]; // @[MemPrimitives.scala 95:29:@12921.4]
  assign Mem1D_4_io_w_en_0 = _T_366[42]; // @[MemPrimitives.scala 96:27:@12922.4]
  assign Mem1D_5_clock = clock; // @[:@12752.4]
  assign Mem1D_5_reset = reset; // @[:@12753.4]
  assign Mem1D_5_io_r_ofs_0 = _T_995[9:0]; // @[MemPrimitives.scala 131:28:@13538.4]
  assign Mem1D_5_io_r_backpressure = _T_995[10]; // @[MemPrimitives.scala 132:32:@13539.4]
  assign Mem1D_5_io_w_ofs_0 = _T_377[9:0]; // @[MemPrimitives.scala 94:28:@12932.4]
  assign Mem1D_5_io_w_data_0 = _T_377[41:10]; // @[MemPrimitives.scala 95:29:@12933.4]
  assign Mem1D_5_io_w_en_0 = _T_377[42]; // @[MemPrimitives.scala 96:27:@12934.4]
  assign Mem1D_6_clock = clock; // @[:@12768.4]
  assign Mem1D_6_reset = reset; // @[:@12769.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1087[9:0]; // @[MemPrimitives.scala 131:28:@13627.4]
  assign Mem1D_6_io_r_backpressure = _T_1087[10]; // @[MemPrimitives.scala 132:32:@13628.4]
  assign Mem1D_6_io_w_ofs_0 = _T_388[9:0]; // @[MemPrimitives.scala 94:28:@12944.4]
  assign Mem1D_6_io_w_data_0 = _T_388[41:10]; // @[MemPrimitives.scala 95:29:@12945.4]
  assign Mem1D_6_io_w_en_0 = _T_388[42]; // @[MemPrimitives.scala 96:27:@12946.4]
  assign Mem1D_7_clock = clock; // @[:@12784.4]
  assign Mem1D_7_reset = reset; // @[:@12785.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1179[9:0]; // @[MemPrimitives.scala 131:28:@13716.4]
  assign Mem1D_7_io_r_backpressure = _T_1179[10]; // @[MemPrimitives.scala 132:32:@13717.4]
  assign Mem1D_7_io_w_ofs_0 = _T_399[9:0]; // @[MemPrimitives.scala 94:28:@12956.4]
  assign Mem1D_7_io_w_data_0 = _T_399[41:10]; // @[MemPrimitives.scala 95:29:@12957.4]
  assign Mem1D_7_io_w_en_0 = _T_399[42]; // @[MemPrimitives.scala 96:27:@12958.4]
  assign Mem1D_8_clock = clock; // @[:@12800.4]
  assign Mem1D_8_reset = reset; // @[:@12801.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1271[9:0]; // @[MemPrimitives.scala 131:28:@13805.4]
  assign Mem1D_8_io_r_backpressure = _T_1271[10]; // @[MemPrimitives.scala 132:32:@13806.4]
  assign Mem1D_8_io_w_ofs_0 = _T_410[9:0]; // @[MemPrimitives.scala 94:28:@12968.4]
  assign Mem1D_8_io_w_data_0 = _T_410[41:10]; // @[MemPrimitives.scala 95:29:@12969.4]
  assign Mem1D_8_io_w_en_0 = _T_410[42]; // @[MemPrimitives.scala 96:27:@12970.4]
  assign Mem1D_9_clock = clock; // @[:@12816.4]
  assign Mem1D_9_reset = reset; // @[:@12817.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1363[9:0]; // @[MemPrimitives.scala 131:28:@13894.4]
  assign Mem1D_9_io_r_backpressure = _T_1363[10]; // @[MemPrimitives.scala 132:32:@13895.4]
  assign Mem1D_9_io_w_ofs_0 = _T_421[9:0]; // @[MemPrimitives.scala 94:28:@12980.4]
  assign Mem1D_9_io_w_data_0 = _T_421[41:10]; // @[MemPrimitives.scala 95:29:@12981.4]
  assign Mem1D_9_io_w_en_0 = _T_421[42]; // @[MemPrimitives.scala 96:27:@12982.4]
  assign Mem1D_10_clock = clock; // @[:@12832.4]
  assign Mem1D_10_reset = reset; // @[:@12833.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1455[9:0]; // @[MemPrimitives.scala 131:28:@13983.4]
  assign Mem1D_10_io_r_backpressure = _T_1455[10]; // @[MemPrimitives.scala 132:32:@13984.4]
  assign Mem1D_10_io_w_ofs_0 = _T_432[9:0]; // @[MemPrimitives.scala 94:28:@12992.4]
  assign Mem1D_10_io_w_data_0 = _T_432[41:10]; // @[MemPrimitives.scala 95:29:@12993.4]
  assign Mem1D_10_io_w_en_0 = _T_432[42]; // @[MemPrimitives.scala 96:27:@12994.4]
  assign Mem1D_11_clock = clock; // @[:@12848.4]
  assign Mem1D_11_reset = reset; // @[:@12849.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1547[9:0]; // @[MemPrimitives.scala 131:28:@14072.4]
  assign Mem1D_11_io_r_backpressure = _T_1547[10]; // @[MemPrimitives.scala 132:32:@14073.4]
  assign Mem1D_11_io_w_ofs_0 = _T_443[9:0]; // @[MemPrimitives.scala 94:28:@13004.4]
  assign Mem1D_11_io_w_data_0 = _T_443[41:10]; // @[MemPrimitives.scala 95:29:@13005.4]
  assign Mem1D_11_io_w_en_0 = _T_443[42]; // @[MemPrimitives.scala 96:27:@13006.4]
  assign StickySelects_clock = clock; // @[:@13044.4]
  assign StickySelects_reset = reset; // @[:@13045.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_451; // @[MemPrimitives.scala 125:64:@13046.4]
  assign StickySelects_io_ins_1 = io_rPort_1_en_0 & _T_457; // @[MemPrimitives.scala 125:64:@13047.4]
  assign StickySelects_io_ins_2 = io_rPort_2_en_0 & _T_463; // @[MemPrimitives.scala 125:64:@13048.4]
  assign StickySelects_io_ins_3 = io_rPort_3_en_0 & _T_469; // @[MemPrimitives.scala 125:64:@13049.4]
  assign StickySelects_io_ins_4 = io_rPort_4_en_0 & _T_475; // @[MemPrimitives.scala 125:64:@13050.4]
  assign StickySelects_io_ins_5 = io_rPort_5_en_0 & _T_481; // @[MemPrimitives.scala 125:64:@13051.4]
  assign StickySelects_io_ins_6 = io_rPort_6_en_0 & _T_487; // @[MemPrimitives.scala 125:64:@13052.4]
  assign StickySelects_io_ins_7 = io_rPort_7_en_0 & _T_493; // @[MemPrimitives.scala 125:64:@13053.4]
  assign StickySelects_io_ins_8 = io_rPort_8_en_0 & _T_499; // @[MemPrimitives.scala 125:64:@13054.4]
  assign StickySelects_1_clock = clock; // @[:@13133.4]
  assign StickySelects_1_reset = reset; // @[:@13134.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_543; // @[MemPrimitives.scala 125:64:@13135.4]
  assign StickySelects_1_io_ins_1 = io_rPort_1_en_0 & _T_549; // @[MemPrimitives.scala 125:64:@13136.4]
  assign StickySelects_1_io_ins_2 = io_rPort_2_en_0 & _T_555; // @[MemPrimitives.scala 125:64:@13137.4]
  assign StickySelects_1_io_ins_3 = io_rPort_3_en_0 & _T_561; // @[MemPrimitives.scala 125:64:@13138.4]
  assign StickySelects_1_io_ins_4 = io_rPort_4_en_0 & _T_567; // @[MemPrimitives.scala 125:64:@13139.4]
  assign StickySelects_1_io_ins_5 = io_rPort_5_en_0 & _T_573; // @[MemPrimitives.scala 125:64:@13140.4]
  assign StickySelects_1_io_ins_6 = io_rPort_6_en_0 & _T_579; // @[MemPrimitives.scala 125:64:@13141.4]
  assign StickySelects_1_io_ins_7 = io_rPort_7_en_0 & _T_585; // @[MemPrimitives.scala 125:64:@13142.4]
  assign StickySelects_1_io_ins_8 = io_rPort_8_en_0 & _T_591; // @[MemPrimitives.scala 125:64:@13143.4]
  assign StickySelects_2_clock = clock; // @[:@13222.4]
  assign StickySelects_2_reset = reset; // @[:@13223.4]
  assign StickySelects_2_io_ins_0 = io_rPort_0_en_0 & _T_635; // @[MemPrimitives.scala 125:64:@13224.4]
  assign StickySelects_2_io_ins_1 = io_rPort_1_en_0 & _T_641; // @[MemPrimitives.scala 125:64:@13225.4]
  assign StickySelects_2_io_ins_2 = io_rPort_2_en_0 & _T_647; // @[MemPrimitives.scala 125:64:@13226.4]
  assign StickySelects_2_io_ins_3 = io_rPort_3_en_0 & _T_653; // @[MemPrimitives.scala 125:64:@13227.4]
  assign StickySelects_2_io_ins_4 = io_rPort_4_en_0 & _T_659; // @[MemPrimitives.scala 125:64:@13228.4]
  assign StickySelects_2_io_ins_5 = io_rPort_5_en_0 & _T_665; // @[MemPrimitives.scala 125:64:@13229.4]
  assign StickySelects_2_io_ins_6 = io_rPort_6_en_0 & _T_671; // @[MemPrimitives.scala 125:64:@13230.4]
  assign StickySelects_2_io_ins_7 = io_rPort_7_en_0 & _T_677; // @[MemPrimitives.scala 125:64:@13231.4]
  assign StickySelects_2_io_ins_8 = io_rPort_8_en_0 & _T_683; // @[MemPrimitives.scala 125:64:@13232.4]
  assign StickySelects_3_clock = clock; // @[:@13311.4]
  assign StickySelects_3_reset = reset; // @[:@13312.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_727; // @[MemPrimitives.scala 125:64:@13313.4]
  assign StickySelects_3_io_ins_1 = io_rPort_1_en_0 & _T_733; // @[MemPrimitives.scala 125:64:@13314.4]
  assign StickySelects_3_io_ins_2 = io_rPort_2_en_0 & _T_739; // @[MemPrimitives.scala 125:64:@13315.4]
  assign StickySelects_3_io_ins_3 = io_rPort_3_en_0 & _T_745; // @[MemPrimitives.scala 125:64:@13316.4]
  assign StickySelects_3_io_ins_4 = io_rPort_4_en_0 & _T_751; // @[MemPrimitives.scala 125:64:@13317.4]
  assign StickySelects_3_io_ins_5 = io_rPort_5_en_0 & _T_757; // @[MemPrimitives.scala 125:64:@13318.4]
  assign StickySelects_3_io_ins_6 = io_rPort_6_en_0 & _T_763; // @[MemPrimitives.scala 125:64:@13319.4]
  assign StickySelects_3_io_ins_7 = io_rPort_7_en_0 & _T_769; // @[MemPrimitives.scala 125:64:@13320.4]
  assign StickySelects_3_io_ins_8 = io_rPort_8_en_0 & _T_775; // @[MemPrimitives.scala 125:64:@13321.4]
  assign StickySelects_4_clock = clock; // @[:@13400.4]
  assign StickySelects_4_reset = reset; // @[:@13401.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_819; // @[MemPrimitives.scala 125:64:@13402.4]
  assign StickySelects_4_io_ins_1 = io_rPort_1_en_0 & _T_825; // @[MemPrimitives.scala 125:64:@13403.4]
  assign StickySelects_4_io_ins_2 = io_rPort_2_en_0 & _T_831; // @[MemPrimitives.scala 125:64:@13404.4]
  assign StickySelects_4_io_ins_3 = io_rPort_3_en_0 & _T_837; // @[MemPrimitives.scala 125:64:@13405.4]
  assign StickySelects_4_io_ins_4 = io_rPort_4_en_0 & _T_843; // @[MemPrimitives.scala 125:64:@13406.4]
  assign StickySelects_4_io_ins_5 = io_rPort_5_en_0 & _T_849; // @[MemPrimitives.scala 125:64:@13407.4]
  assign StickySelects_4_io_ins_6 = io_rPort_6_en_0 & _T_855; // @[MemPrimitives.scala 125:64:@13408.4]
  assign StickySelects_4_io_ins_7 = io_rPort_7_en_0 & _T_861; // @[MemPrimitives.scala 125:64:@13409.4]
  assign StickySelects_4_io_ins_8 = io_rPort_8_en_0 & _T_867; // @[MemPrimitives.scala 125:64:@13410.4]
  assign StickySelects_5_clock = clock; // @[:@13489.4]
  assign StickySelects_5_reset = reset; // @[:@13490.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_911; // @[MemPrimitives.scala 125:64:@13491.4]
  assign StickySelects_5_io_ins_1 = io_rPort_1_en_0 & _T_917; // @[MemPrimitives.scala 125:64:@13492.4]
  assign StickySelects_5_io_ins_2 = io_rPort_2_en_0 & _T_923; // @[MemPrimitives.scala 125:64:@13493.4]
  assign StickySelects_5_io_ins_3 = io_rPort_3_en_0 & _T_929; // @[MemPrimitives.scala 125:64:@13494.4]
  assign StickySelects_5_io_ins_4 = io_rPort_4_en_0 & _T_935; // @[MemPrimitives.scala 125:64:@13495.4]
  assign StickySelects_5_io_ins_5 = io_rPort_5_en_0 & _T_941; // @[MemPrimitives.scala 125:64:@13496.4]
  assign StickySelects_5_io_ins_6 = io_rPort_6_en_0 & _T_947; // @[MemPrimitives.scala 125:64:@13497.4]
  assign StickySelects_5_io_ins_7 = io_rPort_7_en_0 & _T_953; // @[MemPrimitives.scala 125:64:@13498.4]
  assign StickySelects_5_io_ins_8 = io_rPort_8_en_0 & _T_959; // @[MemPrimitives.scala 125:64:@13499.4]
  assign StickySelects_6_clock = clock; // @[:@13578.4]
  assign StickySelects_6_reset = reset; // @[:@13579.4]
  assign StickySelects_6_io_ins_0 = io_rPort_0_en_0 & _T_1003; // @[MemPrimitives.scala 125:64:@13580.4]
  assign StickySelects_6_io_ins_1 = io_rPort_1_en_0 & _T_1009; // @[MemPrimitives.scala 125:64:@13581.4]
  assign StickySelects_6_io_ins_2 = io_rPort_2_en_0 & _T_1015; // @[MemPrimitives.scala 125:64:@13582.4]
  assign StickySelects_6_io_ins_3 = io_rPort_3_en_0 & _T_1021; // @[MemPrimitives.scala 125:64:@13583.4]
  assign StickySelects_6_io_ins_4 = io_rPort_4_en_0 & _T_1027; // @[MemPrimitives.scala 125:64:@13584.4]
  assign StickySelects_6_io_ins_5 = io_rPort_5_en_0 & _T_1033; // @[MemPrimitives.scala 125:64:@13585.4]
  assign StickySelects_6_io_ins_6 = io_rPort_6_en_0 & _T_1039; // @[MemPrimitives.scala 125:64:@13586.4]
  assign StickySelects_6_io_ins_7 = io_rPort_7_en_0 & _T_1045; // @[MemPrimitives.scala 125:64:@13587.4]
  assign StickySelects_6_io_ins_8 = io_rPort_8_en_0 & _T_1051; // @[MemPrimitives.scala 125:64:@13588.4]
  assign StickySelects_7_clock = clock; // @[:@13667.4]
  assign StickySelects_7_reset = reset; // @[:@13668.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_1095; // @[MemPrimitives.scala 125:64:@13669.4]
  assign StickySelects_7_io_ins_1 = io_rPort_1_en_0 & _T_1101; // @[MemPrimitives.scala 125:64:@13670.4]
  assign StickySelects_7_io_ins_2 = io_rPort_2_en_0 & _T_1107; // @[MemPrimitives.scala 125:64:@13671.4]
  assign StickySelects_7_io_ins_3 = io_rPort_3_en_0 & _T_1113; // @[MemPrimitives.scala 125:64:@13672.4]
  assign StickySelects_7_io_ins_4 = io_rPort_4_en_0 & _T_1119; // @[MemPrimitives.scala 125:64:@13673.4]
  assign StickySelects_7_io_ins_5 = io_rPort_5_en_0 & _T_1125; // @[MemPrimitives.scala 125:64:@13674.4]
  assign StickySelects_7_io_ins_6 = io_rPort_6_en_0 & _T_1131; // @[MemPrimitives.scala 125:64:@13675.4]
  assign StickySelects_7_io_ins_7 = io_rPort_7_en_0 & _T_1137; // @[MemPrimitives.scala 125:64:@13676.4]
  assign StickySelects_7_io_ins_8 = io_rPort_8_en_0 & _T_1143; // @[MemPrimitives.scala 125:64:@13677.4]
  assign StickySelects_8_clock = clock; // @[:@13756.4]
  assign StickySelects_8_reset = reset; // @[:@13757.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_1187; // @[MemPrimitives.scala 125:64:@13758.4]
  assign StickySelects_8_io_ins_1 = io_rPort_1_en_0 & _T_1193; // @[MemPrimitives.scala 125:64:@13759.4]
  assign StickySelects_8_io_ins_2 = io_rPort_2_en_0 & _T_1199; // @[MemPrimitives.scala 125:64:@13760.4]
  assign StickySelects_8_io_ins_3 = io_rPort_3_en_0 & _T_1205; // @[MemPrimitives.scala 125:64:@13761.4]
  assign StickySelects_8_io_ins_4 = io_rPort_4_en_0 & _T_1211; // @[MemPrimitives.scala 125:64:@13762.4]
  assign StickySelects_8_io_ins_5 = io_rPort_5_en_0 & _T_1217; // @[MemPrimitives.scala 125:64:@13763.4]
  assign StickySelects_8_io_ins_6 = io_rPort_6_en_0 & _T_1223; // @[MemPrimitives.scala 125:64:@13764.4]
  assign StickySelects_8_io_ins_7 = io_rPort_7_en_0 & _T_1229; // @[MemPrimitives.scala 125:64:@13765.4]
  assign StickySelects_8_io_ins_8 = io_rPort_8_en_0 & _T_1235; // @[MemPrimitives.scala 125:64:@13766.4]
  assign StickySelects_9_clock = clock; // @[:@13845.4]
  assign StickySelects_9_reset = reset; // @[:@13846.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_1279; // @[MemPrimitives.scala 125:64:@13847.4]
  assign StickySelects_9_io_ins_1 = io_rPort_1_en_0 & _T_1285; // @[MemPrimitives.scala 125:64:@13848.4]
  assign StickySelects_9_io_ins_2 = io_rPort_2_en_0 & _T_1291; // @[MemPrimitives.scala 125:64:@13849.4]
  assign StickySelects_9_io_ins_3 = io_rPort_3_en_0 & _T_1297; // @[MemPrimitives.scala 125:64:@13850.4]
  assign StickySelects_9_io_ins_4 = io_rPort_4_en_0 & _T_1303; // @[MemPrimitives.scala 125:64:@13851.4]
  assign StickySelects_9_io_ins_5 = io_rPort_5_en_0 & _T_1309; // @[MemPrimitives.scala 125:64:@13852.4]
  assign StickySelects_9_io_ins_6 = io_rPort_6_en_0 & _T_1315; // @[MemPrimitives.scala 125:64:@13853.4]
  assign StickySelects_9_io_ins_7 = io_rPort_7_en_0 & _T_1321; // @[MemPrimitives.scala 125:64:@13854.4]
  assign StickySelects_9_io_ins_8 = io_rPort_8_en_0 & _T_1327; // @[MemPrimitives.scala 125:64:@13855.4]
  assign StickySelects_10_clock = clock; // @[:@13934.4]
  assign StickySelects_10_reset = reset; // @[:@13935.4]
  assign StickySelects_10_io_ins_0 = io_rPort_0_en_0 & _T_1371; // @[MemPrimitives.scala 125:64:@13936.4]
  assign StickySelects_10_io_ins_1 = io_rPort_1_en_0 & _T_1377; // @[MemPrimitives.scala 125:64:@13937.4]
  assign StickySelects_10_io_ins_2 = io_rPort_2_en_0 & _T_1383; // @[MemPrimitives.scala 125:64:@13938.4]
  assign StickySelects_10_io_ins_3 = io_rPort_3_en_0 & _T_1389; // @[MemPrimitives.scala 125:64:@13939.4]
  assign StickySelects_10_io_ins_4 = io_rPort_4_en_0 & _T_1395; // @[MemPrimitives.scala 125:64:@13940.4]
  assign StickySelects_10_io_ins_5 = io_rPort_5_en_0 & _T_1401; // @[MemPrimitives.scala 125:64:@13941.4]
  assign StickySelects_10_io_ins_6 = io_rPort_6_en_0 & _T_1407; // @[MemPrimitives.scala 125:64:@13942.4]
  assign StickySelects_10_io_ins_7 = io_rPort_7_en_0 & _T_1413; // @[MemPrimitives.scala 125:64:@13943.4]
  assign StickySelects_10_io_ins_8 = io_rPort_8_en_0 & _T_1419; // @[MemPrimitives.scala 125:64:@13944.4]
  assign StickySelects_11_clock = clock; // @[:@14023.4]
  assign StickySelects_11_reset = reset; // @[:@14024.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_1463; // @[MemPrimitives.scala 125:64:@14025.4]
  assign StickySelects_11_io_ins_1 = io_rPort_1_en_0 & _T_1469; // @[MemPrimitives.scala 125:64:@14026.4]
  assign StickySelects_11_io_ins_2 = io_rPort_2_en_0 & _T_1475; // @[MemPrimitives.scala 125:64:@14027.4]
  assign StickySelects_11_io_ins_3 = io_rPort_3_en_0 & _T_1481; // @[MemPrimitives.scala 125:64:@14028.4]
  assign StickySelects_11_io_ins_4 = io_rPort_4_en_0 & _T_1487; // @[MemPrimitives.scala 125:64:@14029.4]
  assign StickySelects_11_io_ins_5 = io_rPort_5_en_0 & _T_1493; // @[MemPrimitives.scala 125:64:@14030.4]
  assign StickySelects_11_io_ins_6 = io_rPort_6_en_0 & _T_1499; // @[MemPrimitives.scala 125:64:@14031.4]
  assign StickySelects_11_io_ins_7 = io_rPort_7_en_0 & _T_1505; // @[MemPrimitives.scala 125:64:@14032.4]
  assign StickySelects_11_io_ins_8 = io_rPort_8_en_0 & _T_1511; // @[MemPrimitives.scala 125:64:@14033.4]
  assign RetimeWrapper_clock = clock; // @[:@14113.4]
  assign RetimeWrapper_reset = reset; // @[:@14114.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14116.4]
  assign RetimeWrapper_io_in = _T_451 & io_rPort_0_en_0; // @[package.scala 94:16:@14115.4]
  assign RetimeWrapper_1_clock = clock; // @[:@14121.4]
  assign RetimeWrapper_1_reset = reset; // @[:@14122.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14124.4]
  assign RetimeWrapper_1_io_in = _T_543 & io_rPort_0_en_0; // @[package.scala 94:16:@14123.4]
  assign RetimeWrapper_2_clock = clock; // @[:@14129.4]
  assign RetimeWrapper_2_reset = reset; // @[:@14130.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14132.4]
  assign RetimeWrapper_2_io_in = _T_635 & io_rPort_0_en_0; // @[package.scala 94:16:@14131.4]
  assign RetimeWrapper_3_clock = clock; // @[:@14137.4]
  assign RetimeWrapper_3_reset = reset; // @[:@14138.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14140.4]
  assign RetimeWrapper_3_io_in = _T_727 & io_rPort_0_en_0; // @[package.scala 94:16:@14139.4]
  assign RetimeWrapper_4_clock = clock; // @[:@14145.4]
  assign RetimeWrapper_4_reset = reset; // @[:@14146.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14148.4]
  assign RetimeWrapper_4_io_in = _T_819 & io_rPort_0_en_0; // @[package.scala 94:16:@14147.4]
  assign RetimeWrapper_5_clock = clock; // @[:@14153.4]
  assign RetimeWrapper_5_reset = reset; // @[:@14154.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14156.4]
  assign RetimeWrapper_5_io_in = _T_911 & io_rPort_0_en_0; // @[package.scala 94:16:@14155.4]
  assign RetimeWrapper_6_clock = clock; // @[:@14161.4]
  assign RetimeWrapper_6_reset = reset; // @[:@14162.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14164.4]
  assign RetimeWrapper_6_io_in = _T_1003 & io_rPort_0_en_0; // @[package.scala 94:16:@14163.4]
  assign RetimeWrapper_7_clock = clock; // @[:@14169.4]
  assign RetimeWrapper_7_reset = reset; // @[:@14170.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14172.4]
  assign RetimeWrapper_7_io_in = _T_1095 & io_rPort_0_en_0; // @[package.scala 94:16:@14171.4]
  assign RetimeWrapper_8_clock = clock; // @[:@14177.4]
  assign RetimeWrapper_8_reset = reset; // @[:@14178.4]
  assign RetimeWrapper_8_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14180.4]
  assign RetimeWrapper_8_io_in = _T_1187 & io_rPort_0_en_0; // @[package.scala 94:16:@14179.4]
  assign RetimeWrapper_9_clock = clock; // @[:@14185.4]
  assign RetimeWrapper_9_reset = reset; // @[:@14186.4]
  assign RetimeWrapper_9_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14188.4]
  assign RetimeWrapper_9_io_in = _T_1279 & io_rPort_0_en_0; // @[package.scala 94:16:@14187.4]
  assign RetimeWrapper_10_clock = clock; // @[:@14193.4]
  assign RetimeWrapper_10_reset = reset; // @[:@14194.4]
  assign RetimeWrapper_10_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14196.4]
  assign RetimeWrapper_10_io_in = _T_1371 & io_rPort_0_en_0; // @[package.scala 94:16:@14195.4]
  assign RetimeWrapper_11_clock = clock; // @[:@14201.4]
  assign RetimeWrapper_11_reset = reset; // @[:@14202.4]
  assign RetimeWrapper_11_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14204.4]
  assign RetimeWrapper_11_io_in = _T_1463 & io_rPort_0_en_0; // @[package.scala 94:16:@14203.4]
  assign RetimeWrapper_12_clock = clock; // @[:@14257.4]
  assign RetimeWrapper_12_reset = reset; // @[:@14258.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14260.4]
  assign RetimeWrapper_12_io_in = _T_457 & io_rPort_1_en_0; // @[package.scala 94:16:@14259.4]
  assign RetimeWrapper_13_clock = clock; // @[:@14265.4]
  assign RetimeWrapper_13_reset = reset; // @[:@14266.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14268.4]
  assign RetimeWrapper_13_io_in = _T_549 & io_rPort_1_en_0; // @[package.scala 94:16:@14267.4]
  assign RetimeWrapper_14_clock = clock; // @[:@14273.4]
  assign RetimeWrapper_14_reset = reset; // @[:@14274.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14276.4]
  assign RetimeWrapper_14_io_in = _T_641 & io_rPort_1_en_0; // @[package.scala 94:16:@14275.4]
  assign RetimeWrapper_15_clock = clock; // @[:@14281.4]
  assign RetimeWrapper_15_reset = reset; // @[:@14282.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14284.4]
  assign RetimeWrapper_15_io_in = _T_733 & io_rPort_1_en_0; // @[package.scala 94:16:@14283.4]
  assign RetimeWrapper_16_clock = clock; // @[:@14289.4]
  assign RetimeWrapper_16_reset = reset; // @[:@14290.4]
  assign RetimeWrapper_16_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14292.4]
  assign RetimeWrapper_16_io_in = _T_825 & io_rPort_1_en_0; // @[package.scala 94:16:@14291.4]
  assign RetimeWrapper_17_clock = clock; // @[:@14297.4]
  assign RetimeWrapper_17_reset = reset; // @[:@14298.4]
  assign RetimeWrapper_17_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14300.4]
  assign RetimeWrapper_17_io_in = _T_917 & io_rPort_1_en_0; // @[package.scala 94:16:@14299.4]
  assign RetimeWrapper_18_clock = clock; // @[:@14305.4]
  assign RetimeWrapper_18_reset = reset; // @[:@14306.4]
  assign RetimeWrapper_18_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14308.4]
  assign RetimeWrapper_18_io_in = _T_1009 & io_rPort_1_en_0; // @[package.scala 94:16:@14307.4]
  assign RetimeWrapper_19_clock = clock; // @[:@14313.4]
  assign RetimeWrapper_19_reset = reset; // @[:@14314.4]
  assign RetimeWrapper_19_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14316.4]
  assign RetimeWrapper_19_io_in = _T_1101 & io_rPort_1_en_0; // @[package.scala 94:16:@14315.4]
  assign RetimeWrapper_20_clock = clock; // @[:@14321.4]
  assign RetimeWrapper_20_reset = reset; // @[:@14322.4]
  assign RetimeWrapper_20_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14324.4]
  assign RetimeWrapper_20_io_in = _T_1193 & io_rPort_1_en_0; // @[package.scala 94:16:@14323.4]
  assign RetimeWrapper_21_clock = clock; // @[:@14329.4]
  assign RetimeWrapper_21_reset = reset; // @[:@14330.4]
  assign RetimeWrapper_21_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14332.4]
  assign RetimeWrapper_21_io_in = _T_1285 & io_rPort_1_en_0; // @[package.scala 94:16:@14331.4]
  assign RetimeWrapper_22_clock = clock; // @[:@14337.4]
  assign RetimeWrapper_22_reset = reset; // @[:@14338.4]
  assign RetimeWrapper_22_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14340.4]
  assign RetimeWrapper_22_io_in = _T_1377 & io_rPort_1_en_0; // @[package.scala 94:16:@14339.4]
  assign RetimeWrapper_23_clock = clock; // @[:@14345.4]
  assign RetimeWrapper_23_reset = reset; // @[:@14346.4]
  assign RetimeWrapper_23_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14348.4]
  assign RetimeWrapper_23_io_in = _T_1469 & io_rPort_1_en_0; // @[package.scala 94:16:@14347.4]
  assign RetimeWrapper_24_clock = clock; // @[:@14401.4]
  assign RetimeWrapper_24_reset = reset; // @[:@14402.4]
  assign RetimeWrapper_24_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14404.4]
  assign RetimeWrapper_24_io_in = _T_463 & io_rPort_2_en_0; // @[package.scala 94:16:@14403.4]
  assign RetimeWrapper_25_clock = clock; // @[:@14409.4]
  assign RetimeWrapper_25_reset = reset; // @[:@14410.4]
  assign RetimeWrapper_25_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14412.4]
  assign RetimeWrapper_25_io_in = _T_555 & io_rPort_2_en_0; // @[package.scala 94:16:@14411.4]
  assign RetimeWrapper_26_clock = clock; // @[:@14417.4]
  assign RetimeWrapper_26_reset = reset; // @[:@14418.4]
  assign RetimeWrapper_26_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14420.4]
  assign RetimeWrapper_26_io_in = _T_647 & io_rPort_2_en_0; // @[package.scala 94:16:@14419.4]
  assign RetimeWrapper_27_clock = clock; // @[:@14425.4]
  assign RetimeWrapper_27_reset = reset; // @[:@14426.4]
  assign RetimeWrapper_27_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14428.4]
  assign RetimeWrapper_27_io_in = _T_739 & io_rPort_2_en_0; // @[package.scala 94:16:@14427.4]
  assign RetimeWrapper_28_clock = clock; // @[:@14433.4]
  assign RetimeWrapper_28_reset = reset; // @[:@14434.4]
  assign RetimeWrapper_28_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14436.4]
  assign RetimeWrapper_28_io_in = _T_831 & io_rPort_2_en_0; // @[package.scala 94:16:@14435.4]
  assign RetimeWrapper_29_clock = clock; // @[:@14441.4]
  assign RetimeWrapper_29_reset = reset; // @[:@14442.4]
  assign RetimeWrapper_29_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14444.4]
  assign RetimeWrapper_29_io_in = _T_923 & io_rPort_2_en_0; // @[package.scala 94:16:@14443.4]
  assign RetimeWrapper_30_clock = clock; // @[:@14449.4]
  assign RetimeWrapper_30_reset = reset; // @[:@14450.4]
  assign RetimeWrapper_30_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14452.4]
  assign RetimeWrapper_30_io_in = _T_1015 & io_rPort_2_en_0; // @[package.scala 94:16:@14451.4]
  assign RetimeWrapper_31_clock = clock; // @[:@14457.4]
  assign RetimeWrapper_31_reset = reset; // @[:@14458.4]
  assign RetimeWrapper_31_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14460.4]
  assign RetimeWrapper_31_io_in = _T_1107 & io_rPort_2_en_0; // @[package.scala 94:16:@14459.4]
  assign RetimeWrapper_32_clock = clock; // @[:@14465.4]
  assign RetimeWrapper_32_reset = reset; // @[:@14466.4]
  assign RetimeWrapper_32_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14468.4]
  assign RetimeWrapper_32_io_in = _T_1199 & io_rPort_2_en_0; // @[package.scala 94:16:@14467.4]
  assign RetimeWrapper_33_clock = clock; // @[:@14473.4]
  assign RetimeWrapper_33_reset = reset; // @[:@14474.4]
  assign RetimeWrapper_33_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14476.4]
  assign RetimeWrapper_33_io_in = _T_1291 & io_rPort_2_en_0; // @[package.scala 94:16:@14475.4]
  assign RetimeWrapper_34_clock = clock; // @[:@14481.4]
  assign RetimeWrapper_34_reset = reset; // @[:@14482.4]
  assign RetimeWrapper_34_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14484.4]
  assign RetimeWrapper_34_io_in = _T_1383 & io_rPort_2_en_0; // @[package.scala 94:16:@14483.4]
  assign RetimeWrapper_35_clock = clock; // @[:@14489.4]
  assign RetimeWrapper_35_reset = reset; // @[:@14490.4]
  assign RetimeWrapper_35_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14492.4]
  assign RetimeWrapper_35_io_in = _T_1475 & io_rPort_2_en_0; // @[package.scala 94:16:@14491.4]
  assign RetimeWrapper_36_clock = clock; // @[:@14545.4]
  assign RetimeWrapper_36_reset = reset; // @[:@14546.4]
  assign RetimeWrapper_36_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14548.4]
  assign RetimeWrapper_36_io_in = _T_469 & io_rPort_3_en_0; // @[package.scala 94:16:@14547.4]
  assign RetimeWrapper_37_clock = clock; // @[:@14553.4]
  assign RetimeWrapper_37_reset = reset; // @[:@14554.4]
  assign RetimeWrapper_37_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14556.4]
  assign RetimeWrapper_37_io_in = _T_561 & io_rPort_3_en_0; // @[package.scala 94:16:@14555.4]
  assign RetimeWrapper_38_clock = clock; // @[:@14561.4]
  assign RetimeWrapper_38_reset = reset; // @[:@14562.4]
  assign RetimeWrapper_38_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14564.4]
  assign RetimeWrapper_38_io_in = _T_653 & io_rPort_3_en_0; // @[package.scala 94:16:@14563.4]
  assign RetimeWrapper_39_clock = clock; // @[:@14569.4]
  assign RetimeWrapper_39_reset = reset; // @[:@14570.4]
  assign RetimeWrapper_39_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14572.4]
  assign RetimeWrapper_39_io_in = _T_745 & io_rPort_3_en_0; // @[package.scala 94:16:@14571.4]
  assign RetimeWrapper_40_clock = clock; // @[:@14577.4]
  assign RetimeWrapper_40_reset = reset; // @[:@14578.4]
  assign RetimeWrapper_40_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14580.4]
  assign RetimeWrapper_40_io_in = _T_837 & io_rPort_3_en_0; // @[package.scala 94:16:@14579.4]
  assign RetimeWrapper_41_clock = clock; // @[:@14585.4]
  assign RetimeWrapper_41_reset = reset; // @[:@14586.4]
  assign RetimeWrapper_41_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14588.4]
  assign RetimeWrapper_41_io_in = _T_929 & io_rPort_3_en_0; // @[package.scala 94:16:@14587.4]
  assign RetimeWrapper_42_clock = clock; // @[:@14593.4]
  assign RetimeWrapper_42_reset = reset; // @[:@14594.4]
  assign RetimeWrapper_42_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14596.4]
  assign RetimeWrapper_42_io_in = _T_1021 & io_rPort_3_en_0; // @[package.scala 94:16:@14595.4]
  assign RetimeWrapper_43_clock = clock; // @[:@14601.4]
  assign RetimeWrapper_43_reset = reset; // @[:@14602.4]
  assign RetimeWrapper_43_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14604.4]
  assign RetimeWrapper_43_io_in = _T_1113 & io_rPort_3_en_0; // @[package.scala 94:16:@14603.4]
  assign RetimeWrapper_44_clock = clock; // @[:@14609.4]
  assign RetimeWrapper_44_reset = reset; // @[:@14610.4]
  assign RetimeWrapper_44_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14612.4]
  assign RetimeWrapper_44_io_in = _T_1205 & io_rPort_3_en_0; // @[package.scala 94:16:@14611.4]
  assign RetimeWrapper_45_clock = clock; // @[:@14617.4]
  assign RetimeWrapper_45_reset = reset; // @[:@14618.4]
  assign RetimeWrapper_45_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14620.4]
  assign RetimeWrapper_45_io_in = _T_1297 & io_rPort_3_en_0; // @[package.scala 94:16:@14619.4]
  assign RetimeWrapper_46_clock = clock; // @[:@14625.4]
  assign RetimeWrapper_46_reset = reset; // @[:@14626.4]
  assign RetimeWrapper_46_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14628.4]
  assign RetimeWrapper_46_io_in = _T_1389 & io_rPort_3_en_0; // @[package.scala 94:16:@14627.4]
  assign RetimeWrapper_47_clock = clock; // @[:@14633.4]
  assign RetimeWrapper_47_reset = reset; // @[:@14634.4]
  assign RetimeWrapper_47_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14636.4]
  assign RetimeWrapper_47_io_in = _T_1481 & io_rPort_3_en_0; // @[package.scala 94:16:@14635.4]
  assign RetimeWrapper_48_clock = clock; // @[:@14689.4]
  assign RetimeWrapper_48_reset = reset; // @[:@14690.4]
  assign RetimeWrapper_48_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14692.4]
  assign RetimeWrapper_48_io_in = _T_475 & io_rPort_4_en_0; // @[package.scala 94:16:@14691.4]
  assign RetimeWrapper_49_clock = clock; // @[:@14697.4]
  assign RetimeWrapper_49_reset = reset; // @[:@14698.4]
  assign RetimeWrapper_49_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14700.4]
  assign RetimeWrapper_49_io_in = _T_567 & io_rPort_4_en_0; // @[package.scala 94:16:@14699.4]
  assign RetimeWrapper_50_clock = clock; // @[:@14705.4]
  assign RetimeWrapper_50_reset = reset; // @[:@14706.4]
  assign RetimeWrapper_50_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14708.4]
  assign RetimeWrapper_50_io_in = _T_659 & io_rPort_4_en_0; // @[package.scala 94:16:@14707.4]
  assign RetimeWrapper_51_clock = clock; // @[:@14713.4]
  assign RetimeWrapper_51_reset = reset; // @[:@14714.4]
  assign RetimeWrapper_51_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14716.4]
  assign RetimeWrapper_51_io_in = _T_751 & io_rPort_4_en_0; // @[package.scala 94:16:@14715.4]
  assign RetimeWrapper_52_clock = clock; // @[:@14721.4]
  assign RetimeWrapper_52_reset = reset; // @[:@14722.4]
  assign RetimeWrapper_52_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14724.4]
  assign RetimeWrapper_52_io_in = _T_843 & io_rPort_4_en_0; // @[package.scala 94:16:@14723.4]
  assign RetimeWrapper_53_clock = clock; // @[:@14729.4]
  assign RetimeWrapper_53_reset = reset; // @[:@14730.4]
  assign RetimeWrapper_53_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14732.4]
  assign RetimeWrapper_53_io_in = _T_935 & io_rPort_4_en_0; // @[package.scala 94:16:@14731.4]
  assign RetimeWrapper_54_clock = clock; // @[:@14737.4]
  assign RetimeWrapper_54_reset = reset; // @[:@14738.4]
  assign RetimeWrapper_54_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14740.4]
  assign RetimeWrapper_54_io_in = _T_1027 & io_rPort_4_en_0; // @[package.scala 94:16:@14739.4]
  assign RetimeWrapper_55_clock = clock; // @[:@14745.4]
  assign RetimeWrapper_55_reset = reset; // @[:@14746.4]
  assign RetimeWrapper_55_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14748.4]
  assign RetimeWrapper_55_io_in = _T_1119 & io_rPort_4_en_0; // @[package.scala 94:16:@14747.4]
  assign RetimeWrapper_56_clock = clock; // @[:@14753.4]
  assign RetimeWrapper_56_reset = reset; // @[:@14754.4]
  assign RetimeWrapper_56_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14756.4]
  assign RetimeWrapper_56_io_in = _T_1211 & io_rPort_4_en_0; // @[package.scala 94:16:@14755.4]
  assign RetimeWrapper_57_clock = clock; // @[:@14761.4]
  assign RetimeWrapper_57_reset = reset; // @[:@14762.4]
  assign RetimeWrapper_57_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14764.4]
  assign RetimeWrapper_57_io_in = _T_1303 & io_rPort_4_en_0; // @[package.scala 94:16:@14763.4]
  assign RetimeWrapper_58_clock = clock; // @[:@14769.4]
  assign RetimeWrapper_58_reset = reset; // @[:@14770.4]
  assign RetimeWrapper_58_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14772.4]
  assign RetimeWrapper_58_io_in = _T_1395 & io_rPort_4_en_0; // @[package.scala 94:16:@14771.4]
  assign RetimeWrapper_59_clock = clock; // @[:@14777.4]
  assign RetimeWrapper_59_reset = reset; // @[:@14778.4]
  assign RetimeWrapper_59_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14780.4]
  assign RetimeWrapper_59_io_in = _T_1487 & io_rPort_4_en_0; // @[package.scala 94:16:@14779.4]
  assign RetimeWrapper_60_clock = clock; // @[:@14833.4]
  assign RetimeWrapper_60_reset = reset; // @[:@14834.4]
  assign RetimeWrapper_60_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14836.4]
  assign RetimeWrapper_60_io_in = _T_481 & io_rPort_5_en_0; // @[package.scala 94:16:@14835.4]
  assign RetimeWrapper_61_clock = clock; // @[:@14841.4]
  assign RetimeWrapper_61_reset = reset; // @[:@14842.4]
  assign RetimeWrapper_61_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14844.4]
  assign RetimeWrapper_61_io_in = _T_573 & io_rPort_5_en_0; // @[package.scala 94:16:@14843.4]
  assign RetimeWrapper_62_clock = clock; // @[:@14849.4]
  assign RetimeWrapper_62_reset = reset; // @[:@14850.4]
  assign RetimeWrapper_62_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14852.4]
  assign RetimeWrapper_62_io_in = _T_665 & io_rPort_5_en_0; // @[package.scala 94:16:@14851.4]
  assign RetimeWrapper_63_clock = clock; // @[:@14857.4]
  assign RetimeWrapper_63_reset = reset; // @[:@14858.4]
  assign RetimeWrapper_63_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14860.4]
  assign RetimeWrapper_63_io_in = _T_757 & io_rPort_5_en_0; // @[package.scala 94:16:@14859.4]
  assign RetimeWrapper_64_clock = clock; // @[:@14865.4]
  assign RetimeWrapper_64_reset = reset; // @[:@14866.4]
  assign RetimeWrapper_64_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14868.4]
  assign RetimeWrapper_64_io_in = _T_849 & io_rPort_5_en_0; // @[package.scala 94:16:@14867.4]
  assign RetimeWrapper_65_clock = clock; // @[:@14873.4]
  assign RetimeWrapper_65_reset = reset; // @[:@14874.4]
  assign RetimeWrapper_65_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14876.4]
  assign RetimeWrapper_65_io_in = _T_941 & io_rPort_5_en_0; // @[package.scala 94:16:@14875.4]
  assign RetimeWrapper_66_clock = clock; // @[:@14881.4]
  assign RetimeWrapper_66_reset = reset; // @[:@14882.4]
  assign RetimeWrapper_66_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14884.4]
  assign RetimeWrapper_66_io_in = _T_1033 & io_rPort_5_en_0; // @[package.scala 94:16:@14883.4]
  assign RetimeWrapper_67_clock = clock; // @[:@14889.4]
  assign RetimeWrapper_67_reset = reset; // @[:@14890.4]
  assign RetimeWrapper_67_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14892.4]
  assign RetimeWrapper_67_io_in = _T_1125 & io_rPort_5_en_0; // @[package.scala 94:16:@14891.4]
  assign RetimeWrapper_68_clock = clock; // @[:@14897.4]
  assign RetimeWrapper_68_reset = reset; // @[:@14898.4]
  assign RetimeWrapper_68_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14900.4]
  assign RetimeWrapper_68_io_in = _T_1217 & io_rPort_5_en_0; // @[package.scala 94:16:@14899.4]
  assign RetimeWrapper_69_clock = clock; // @[:@14905.4]
  assign RetimeWrapper_69_reset = reset; // @[:@14906.4]
  assign RetimeWrapper_69_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14908.4]
  assign RetimeWrapper_69_io_in = _T_1309 & io_rPort_5_en_0; // @[package.scala 94:16:@14907.4]
  assign RetimeWrapper_70_clock = clock; // @[:@14913.4]
  assign RetimeWrapper_70_reset = reset; // @[:@14914.4]
  assign RetimeWrapper_70_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14916.4]
  assign RetimeWrapper_70_io_in = _T_1401 & io_rPort_5_en_0; // @[package.scala 94:16:@14915.4]
  assign RetimeWrapper_71_clock = clock; // @[:@14921.4]
  assign RetimeWrapper_71_reset = reset; // @[:@14922.4]
  assign RetimeWrapper_71_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14924.4]
  assign RetimeWrapper_71_io_in = _T_1493 & io_rPort_5_en_0; // @[package.scala 94:16:@14923.4]
  assign RetimeWrapper_72_clock = clock; // @[:@14977.4]
  assign RetimeWrapper_72_reset = reset; // @[:@14978.4]
  assign RetimeWrapper_72_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14980.4]
  assign RetimeWrapper_72_io_in = _T_487 & io_rPort_6_en_0; // @[package.scala 94:16:@14979.4]
  assign RetimeWrapper_73_clock = clock; // @[:@14985.4]
  assign RetimeWrapper_73_reset = reset; // @[:@14986.4]
  assign RetimeWrapper_73_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14988.4]
  assign RetimeWrapper_73_io_in = _T_579 & io_rPort_6_en_0; // @[package.scala 94:16:@14987.4]
  assign RetimeWrapper_74_clock = clock; // @[:@14993.4]
  assign RetimeWrapper_74_reset = reset; // @[:@14994.4]
  assign RetimeWrapper_74_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14996.4]
  assign RetimeWrapper_74_io_in = _T_671 & io_rPort_6_en_0; // @[package.scala 94:16:@14995.4]
  assign RetimeWrapper_75_clock = clock; // @[:@15001.4]
  assign RetimeWrapper_75_reset = reset; // @[:@15002.4]
  assign RetimeWrapper_75_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15004.4]
  assign RetimeWrapper_75_io_in = _T_763 & io_rPort_6_en_0; // @[package.scala 94:16:@15003.4]
  assign RetimeWrapper_76_clock = clock; // @[:@15009.4]
  assign RetimeWrapper_76_reset = reset; // @[:@15010.4]
  assign RetimeWrapper_76_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15012.4]
  assign RetimeWrapper_76_io_in = _T_855 & io_rPort_6_en_0; // @[package.scala 94:16:@15011.4]
  assign RetimeWrapper_77_clock = clock; // @[:@15017.4]
  assign RetimeWrapper_77_reset = reset; // @[:@15018.4]
  assign RetimeWrapper_77_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15020.4]
  assign RetimeWrapper_77_io_in = _T_947 & io_rPort_6_en_0; // @[package.scala 94:16:@15019.4]
  assign RetimeWrapper_78_clock = clock; // @[:@15025.4]
  assign RetimeWrapper_78_reset = reset; // @[:@15026.4]
  assign RetimeWrapper_78_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15028.4]
  assign RetimeWrapper_78_io_in = _T_1039 & io_rPort_6_en_0; // @[package.scala 94:16:@15027.4]
  assign RetimeWrapper_79_clock = clock; // @[:@15033.4]
  assign RetimeWrapper_79_reset = reset; // @[:@15034.4]
  assign RetimeWrapper_79_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15036.4]
  assign RetimeWrapper_79_io_in = _T_1131 & io_rPort_6_en_0; // @[package.scala 94:16:@15035.4]
  assign RetimeWrapper_80_clock = clock; // @[:@15041.4]
  assign RetimeWrapper_80_reset = reset; // @[:@15042.4]
  assign RetimeWrapper_80_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15044.4]
  assign RetimeWrapper_80_io_in = _T_1223 & io_rPort_6_en_0; // @[package.scala 94:16:@15043.4]
  assign RetimeWrapper_81_clock = clock; // @[:@15049.4]
  assign RetimeWrapper_81_reset = reset; // @[:@15050.4]
  assign RetimeWrapper_81_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15052.4]
  assign RetimeWrapper_81_io_in = _T_1315 & io_rPort_6_en_0; // @[package.scala 94:16:@15051.4]
  assign RetimeWrapper_82_clock = clock; // @[:@15057.4]
  assign RetimeWrapper_82_reset = reset; // @[:@15058.4]
  assign RetimeWrapper_82_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15060.4]
  assign RetimeWrapper_82_io_in = _T_1407 & io_rPort_6_en_0; // @[package.scala 94:16:@15059.4]
  assign RetimeWrapper_83_clock = clock; // @[:@15065.4]
  assign RetimeWrapper_83_reset = reset; // @[:@15066.4]
  assign RetimeWrapper_83_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15068.4]
  assign RetimeWrapper_83_io_in = _T_1499 & io_rPort_6_en_0; // @[package.scala 94:16:@15067.4]
  assign RetimeWrapper_84_clock = clock; // @[:@15121.4]
  assign RetimeWrapper_84_reset = reset; // @[:@15122.4]
  assign RetimeWrapper_84_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15124.4]
  assign RetimeWrapper_84_io_in = _T_493 & io_rPort_7_en_0; // @[package.scala 94:16:@15123.4]
  assign RetimeWrapper_85_clock = clock; // @[:@15129.4]
  assign RetimeWrapper_85_reset = reset; // @[:@15130.4]
  assign RetimeWrapper_85_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15132.4]
  assign RetimeWrapper_85_io_in = _T_585 & io_rPort_7_en_0; // @[package.scala 94:16:@15131.4]
  assign RetimeWrapper_86_clock = clock; // @[:@15137.4]
  assign RetimeWrapper_86_reset = reset; // @[:@15138.4]
  assign RetimeWrapper_86_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15140.4]
  assign RetimeWrapper_86_io_in = _T_677 & io_rPort_7_en_0; // @[package.scala 94:16:@15139.4]
  assign RetimeWrapper_87_clock = clock; // @[:@15145.4]
  assign RetimeWrapper_87_reset = reset; // @[:@15146.4]
  assign RetimeWrapper_87_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15148.4]
  assign RetimeWrapper_87_io_in = _T_769 & io_rPort_7_en_0; // @[package.scala 94:16:@15147.4]
  assign RetimeWrapper_88_clock = clock; // @[:@15153.4]
  assign RetimeWrapper_88_reset = reset; // @[:@15154.4]
  assign RetimeWrapper_88_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15156.4]
  assign RetimeWrapper_88_io_in = _T_861 & io_rPort_7_en_0; // @[package.scala 94:16:@15155.4]
  assign RetimeWrapper_89_clock = clock; // @[:@15161.4]
  assign RetimeWrapper_89_reset = reset; // @[:@15162.4]
  assign RetimeWrapper_89_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15164.4]
  assign RetimeWrapper_89_io_in = _T_953 & io_rPort_7_en_0; // @[package.scala 94:16:@15163.4]
  assign RetimeWrapper_90_clock = clock; // @[:@15169.4]
  assign RetimeWrapper_90_reset = reset; // @[:@15170.4]
  assign RetimeWrapper_90_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15172.4]
  assign RetimeWrapper_90_io_in = _T_1045 & io_rPort_7_en_0; // @[package.scala 94:16:@15171.4]
  assign RetimeWrapper_91_clock = clock; // @[:@15177.4]
  assign RetimeWrapper_91_reset = reset; // @[:@15178.4]
  assign RetimeWrapper_91_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15180.4]
  assign RetimeWrapper_91_io_in = _T_1137 & io_rPort_7_en_0; // @[package.scala 94:16:@15179.4]
  assign RetimeWrapper_92_clock = clock; // @[:@15185.4]
  assign RetimeWrapper_92_reset = reset; // @[:@15186.4]
  assign RetimeWrapper_92_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15188.4]
  assign RetimeWrapper_92_io_in = _T_1229 & io_rPort_7_en_0; // @[package.scala 94:16:@15187.4]
  assign RetimeWrapper_93_clock = clock; // @[:@15193.4]
  assign RetimeWrapper_93_reset = reset; // @[:@15194.4]
  assign RetimeWrapper_93_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15196.4]
  assign RetimeWrapper_93_io_in = _T_1321 & io_rPort_7_en_0; // @[package.scala 94:16:@15195.4]
  assign RetimeWrapper_94_clock = clock; // @[:@15201.4]
  assign RetimeWrapper_94_reset = reset; // @[:@15202.4]
  assign RetimeWrapper_94_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15204.4]
  assign RetimeWrapper_94_io_in = _T_1413 & io_rPort_7_en_0; // @[package.scala 94:16:@15203.4]
  assign RetimeWrapper_95_clock = clock; // @[:@15209.4]
  assign RetimeWrapper_95_reset = reset; // @[:@15210.4]
  assign RetimeWrapper_95_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15212.4]
  assign RetimeWrapper_95_io_in = _T_1505 & io_rPort_7_en_0; // @[package.scala 94:16:@15211.4]
  assign RetimeWrapper_96_clock = clock; // @[:@15265.4]
  assign RetimeWrapper_96_reset = reset; // @[:@15266.4]
  assign RetimeWrapper_96_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15268.4]
  assign RetimeWrapper_96_io_in = _T_499 & io_rPort_8_en_0; // @[package.scala 94:16:@15267.4]
  assign RetimeWrapper_97_clock = clock; // @[:@15273.4]
  assign RetimeWrapper_97_reset = reset; // @[:@15274.4]
  assign RetimeWrapper_97_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15276.4]
  assign RetimeWrapper_97_io_in = _T_591 & io_rPort_8_en_0; // @[package.scala 94:16:@15275.4]
  assign RetimeWrapper_98_clock = clock; // @[:@15281.4]
  assign RetimeWrapper_98_reset = reset; // @[:@15282.4]
  assign RetimeWrapper_98_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15284.4]
  assign RetimeWrapper_98_io_in = _T_683 & io_rPort_8_en_0; // @[package.scala 94:16:@15283.4]
  assign RetimeWrapper_99_clock = clock; // @[:@15289.4]
  assign RetimeWrapper_99_reset = reset; // @[:@15290.4]
  assign RetimeWrapper_99_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15292.4]
  assign RetimeWrapper_99_io_in = _T_775 & io_rPort_8_en_0; // @[package.scala 94:16:@15291.4]
  assign RetimeWrapper_100_clock = clock; // @[:@15297.4]
  assign RetimeWrapper_100_reset = reset; // @[:@15298.4]
  assign RetimeWrapper_100_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15300.4]
  assign RetimeWrapper_100_io_in = _T_867 & io_rPort_8_en_0; // @[package.scala 94:16:@15299.4]
  assign RetimeWrapper_101_clock = clock; // @[:@15305.4]
  assign RetimeWrapper_101_reset = reset; // @[:@15306.4]
  assign RetimeWrapper_101_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15308.4]
  assign RetimeWrapper_101_io_in = _T_959 & io_rPort_8_en_0; // @[package.scala 94:16:@15307.4]
  assign RetimeWrapper_102_clock = clock; // @[:@15313.4]
  assign RetimeWrapper_102_reset = reset; // @[:@15314.4]
  assign RetimeWrapper_102_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15316.4]
  assign RetimeWrapper_102_io_in = _T_1051 & io_rPort_8_en_0; // @[package.scala 94:16:@15315.4]
  assign RetimeWrapper_103_clock = clock; // @[:@15321.4]
  assign RetimeWrapper_103_reset = reset; // @[:@15322.4]
  assign RetimeWrapper_103_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15324.4]
  assign RetimeWrapper_103_io_in = _T_1143 & io_rPort_8_en_0; // @[package.scala 94:16:@15323.4]
  assign RetimeWrapper_104_clock = clock; // @[:@15329.4]
  assign RetimeWrapper_104_reset = reset; // @[:@15330.4]
  assign RetimeWrapper_104_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15332.4]
  assign RetimeWrapper_104_io_in = _T_1235 & io_rPort_8_en_0; // @[package.scala 94:16:@15331.4]
  assign RetimeWrapper_105_clock = clock; // @[:@15337.4]
  assign RetimeWrapper_105_reset = reset; // @[:@15338.4]
  assign RetimeWrapper_105_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15340.4]
  assign RetimeWrapper_105_io_in = _T_1327 & io_rPort_8_en_0; // @[package.scala 94:16:@15339.4]
  assign RetimeWrapper_106_clock = clock; // @[:@15345.4]
  assign RetimeWrapper_106_reset = reset; // @[:@15346.4]
  assign RetimeWrapper_106_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15348.4]
  assign RetimeWrapper_106_io_in = _T_1419 & io_rPort_8_en_0; // @[package.scala 94:16:@15347.4]
  assign RetimeWrapper_107_clock = clock; // @[:@15353.4]
  assign RetimeWrapper_107_reset = reset; // @[:@15354.4]
  assign RetimeWrapper_107_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15356.4]
  assign RetimeWrapper_107_io_in = _T_1511 & io_rPort_8_en_0; // @[package.scala 94:16:@15355.4]
endmodule
module Divider( // @[:@16978.2]
  input         clock, // @[:@16979.4]
  input         io_flow, // @[:@16981.4]
  input  [31:0] io_dividend, // @[:@16981.4]
  input  [31:0] io_divisor, // @[:@16981.4]
  output [31:0] io_out // @[:@16981.4]
);
  wire [31:0] m_m_axis_dout_tdata; // @[ZynqBlackBoxes.scala 26:19:@16983.4]
  wire  m_m_axis_dout_tvalid; // @[ZynqBlackBoxes.scala 26:19:@16983.4]
  wire [31:0] m_s_axis_divisor_tdata; // @[ZynqBlackBoxes.scala 26:19:@16983.4]
  wire  m_s_axis_divisor_tvalid; // @[ZynqBlackBoxes.scala 26:19:@16983.4]
  wire [31:0] m_s_axis_dividend_tdata; // @[ZynqBlackBoxes.scala 26:19:@16983.4]
  wire  m_s_axis_dividend_tvalid; // @[ZynqBlackBoxes.scala 26:19:@16983.4]
  wire  m_aclken; // @[ZynqBlackBoxes.scala 26:19:@16983.4]
  wire  m_aclk; // @[ZynqBlackBoxes.scala 26:19:@16983.4]
  wire [29:0] _T_15; // @[ZynqBlackBoxes.scala 34:37:@16999.4]
  div_32_32_20_Signed_Fractional m ( // @[ZynqBlackBoxes.scala 26:19:@16983.4]
    .m_axis_dout_tdata(m_m_axis_dout_tdata),
    .m_axis_dout_tvalid(m_m_axis_dout_tvalid),
    .s_axis_divisor_tdata(m_s_axis_divisor_tdata),
    .s_axis_divisor_tvalid(m_s_axis_divisor_tvalid),
    .s_axis_dividend_tdata(m_s_axis_dividend_tdata),
    .s_axis_dividend_tvalid(m_s_axis_dividend_tvalid),
    .aclken(m_aclken),
    .aclk(m_aclk)
  );
  assign _T_15 = m_m_axis_dout_tdata[31:2]; // @[ZynqBlackBoxes.scala 34:37:@16999.4]
  assign io_out = {{2'd0}, _T_15}; // @[ZynqBlackBoxes.scala 34:12:@17000.4]
  assign m_s_axis_divisor_tdata = io_divisor; // @[ZynqBlackBoxes.scala 32:31:@16997.4]
  assign m_s_axis_divisor_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 31:32:@16996.4]
  assign m_s_axis_dividend_tdata = io_dividend; // @[ZynqBlackBoxes.scala 30:32:@16995.4]
  assign m_s_axis_dividend_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 29:33:@16994.4]
  assign m_aclken = io_flow; // @[ZynqBlackBoxes.scala 28:17:@16993.4 ZynqBlackBoxes.scala 33:17:@16998.4]
  assign m_aclk = clock; // @[ZynqBlackBoxes.scala 27:15:@16992.4]
endmodule
module x225_div( // @[:@17038.2]
  input         clock, // @[:@17039.4]
  input  [31:0] io_a, // @[:@17041.4]
  input         io_flow, // @[:@17041.4]
  output [31:0] io_result // @[:@17041.4]
);
  wire  x225_div_clock; // @[BigIPZynq.scala 25:21:@17049.4]
  wire  x225_div_io_flow; // @[BigIPZynq.scala 25:21:@17049.4]
  wire [31:0] x225_div_io_dividend; // @[BigIPZynq.scala 25:21:@17049.4]
  wire [31:0] x225_div_io_divisor; // @[BigIPZynq.scala 25:21:@17049.4]
  wire [31:0] x225_div_io_out; // @[BigIPZynq.scala 25:21:@17049.4]
  wire [31:0] __io_b; // @[Math.scala 720:24:@17062.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@17062.4]
  wire [31:0] _T_15; // @[FixedPoint.scala 24:59:@17047.4]
  wire [31:0] _T_19; // @[BigIPZynq.scala 29:16:@17057.4]
  Divider x225_div ( // @[BigIPZynq.scala 25:21:@17049.4]
    .clock(x225_div_clock),
    .io_flow(x225_div_io_flow),
    .io_dividend(x225_div_io_dividend),
    .io_divisor(x225_div_io_divisor),
    .io_out(x225_div_io_out)
  );
  _ _ ( // @[Math.scala 720:24:@17062.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  assign _T_15 = $signed(io_a); // @[FixedPoint.scala 24:59:@17047.4]
  assign _T_19 = $signed(x225_div_io_out); // @[BigIPZynq.scala 29:16:@17057.4]
  assign io_result = __io_result; // @[Math.scala 290:34:@17070.4]
  assign x225_div_clock = clock; // @[:@17050.4]
  assign x225_div_io_flow = io_flow; // @[BigIPZynq.scala 28:17:@17056.4]
  assign x225_div_io_dividend = $unsigned(_T_15); // @[BigIPZynq.scala 26:21:@17053.4]
  assign x225_div_io_divisor = 32'h3; // @[BigIPZynq.scala 27:20:@17055.4]
  assign __io_b = $unsigned(_T_19); // @[Math.scala 721:17:@17065.4]
endmodule
module RetimeWrapper_184( // @[:@17084.2]
  input         clock, // @[:@17085.4]
  input         reset, // @[:@17086.4]
  input         io_flow, // @[:@17087.4]
  input  [31:0] io_in, // @[:@17087.4]
  output [31:0] io_out // @[:@17087.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17089.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17089.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17089.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17089.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17089.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17089.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(19)) sr ( // @[RetimeShiftRegister.scala 15:20:@17089.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17102.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17101.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17100.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17099.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17098.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17096.4]
endmodule
module RetimeWrapper_186( // @[:@17295.2]
  input         clock, // @[:@17296.4]
  input         reset, // @[:@17297.4]
  input         io_flow, // @[:@17298.4]
  input  [31:0] io_in, // @[:@17298.4]
  output [31:0] io_out // @[:@17298.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17300.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17300.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17300.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17300.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17300.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17300.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(13)) sr ( // @[RetimeShiftRegister.scala 15:20:@17300.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17313.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17312.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17311.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17310.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17309.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17307.4]
endmodule
module RetimeWrapper_187( // @[:@17327.2]
  input         clock, // @[:@17328.4]
  input         reset, // @[:@17329.4]
  input         io_flow, // @[:@17330.4]
  input  [31:0] io_in, // @[:@17330.4]
  output [31:0] io_out // @[:@17330.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17332.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17332.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17332.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17332.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17332.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17332.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@17332.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17345.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17344.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17343.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17342.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17341.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17339.4]
endmodule
module RetimeWrapper_188( // @[:@17359.2]
  input         clock, // @[:@17360.4]
  input         reset, // @[:@17361.4]
  input         io_flow, // @[:@17362.4]
  input  [31:0] io_in, // @[:@17362.4]
  output [31:0] io_out // @[:@17362.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17364.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17364.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17364.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17364.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17364.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17364.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@17364.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17377.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17376.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17375.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17374.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17373.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17371.4]
endmodule
module RetimeWrapper_189( // @[:@17391.2]
  input   clock, // @[:@17392.4]
  input   reset, // @[:@17393.4]
  input   io_flow, // @[:@17394.4]
  input   io_in, // @[:@17394.4]
  output  io_out // @[:@17394.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@17396.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@17396.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@17396.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17396.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17396.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17396.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@17396.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17409.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17408.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@17407.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17406.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17405.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17403.4]
endmodule
module RetimeWrapper_192( // @[:@17487.2]
  input         clock, // @[:@17488.4]
  input         reset, // @[:@17489.4]
  input         io_flow, // @[:@17490.4]
  input  [31:0] io_in, // @[:@17490.4]
  output [31:0] io_out // @[:@17490.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17492.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17492.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17492.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17492.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17492.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17492.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(23)) sr ( // @[RetimeShiftRegister.scala 15:20:@17492.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17505.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17504.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17503.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17502.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17501.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17499.4]
endmodule
module RetimeWrapper_196( // @[:@17615.2]
  input         clock, // @[:@17616.4]
  input         reset, // @[:@17617.4]
  input         io_flow, // @[:@17618.4]
  input  [31:0] io_in, // @[:@17618.4]
  output [31:0] io_out // @[:@17618.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17620.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17620.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17620.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17620.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17620.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17620.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(37)) sr ( // @[RetimeShiftRegister.scala 15:20:@17620.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17633.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17632.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17631.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17630.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17629.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17627.4]
endmodule
module RetimeWrapper_197( // @[:@17647.2]
  input         clock, // @[:@17648.4]
  input         reset, // @[:@17649.4]
  input         io_flow, // @[:@17650.4]
  input  [31:0] io_in, // @[:@17650.4]
  output [31:0] io_out // @[:@17650.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17652.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17652.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17652.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17652.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17652.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17652.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(45)) sr ( // @[RetimeShiftRegister.scala 15:20:@17652.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17665.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17664.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17663.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17662.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17661.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17659.4]
endmodule
module RetimeWrapper_198( // @[:@17679.2]
  input   clock, // @[:@17680.4]
  input   reset, // @[:@17681.4]
  input   io_flow, // @[:@17682.4]
  input   io_in, // @[:@17682.4]
  output  io_out // @[:@17682.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@17684.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@17684.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@17684.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17684.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17684.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17684.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(45)) sr ( // @[RetimeShiftRegister.scala 15:20:@17684.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17697.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17696.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@17695.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17694.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17693.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17691.4]
endmodule
module RetimeWrapper_199( // @[:@17711.2]
  input         clock, // @[:@17712.4]
  input         reset, // @[:@17713.4]
  input         io_flow, // @[:@17714.4]
  input  [31:0] io_in, // @[:@17714.4]
  output [31:0] io_out // @[:@17714.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17716.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17716.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17716.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17716.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17716.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17716.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(24)) sr ( // @[RetimeShiftRegister.scala 15:20:@17716.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17729.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17728.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17727.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17726.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17725.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17723.4]
endmodule
module RetimeWrapper_218( // @[:@19604.2]
  input         clock, // @[:@19605.4]
  input         reset, // @[:@19606.4]
  input         io_flow, // @[:@19607.4]
  input  [31:0] io_in, // @[:@19607.4]
  output [31:0] io_out // @[:@19607.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@19609.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@19609.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@19609.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@19609.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@19609.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@19609.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(43)) sr ( // @[RetimeShiftRegister.scala 15:20:@19609.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@19622.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@19621.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@19620.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@19619.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@19618.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@19616.4]
endmodule
module RetimeWrapper_220( // @[:@19815.2]
  input   clock, // @[:@19816.4]
  input   reset, // @[:@19817.4]
  input   io_flow, // @[:@19818.4]
  input   io_in, // @[:@19818.4]
  output  io_out // @[:@19818.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@19820.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@19820.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@19820.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@19820.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@19820.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@19820.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@19820.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@19833.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@19832.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@19831.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@19830.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@19829.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@19827.4]
endmodule
module RetimeWrapper_248( // @[:@22438.2]
  input         clock, // @[:@22439.4]
  input         reset, // @[:@22440.4]
  input         io_flow, // @[:@22441.4]
  input  [31:0] io_in, // @[:@22441.4]
  output [31:0] io_out // @[:@22441.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@22443.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@22443.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@22443.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22443.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22443.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22443.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(17)) sr ( // @[RetimeShiftRegister.scala 15:20:@22443.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22456.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22455.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@22454.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22453.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22452.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22450.4]
endmodule
module RetimeWrapper_254( // @[:@22777.2]
  input         clock, // @[:@22778.4]
  input         reset, // @[:@22779.4]
  input         io_flow, // @[:@22780.4]
  input  [31:0] io_in, // @[:@22780.4]
  output [31:0] io_out // @[:@22780.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@22782.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@22782.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@22782.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@22782.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@22782.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@22782.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(18)) sr ( // @[RetimeShiftRegister.scala 15:20:@22782.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@22795.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@22794.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@22793.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@22792.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@22791.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@22789.4]
endmodule
module Multiplier( // @[:@24605.2]
  input         clock, // @[:@24606.4]
  input         io_flow, // @[:@24608.4]
  input  [31:0] io_a, // @[:@24608.4]
  input  [31:0] io_b, // @[:@24608.4]
  output [31:0] io_out // @[:@24608.4]
);
  wire [31:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@24610.4]
  wire [31:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@24610.4]
  wire [31:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@24610.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@24610.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@24610.4]
  mul_32_32_32_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@24610.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@24620.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@24618.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@24617.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@24619.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@24616.4]
endmodule
module x295( // @[:@24640.2]
  input         clock, // @[:@24641.4]
  input  [31:0] io_a, // @[:@24643.4]
  input  [31:0] io_b, // @[:@24643.4]
  input         io_flow, // @[:@24643.4]
  output [31:0] io_result // @[:@24643.4]
);
  wire  x295_clock; // @[BigIPZynq.scala 63:21:@24650.4]
  wire  x295_io_flow; // @[BigIPZynq.scala 63:21:@24650.4]
  wire [31:0] x295_io_a; // @[BigIPZynq.scala 63:21:@24650.4]
  wire [31:0] x295_io_b; // @[BigIPZynq.scala 63:21:@24650.4]
  wire [31:0] x295_io_out; // @[BigIPZynq.scala 63:21:@24650.4]
  wire [31:0] fix2fixBox_io_a; // @[Math.scala 253:30:@24659.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@24659.4]
  Multiplier x295 ( // @[BigIPZynq.scala 63:21:@24650.4]
    .clock(x295_clock),
    .io_flow(x295_io_flow),
    .io_a(x295_io_a),
    .io_b(x295_io_b),
    .io_out(x295_io_out)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 253:30:@24659.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@24667.4]
  assign x295_clock = clock; // @[:@24651.4]
  assign x295_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@24655.4]
  assign x295_io_a = io_a; // @[BigIPZynq.scala 64:14:@24653.4]
  assign x295_io_b = io_b; // @[BigIPZynq.scala 65:14:@24654.4]
  assign fix2fixBox_io_a = x295_io_out; // @[Math.scala 254:23:@24662.4]
endmodule
module fix2fixBox_140( // @[:@25261.2]
  input  [31:0] io_a, // @[:@25264.4]
  output [32:0] io_b // @[:@25264.4]
);
  assign io_b = {1'h0,io_a}; // @[Converter.scala 95:38:@25278.4]
endmodule
module __89( // @[:@25280.2]
  input  [31:0] io_b, // @[:@25283.4]
  output [32:0] io_result // @[:@25283.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@25288.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@25288.4]
  fix2fixBox_140 fix2fixBox ( // @[BigIPZynq.scala 219:30:@25288.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@25296.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@25291.4]
endmodule
module x304_x3( // @[:@25392.2]
  input         clock, // @[:@25393.4]
  input         reset, // @[:@25394.4]
  input  [31:0] io_a, // @[:@25395.4]
  input  [31:0] io_b, // @[:@25395.4]
  input         io_flow, // @[:@25395.4]
  output [31:0] io_result // @[:@25395.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@25403.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@25403.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@25410.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@25410.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@25420.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@25420.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@25420.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@25420.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@25420.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@25408.4 Math.scala 724:14:@25409.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@25415.4 Math.scala 724:14:@25416.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@25417.4]
  __89 _ ( // @[Math.scala 720:24:@25403.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __89 __1 ( // @[Math.scala 720:24:@25410.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@25420.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@25408.4 Math.scala 724:14:@25409.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@25415.4 Math.scala 724:14:@25416.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@25417.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@25428.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@25406.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@25413.4]
  assign fix2fixBox_clock = clock; // @[:@25421.4]
  assign fix2fixBox_reset = reset; // @[:@25422.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@25423.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@25426.4]
endmodule
module RetimeWrapper_286( // @[:@26456.2]
  input         clock, // @[:@26457.4]
  input         reset, // @[:@26458.4]
  input         io_flow, // @[:@26459.4]
  input  [31:0] io_in, // @[:@26459.4]
  output [31:0] io_out // @[:@26459.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26461.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26461.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26461.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26461.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26461.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26461.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@26461.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26474.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26473.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@26472.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26471.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26470.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26468.4]
endmodule
module fix2fixBox_164( // @[:@26645.2]
  input  [31:0] io_a, // @[:@26648.4]
  output [31:0] io_b // @[:@26648.4]
);
  wire [24:0] new_dec; // @[Converter.scala 63:26:@26658.4]
  assign new_dec = io_a[24:0]; // @[Converter.scala 63:26:@26658.4]
  assign io_b = {new_dec,7'h0}; // @[Converter.scala 94:38:@26661.4]
endmodule
module x312( // @[:@26663.2]
  input  [31:0] io_b, // @[:@26666.4]
  output [31:0] io_result // @[:@26666.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@26671.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@26671.4]
  fix2fixBox_164 fix2fixBox ( // @[BigIPZynq.scala 219:30:@26671.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@26679.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@26674.4]
endmodule
module Multiplier_9( // @[:@26691.2]
  input         clock, // @[:@26692.4]
  input         io_flow, // @[:@26694.4]
  input  [38:0] io_a, // @[:@26694.4]
  output [38:0] io_out // @[:@26694.4]
);
  wire [38:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@26696.4]
  wire [38:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@26696.4]
  wire [38:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@26696.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@26696.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@26696.4]
  mul_39_39_39_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@26696.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@26706.4]
  assign m_B = 39'h8; // @[ZynqBlackBoxes.scala 107:12:@26704.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@26703.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@26705.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@26702.4]
endmodule
module fix2fixBox_165( // @[:@26708.2]
  input  [38:0] io_a, // @[:@26711.4]
  output [31:0] io_b // @[:@26711.4]
);
  wire [6:0] tmp_frac; // @[Converter.scala 38:42:@26719.4]
  wire [24:0] new_dec; // @[Converter.scala 88:34:@26722.4]
  assign tmp_frac = io_a[13:7]; // @[Converter.scala 38:42:@26719.4]
  assign new_dec = io_a[38:14]; // @[Converter.scala 88:34:@26722.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@26725.4]
endmodule
module x313_mul( // @[:@26727.2]
  input         clock, // @[:@26728.4]
  input  [31:0] io_a, // @[:@26730.4]
  input         io_flow, // @[:@26730.4]
  output [31:0] io_result // @[:@26730.4]
);
  wire  x313_mul_clock; // @[BigIPZynq.scala 63:21:@26745.4]
  wire  x313_mul_io_flow; // @[BigIPZynq.scala 63:21:@26745.4]
  wire [38:0] x313_mul_io_a; // @[BigIPZynq.scala 63:21:@26745.4]
  wire [38:0] x313_mul_io_out; // @[BigIPZynq.scala 63:21:@26745.4]
  wire [38:0] fix2fixBox_io_a; // @[Math.scala 253:30:@26753.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@26753.4]
  wire  _T_16; // @[FixedPoint.scala 50:25:@26737.4]
  wire [6:0] _T_20; // @[Bitwise.scala 72:12:@26739.4]
  Multiplier_9 x313_mul ( // @[BigIPZynq.scala 63:21:@26745.4]
    .clock(x313_mul_clock),
    .io_flow(x313_mul_io_flow),
    .io_a(x313_mul_io_a),
    .io_out(x313_mul_io_out)
  );
  fix2fixBox_165 fix2fixBox ( // @[Math.scala 253:30:@26753.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_16 = io_a[31]; // @[FixedPoint.scala 50:25:@26737.4]
  assign _T_20 = _T_16 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@26739.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@26761.4]
  assign x313_mul_clock = clock; // @[:@26746.4]
  assign x313_mul_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@26750.4]
  assign x313_mul_io_a = {_T_20,io_a}; // @[BigIPZynq.scala 64:14:@26748.4]
  assign fix2fixBox_io_a = x313_mul_io_out; // @[Math.scala 254:23:@26756.4]
endmodule
module fix2fixBox_166( // @[:@26763.2]
  input  [31:0] io_a, // @[:@26766.4]
  output [31:0] io_b // @[:@26766.4]
);
  wire [24:0] _T_25; // @[Converter.scala 84:75:@26778.4]
  assign _T_25 = io_a[31:7]; // @[Converter.scala 84:75:@26778.4]
  assign io_b = {7'h0,_T_25}; // @[Converter.scala 95:38:@26781.4]
endmodule
module x314( // @[:@26783.2]
  input  [31:0] io_b, // @[:@26786.4]
  output [31:0] io_result // @[:@26786.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@26791.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@26791.4]
  fix2fixBox_166 fix2fixBox ( // @[BigIPZynq.scala 219:30:@26791.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@26799.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@26794.4]
endmodule
module x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@26929.2]
  input          clock, // @[:@26930.4]
  input          reset, // @[:@26931.4]
  output         io_in_x185_TVALID, // @[:@26932.4]
  input          io_in_x185_TREADY, // @[:@26932.4]
  output [255:0] io_in_x185_TDATA, // @[:@26932.4]
  output         io_in_x184_TREADY, // @[:@26932.4]
  input  [255:0] io_in_x184_TDATA, // @[:@26932.4]
  input  [7:0]   io_in_x184_TID, // @[:@26932.4]
  input  [7:0]   io_in_x184_TDEST, // @[:@26932.4]
  input          io_sigsIn_backpressure, // @[:@26932.4]
  input          io_sigsIn_datapathEn, // @[:@26932.4]
  input          io_sigsIn_break, // @[:@26932.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@26932.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@26932.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@26932.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@26932.4]
  input          io_rr // @[:@26932.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@26946.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@26946.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@26958.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@26958.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@26981.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@26981.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@26981.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@26981.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@26981.4]
  wire  x217_lb_0_clock; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_reset; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [1:0] x217_lb_0_io_rPort_8_banks_1; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [2:0] x217_lb_0_io_rPort_8_banks_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [9:0] x217_lb_0_io_rPort_8_ofs_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_rPort_8_en_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_rPort_8_backpressure; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [31:0] x217_lb_0_io_rPort_8_output_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [1:0] x217_lb_0_io_rPort_7_banks_1; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [2:0] x217_lb_0_io_rPort_7_banks_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [9:0] x217_lb_0_io_rPort_7_ofs_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_rPort_7_en_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_rPort_7_backpressure; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [31:0] x217_lb_0_io_rPort_7_output_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [1:0] x217_lb_0_io_rPort_6_banks_1; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [2:0] x217_lb_0_io_rPort_6_banks_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [9:0] x217_lb_0_io_rPort_6_ofs_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_rPort_6_en_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_rPort_6_backpressure; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [31:0] x217_lb_0_io_rPort_6_output_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [1:0] x217_lb_0_io_rPort_5_banks_1; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [2:0] x217_lb_0_io_rPort_5_banks_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [9:0] x217_lb_0_io_rPort_5_ofs_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_rPort_5_en_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_rPort_5_backpressure; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [31:0] x217_lb_0_io_rPort_5_output_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [1:0] x217_lb_0_io_rPort_4_banks_1; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [2:0] x217_lb_0_io_rPort_4_banks_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [9:0] x217_lb_0_io_rPort_4_ofs_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_rPort_4_en_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_rPort_4_backpressure; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [31:0] x217_lb_0_io_rPort_4_output_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [1:0] x217_lb_0_io_rPort_3_banks_1; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [2:0] x217_lb_0_io_rPort_3_banks_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [9:0] x217_lb_0_io_rPort_3_ofs_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_rPort_3_en_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_rPort_3_backpressure; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [31:0] x217_lb_0_io_rPort_3_output_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [1:0] x217_lb_0_io_rPort_2_banks_1; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [2:0] x217_lb_0_io_rPort_2_banks_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [9:0] x217_lb_0_io_rPort_2_ofs_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_rPort_2_en_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_rPort_2_backpressure; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [31:0] x217_lb_0_io_rPort_2_output_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [1:0] x217_lb_0_io_rPort_1_banks_1; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [2:0] x217_lb_0_io_rPort_1_banks_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [9:0] x217_lb_0_io_rPort_1_ofs_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_rPort_1_en_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_rPort_1_backpressure; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [31:0] x217_lb_0_io_rPort_1_output_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [1:0] x217_lb_0_io_rPort_0_banks_1; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [2:0] x217_lb_0_io_rPort_0_banks_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [9:0] x217_lb_0_io_rPort_0_ofs_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_rPort_0_en_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_rPort_0_backpressure; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [31:0] x217_lb_0_io_rPort_0_output_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [1:0] x217_lb_0_io_wPort_0_banks_1; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [2:0] x217_lb_0_io_wPort_0_banks_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [9:0] x217_lb_0_io_wPort_0_ofs_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire [31:0] x217_lb_0_io_wPort_0_data_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x217_lb_0_io_wPort_0_en_0; // @[m_x217_lb_0.scala 35:17:@26991.4]
  wire  x378_sum_1_clock; // @[Math.scala 150:24:@27116.4]
  wire  x378_sum_1_reset; // @[Math.scala 150:24:@27116.4]
  wire [31:0] x378_sum_1_io_a; // @[Math.scala 150:24:@27116.4]
  wire [31:0] x378_sum_1_io_b; // @[Math.scala 150:24:@27116.4]
  wire  x378_sum_1_io_flow; // @[Math.scala 150:24:@27116.4]
  wire [31:0] x378_sum_1_io_result; // @[Math.scala 150:24:@27116.4]
  wire  x381_sum_1_clock; // @[Math.scala 150:24:@27154.4]
  wire  x381_sum_1_reset; // @[Math.scala 150:24:@27154.4]
  wire [31:0] x381_sum_1_io_a; // @[Math.scala 150:24:@27154.4]
  wire [31:0] x381_sum_1_io_b; // @[Math.scala 150:24:@27154.4]
  wire  x381_sum_1_io_flow; // @[Math.scala 150:24:@27154.4]
  wire [31:0] x381_sum_1_io_result; // @[Math.scala 150:24:@27154.4]
  wire  x384_sum_1_clock; // @[Math.scala 150:24:@27192.4]
  wire  x384_sum_1_reset; // @[Math.scala 150:24:@27192.4]
  wire [31:0] x384_sum_1_io_a; // @[Math.scala 150:24:@27192.4]
  wire [31:0] x384_sum_1_io_b; // @[Math.scala 150:24:@27192.4]
  wire  x384_sum_1_io_flow; // @[Math.scala 150:24:@27192.4]
  wire [31:0] x384_sum_1_io_result; // @[Math.scala 150:24:@27192.4]
  wire  x387_sum_1_clock; // @[Math.scala 150:24:@27230.4]
  wire  x387_sum_1_reset; // @[Math.scala 150:24:@27230.4]
  wire [31:0] x387_sum_1_io_a; // @[Math.scala 150:24:@27230.4]
  wire [31:0] x387_sum_1_io_b; // @[Math.scala 150:24:@27230.4]
  wire  x387_sum_1_io_flow; // @[Math.scala 150:24:@27230.4]
  wire [31:0] x387_sum_1_io_result; // @[Math.scala 150:24:@27230.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@27253.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@27253.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@27253.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@27253.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@27253.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@27271.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@27271.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@27271.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@27271.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@27271.4]
  wire  x390_sum_1_clock; // @[Math.scala 150:24:@27284.4]
  wire  x390_sum_1_reset; // @[Math.scala 150:24:@27284.4]
  wire [31:0] x390_sum_1_io_a; // @[Math.scala 150:24:@27284.4]
  wire [31:0] x390_sum_1_io_b; // @[Math.scala 150:24:@27284.4]
  wire  x390_sum_1_io_flow; // @[Math.scala 150:24:@27284.4]
  wire [31:0] x390_sum_1_io_result; // @[Math.scala 150:24:@27284.4]
  wire  x393_sum_1_clock; // @[Math.scala 150:24:@27322.4]
  wire  x393_sum_1_reset; // @[Math.scala 150:24:@27322.4]
  wire [31:0] x393_sum_1_io_a; // @[Math.scala 150:24:@27322.4]
  wire [31:0] x393_sum_1_io_b; // @[Math.scala 150:24:@27322.4]
  wire  x393_sum_1_io_flow; // @[Math.scala 150:24:@27322.4]
  wire [31:0] x393_sum_1_io_result; // @[Math.scala 150:24:@27322.4]
  wire  x396_sub_1_clock; // @[Math.scala 191:24:@27348.4]
  wire  x396_sub_1_reset; // @[Math.scala 191:24:@27348.4]
  wire [31:0] x396_sub_1_io_a; // @[Math.scala 191:24:@27348.4]
  wire [31:0] x396_sub_1_io_b; // @[Math.scala 191:24:@27348.4]
  wire  x396_sub_1_io_flow; // @[Math.scala 191:24:@27348.4]
  wire [31:0] x396_sub_1_io_result; // @[Math.scala 191:24:@27348.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@27358.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@27358.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@27358.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@27358.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@27358.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@27367.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@27367.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@27367.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@27367.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@27367.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@27376.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@27376.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@27376.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@27376.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@27376.4]
  wire  x400_sum_1_clock; // @[Math.scala 150:24:@27415.4]
  wire  x400_sum_1_reset; // @[Math.scala 150:24:@27415.4]
  wire [31:0] x400_sum_1_io_a; // @[Math.scala 150:24:@27415.4]
  wire [31:0] x400_sum_1_io_b; // @[Math.scala 150:24:@27415.4]
  wire  x400_sum_1_io_flow; // @[Math.scala 150:24:@27415.4]
  wire [31:0] x400_sum_1_io_result; // @[Math.scala 150:24:@27415.4]
  wire  x225_div_1_clock; // @[Math.scala 327:24:@27427.4]
  wire [31:0] x225_div_1_io_a; // @[Math.scala 327:24:@27427.4]
  wire  x225_div_1_io_flow; // @[Math.scala 327:24:@27427.4]
  wire [31:0] x225_div_1_io_result; // @[Math.scala 327:24:@27427.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@27437.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@27437.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@27437.4]
  wire [31:0] RetimeWrapper_6_io_in; // @[package.scala 93:22:@27437.4]
  wire [31:0] RetimeWrapper_6_io_out; // @[package.scala 93:22:@27437.4]
  wire  x226_sum_1_clock; // @[Math.scala 150:24:@27446.4]
  wire  x226_sum_1_reset; // @[Math.scala 150:24:@27446.4]
  wire [31:0] x226_sum_1_io_a; // @[Math.scala 150:24:@27446.4]
  wire [31:0] x226_sum_1_io_b; // @[Math.scala 150:24:@27446.4]
  wire  x226_sum_1_io_flow; // @[Math.scala 150:24:@27446.4]
  wire [31:0] x226_sum_1_io_result; // @[Math.scala 150:24:@27446.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@27456.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@27456.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@27456.4]
  wire [31:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@27456.4]
  wire [31:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@27456.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@27465.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@27465.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@27465.4]
  wire [31:0] RetimeWrapper_8_io_in; // @[package.scala 93:22:@27465.4]
  wire [31:0] RetimeWrapper_8_io_out; // @[package.scala 93:22:@27465.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@27474.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@27474.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@27474.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@27474.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@27474.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@27483.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@27483.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@27483.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@27483.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@27483.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@27492.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@27492.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@27492.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@27492.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@27492.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@27503.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@27503.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@27503.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@27503.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@27503.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@27524.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@27524.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@27524.4]
  wire [31:0] RetimeWrapper_13_io_in; // @[package.scala 93:22:@27524.4]
  wire [31:0] RetimeWrapper_13_io_out; // @[package.scala 93:22:@27524.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@27538.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@27538.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@27538.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@27538.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@27538.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@27547.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@27547.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@27547.4]
  wire [31:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@27547.4]
  wire [31:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@27547.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@27563.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@27563.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@27563.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@27563.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@27563.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@27578.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@27578.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@27578.4]
  wire [31:0] RetimeWrapper_17_io_in; // @[package.scala 93:22:@27578.4]
  wire [31:0] RetimeWrapper_17_io_out; // @[package.scala 93:22:@27578.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@27587.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@27587.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@27587.4]
  wire [31:0] RetimeWrapper_18_io_in; // @[package.scala 93:22:@27587.4]
  wire [31:0] RetimeWrapper_18_io_out; // @[package.scala 93:22:@27587.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@27596.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@27596.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@27596.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@27596.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@27596.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@27605.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@27605.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@27605.4]
  wire [31:0] RetimeWrapper_20_io_in; // @[package.scala 93:22:@27605.4]
  wire [31:0] RetimeWrapper_20_io_out; // @[package.scala 93:22:@27605.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@27614.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@27614.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@27614.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@27614.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@27614.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@27623.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@27623.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@27623.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@27623.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@27623.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@27635.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@27635.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@27635.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@27635.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@27635.4]
  wire  x235_rdcol_1_clock; // @[Math.scala 191:24:@27658.4]
  wire  x235_rdcol_1_reset; // @[Math.scala 191:24:@27658.4]
  wire [31:0] x235_rdcol_1_io_a; // @[Math.scala 191:24:@27658.4]
  wire [31:0] x235_rdcol_1_io_b; // @[Math.scala 191:24:@27658.4]
  wire  x235_rdcol_1_io_flow; // @[Math.scala 191:24:@27658.4]
  wire [31:0] x235_rdcol_1_io_result; // @[Math.scala 191:24:@27658.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@27673.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@27673.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@27673.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@27673.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@27673.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@27682.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@27682.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@27682.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@27682.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@27682.4]
  wire  x403_sum_1_clock; // @[Math.scala 150:24:@27725.4]
  wire  x403_sum_1_reset; // @[Math.scala 150:24:@27725.4]
  wire [31:0] x403_sum_1_io_a; // @[Math.scala 150:24:@27725.4]
  wire [31:0] x403_sum_1_io_b; // @[Math.scala 150:24:@27725.4]
  wire  x403_sum_1_io_flow; // @[Math.scala 150:24:@27725.4]
  wire [31:0] x403_sum_1_io_result; // @[Math.scala 150:24:@27725.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@27748.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@27748.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@27748.4]
  wire [31:0] RetimeWrapper_26_io_in; // @[package.scala 93:22:@27748.4]
  wire [31:0] RetimeWrapper_26_io_out; // @[package.scala 93:22:@27748.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@27766.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@27766.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@27766.4]
  wire [31:0] RetimeWrapper_27_io_in; // @[package.scala 93:22:@27766.4]
  wire [31:0] RetimeWrapper_27_io_out; // @[package.scala 93:22:@27766.4]
  wire  x406_sum_1_clock; // @[Math.scala 150:24:@27779.4]
  wire  x406_sum_1_reset; // @[Math.scala 150:24:@27779.4]
  wire [31:0] x406_sum_1_io_a; // @[Math.scala 150:24:@27779.4]
  wire [31:0] x406_sum_1_io_b; // @[Math.scala 150:24:@27779.4]
  wire  x406_sum_1_io_flow; // @[Math.scala 150:24:@27779.4]
  wire [31:0] x406_sum_1_io_result; // @[Math.scala 150:24:@27779.4]
  wire  x409_sum_1_clock; // @[Math.scala 150:24:@27817.4]
  wire  x409_sum_1_reset; // @[Math.scala 150:24:@27817.4]
  wire [31:0] x409_sum_1_io_a; // @[Math.scala 150:24:@27817.4]
  wire [31:0] x409_sum_1_io_b; // @[Math.scala 150:24:@27817.4]
  wire  x409_sum_1_io_flow; // @[Math.scala 150:24:@27817.4]
  wire [31:0] x409_sum_1_io_result; // @[Math.scala 150:24:@27817.4]
  wire  x412_sum_1_clock; // @[Math.scala 150:24:@27855.4]
  wire  x412_sum_1_reset; // @[Math.scala 150:24:@27855.4]
  wire [31:0] x412_sum_1_io_a; // @[Math.scala 150:24:@27855.4]
  wire [31:0] x412_sum_1_io_b; // @[Math.scala 150:24:@27855.4]
  wire  x412_sum_1_io_flow; // @[Math.scala 150:24:@27855.4]
  wire [31:0] x412_sum_1_io_result; // @[Math.scala 150:24:@27855.4]
  wire  x415_sum_1_clock; // @[Math.scala 150:24:@27893.4]
  wire  x415_sum_1_reset; // @[Math.scala 150:24:@27893.4]
  wire [31:0] x415_sum_1_io_a; // @[Math.scala 150:24:@27893.4]
  wire [31:0] x415_sum_1_io_b; // @[Math.scala 150:24:@27893.4]
  wire  x415_sum_1_io_flow; // @[Math.scala 150:24:@27893.4]
  wire [31:0] x415_sum_1_io_result; // @[Math.scala 150:24:@27893.4]
  wire  x418_sum_1_clock; // @[Math.scala 150:24:@27931.4]
  wire  x418_sum_1_reset; // @[Math.scala 150:24:@27931.4]
  wire [31:0] x418_sum_1_io_a; // @[Math.scala 150:24:@27931.4]
  wire [31:0] x418_sum_1_io_b; // @[Math.scala 150:24:@27931.4]
  wire  x418_sum_1_io_flow; // @[Math.scala 150:24:@27931.4]
  wire [31:0] x418_sum_1_io_result; // @[Math.scala 150:24:@27931.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@27946.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@27946.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@27946.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@27946.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@27946.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@27960.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@27960.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@27960.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@27960.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@27960.4]
  wire  x421_sub_1_clock; // @[Math.scala 191:24:@27971.4]
  wire  x421_sub_1_reset; // @[Math.scala 191:24:@27971.4]
  wire [31:0] x421_sub_1_io_a; // @[Math.scala 191:24:@27971.4]
  wire [31:0] x421_sub_1_io_b; // @[Math.scala 191:24:@27971.4]
  wire  x421_sub_1_io_flow; // @[Math.scala 191:24:@27971.4]
  wire [31:0] x421_sub_1_io_result; // @[Math.scala 191:24:@27971.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@27981.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@27981.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@27981.4]
  wire [31:0] RetimeWrapper_30_io_in; // @[package.scala 93:22:@27981.4]
  wire [31:0] RetimeWrapper_30_io_out; // @[package.scala 93:22:@27981.4]
  wire  x240_div_1_clock; // @[Math.scala 327:24:@27995.4]
  wire [31:0] x240_div_1_io_a; // @[Math.scala 327:24:@27995.4]
  wire  x240_div_1_io_flow; // @[Math.scala 327:24:@27995.4]
  wire [31:0] x240_div_1_io_result; // @[Math.scala 327:24:@27995.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@28005.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@28005.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@28005.4]
  wire [31:0] RetimeWrapper_31_io_in; // @[package.scala 93:22:@28005.4]
  wire [31:0] RetimeWrapper_31_io_out; // @[package.scala 93:22:@28005.4]
  wire  x241_sum_1_clock; // @[Math.scala 150:24:@28014.4]
  wire  x241_sum_1_reset; // @[Math.scala 150:24:@28014.4]
  wire [31:0] x241_sum_1_io_a; // @[Math.scala 150:24:@28014.4]
  wire [31:0] x241_sum_1_io_b; // @[Math.scala 150:24:@28014.4]
  wire  x241_sum_1_io_flow; // @[Math.scala 150:24:@28014.4]
  wire [31:0] x241_sum_1_io_result; // @[Math.scala 150:24:@28014.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@28024.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@28024.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@28024.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@28024.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@28024.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@28033.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@28033.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@28033.4]
  wire [31:0] RetimeWrapper_33_io_in; // @[package.scala 93:22:@28033.4]
  wire [31:0] RetimeWrapper_33_io_out; // @[package.scala 93:22:@28033.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@28045.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@28045.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@28045.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@28045.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@28045.4]
  wire  x244_rdcol_1_clock; // @[Math.scala 191:24:@28068.4]
  wire  x244_rdcol_1_reset; // @[Math.scala 191:24:@28068.4]
  wire [31:0] x244_rdcol_1_io_a; // @[Math.scala 191:24:@28068.4]
  wire [31:0] x244_rdcol_1_io_b; // @[Math.scala 191:24:@28068.4]
  wire  x244_rdcol_1_io_flow; // @[Math.scala 191:24:@28068.4]
  wire [31:0] x244_rdcol_1_io_result; // @[Math.scala 191:24:@28068.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@28083.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@28083.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@28083.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@28083.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@28083.4]
  wire  x425_sum_1_clock; // @[Math.scala 150:24:@28128.4]
  wire  x425_sum_1_reset; // @[Math.scala 150:24:@28128.4]
  wire [31:0] x425_sum_1_io_a; // @[Math.scala 150:24:@28128.4]
  wire [31:0] x425_sum_1_io_b; // @[Math.scala 150:24:@28128.4]
  wire  x425_sum_1_io_flow; // @[Math.scala 150:24:@28128.4]
  wire [31:0] x425_sum_1_io_result; // @[Math.scala 150:24:@28128.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@28151.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@28151.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@28151.4]
  wire [31:0] RetimeWrapper_36_io_in; // @[package.scala 93:22:@28151.4]
  wire [31:0] RetimeWrapper_36_io_out; // @[package.scala 93:22:@28151.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@28169.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@28169.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@28169.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@28169.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@28169.4]
  wire  x428_sum_1_clock; // @[Math.scala 150:24:@28182.4]
  wire  x428_sum_1_reset; // @[Math.scala 150:24:@28182.4]
  wire [31:0] x428_sum_1_io_a; // @[Math.scala 150:24:@28182.4]
  wire [31:0] x428_sum_1_io_b; // @[Math.scala 150:24:@28182.4]
  wire  x428_sum_1_io_flow; // @[Math.scala 150:24:@28182.4]
  wire [31:0] x428_sum_1_io_result; // @[Math.scala 150:24:@28182.4]
  wire  x431_sum_1_clock; // @[Math.scala 150:24:@28220.4]
  wire  x431_sum_1_reset; // @[Math.scala 150:24:@28220.4]
  wire [31:0] x431_sum_1_io_a; // @[Math.scala 150:24:@28220.4]
  wire [31:0] x431_sum_1_io_b; // @[Math.scala 150:24:@28220.4]
  wire  x431_sum_1_io_flow; // @[Math.scala 150:24:@28220.4]
  wire [31:0] x431_sum_1_io_result; // @[Math.scala 150:24:@28220.4]
  wire  x434_sum_1_clock; // @[Math.scala 150:24:@28258.4]
  wire  x434_sum_1_reset; // @[Math.scala 150:24:@28258.4]
  wire [31:0] x434_sum_1_io_a; // @[Math.scala 150:24:@28258.4]
  wire [31:0] x434_sum_1_io_b; // @[Math.scala 150:24:@28258.4]
  wire  x434_sum_1_io_flow; // @[Math.scala 150:24:@28258.4]
  wire [31:0] x434_sum_1_io_result; // @[Math.scala 150:24:@28258.4]
  wire  x437_sum_1_clock; // @[Math.scala 150:24:@28296.4]
  wire  x437_sum_1_reset; // @[Math.scala 150:24:@28296.4]
  wire [31:0] x437_sum_1_io_a; // @[Math.scala 150:24:@28296.4]
  wire [31:0] x437_sum_1_io_b; // @[Math.scala 150:24:@28296.4]
  wire  x437_sum_1_io_flow; // @[Math.scala 150:24:@28296.4]
  wire [31:0] x437_sum_1_io_result; // @[Math.scala 150:24:@28296.4]
  wire  x440_sum_1_clock; // @[Math.scala 150:24:@28334.4]
  wire  x440_sum_1_reset; // @[Math.scala 150:24:@28334.4]
  wire [31:0] x440_sum_1_io_a; // @[Math.scala 150:24:@28334.4]
  wire [31:0] x440_sum_1_io_b; // @[Math.scala 150:24:@28334.4]
  wire  x440_sum_1_io_flow; // @[Math.scala 150:24:@28334.4]
  wire [31:0] x440_sum_1_io_result; // @[Math.scala 150:24:@28334.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@28349.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@28349.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@28349.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@28349.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@28349.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@28363.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@28363.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@28363.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@28363.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@28363.4]
  wire  x443_sub_1_clock; // @[Math.scala 191:24:@28374.4]
  wire  x443_sub_1_reset; // @[Math.scala 191:24:@28374.4]
  wire [31:0] x443_sub_1_io_a; // @[Math.scala 191:24:@28374.4]
  wire [31:0] x443_sub_1_io_b; // @[Math.scala 191:24:@28374.4]
  wire  x443_sub_1_io_flow; // @[Math.scala 191:24:@28374.4]
  wire [31:0] x443_sub_1_io_result; // @[Math.scala 191:24:@28374.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@28384.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@28384.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@28384.4]
  wire [31:0] RetimeWrapper_40_io_in; // @[package.scala 93:22:@28384.4]
  wire [31:0] RetimeWrapper_40_io_out; // @[package.scala 93:22:@28384.4]
  wire  x249_div_1_clock; // @[Math.scala 327:24:@28398.4]
  wire [31:0] x249_div_1_io_a; // @[Math.scala 327:24:@28398.4]
  wire  x249_div_1_io_flow; // @[Math.scala 327:24:@28398.4]
  wire [31:0] x249_div_1_io_result; // @[Math.scala 327:24:@28398.4]
  wire  x250_sum_1_clock; // @[Math.scala 150:24:@28408.4]
  wire  x250_sum_1_reset; // @[Math.scala 150:24:@28408.4]
  wire [31:0] x250_sum_1_io_a; // @[Math.scala 150:24:@28408.4]
  wire [31:0] x250_sum_1_io_b; // @[Math.scala 150:24:@28408.4]
  wire  x250_sum_1_io_flow; // @[Math.scala 150:24:@28408.4]
  wire [31:0] x250_sum_1_io_result; // @[Math.scala 150:24:@28408.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@28418.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@28418.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@28418.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@28418.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@28418.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@28427.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@28427.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@28427.4]
  wire [31:0] RetimeWrapper_42_io_in; // @[package.scala 93:22:@28427.4]
  wire [31:0] RetimeWrapper_42_io_out; // @[package.scala 93:22:@28427.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@28439.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@28439.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@28439.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@28439.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@28439.4]
  wire  x253_rdrow_1_clock; // @[Math.scala 191:24:@28462.4]
  wire  x253_rdrow_1_reset; // @[Math.scala 191:24:@28462.4]
  wire [31:0] x253_rdrow_1_io_a; // @[Math.scala 191:24:@28462.4]
  wire [31:0] x253_rdrow_1_io_b; // @[Math.scala 191:24:@28462.4]
  wire  x253_rdrow_1_io_flow; // @[Math.scala 191:24:@28462.4]
  wire [31:0] x253_rdrow_1_io_result; // @[Math.scala 191:24:@28462.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@28488.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@28488.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@28488.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@28488.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@28488.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@28497.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@28497.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@28497.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@28497.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@28497.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@28519.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@28519.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@28519.4]
  wire [31:0] RetimeWrapper_46_io_in; // @[package.scala 93:22:@28519.4]
  wire [31:0] RetimeWrapper_46_io_out; // @[package.scala 93:22:@28519.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@28545.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@28545.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@28545.4]
  wire [31:0] RetimeWrapper_47_io_in; // @[package.scala 93:22:@28545.4]
  wire [31:0] RetimeWrapper_47_io_out; // @[package.scala 93:22:@28545.4]
  wire  x449_sum_1_clock; // @[Math.scala 150:24:@28566.4]
  wire  x449_sum_1_reset; // @[Math.scala 150:24:@28566.4]
  wire [31:0] x449_sum_1_io_a; // @[Math.scala 150:24:@28566.4]
  wire [31:0] x449_sum_1_io_b; // @[Math.scala 150:24:@28566.4]
  wire  x449_sum_1_io_flow; // @[Math.scala 150:24:@28566.4]
  wire [31:0] x449_sum_1_io_result; // @[Math.scala 150:24:@28566.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@28576.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@28576.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@28576.4]
  wire [31:0] RetimeWrapper_48_io_in; // @[package.scala 93:22:@28576.4]
  wire [31:0] RetimeWrapper_48_io_out; // @[package.scala 93:22:@28576.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@28585.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@28585.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@28585.4]
  wire [31:0] RetimeWrapper_49_io_in; // @[package.scala 93:22:@28585.4]
  wire [31:0] RetimeWrapper_49_io_out; // @[package.scala 93:22:@28585.4]
  wire  x261_sum_1_clock; // @[Math.scala 150:24:@28594.4]
  wire  x261_sum_1_reset; // @[Math.scala 150:24:@28594.4]
  wire [31:0] x261_sum_1_io_a; // @[Math.scala 150:24:@28594.4]
  wire [31:0] x261_sum_1_io_b; // @[Math.scala 150:24:@28594.4]
  wire  x261_sum_1_io_flow; // @[Math.scala 150:24:@28594.4]
  wire [31:0] x261_sum_1_io_result; // @[Math.scala 150:24:@28594.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@28604.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@28604.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@28604.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@28604.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@28604.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@28613.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@28613.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@28613.4]
  wire [31:0] RetimeWrapper_51_io_in; // @[package.scala 93:22:@28613.4]
  wire [31:0] RetimeWrapper_51_io_out; // @[package.scala 93:22:@28613.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@28622.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@28622.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@28622.4]
  wire [31:0] RetimeWrapper_52_io_in; // @[package.scala 93:22:@28622.4]
  wire [31:0] RetimeWrapper_52_io_out; // @[package.scala 93:22:@28622.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@28634.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@28634.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@28634.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@28634.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@28634.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@28661.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@28661.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@28661.4]
  wire [31:0] RetimeWrapper_54_io_in; // @[package.scala 93:22:@28661.4]
  wire [31:0] RetimeWrapper_54_io_out; // @[package.scala 93:22:@28661.4]
  wire  x266_sum_1_clock; // @[Math.scala 150:24:@28672.4]
  wire  x266_sum_1_reset; // @[Math.scala 150:24:@28672.4]
  wire [31:0] x266_sum_1_io_a; // @[Math.scala 150:24:@28672.4]
  wire [31:0] x266_sum_1_io_b; // @[Math.scala 150:24:@28672.4]
  wire  x266_sum_1_io_flow; // @[Math.scala 150:24:@28672.4]
  wire [31:0] x266_sum_1_io_result; // @[Math.scala 150:24:@28672.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@28682.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@28682.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@28682.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@28682.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@28682.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@28694.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@28694.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@28694.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@28694.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@28694.4]
  wire  x271_sum_1_clock; // @[Math.scala 150:24:@28721.4]
  wire  x271_sum_1_reset; // @[Math.scala 150:24:@28721.4]
  wire [31:0] x271_sum_1_io_a; // @[Math.scala 150:24:@28721.4]
  wire [31:0] x271_sum_1_io_b; // @[Math.scala 150:24:@28721.4]
  wire  x271_sum_1_io_flow; // @[Math.scala 150:24:@28721.4]
  wire [31:0] x271_sum_1_io_result; // @[Math.scala 150:24:@28721.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@28731.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@28731.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@28731.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@28731.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@28731.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@28743.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@28743.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@28743.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@28743.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@28743.4]
  wire  x274_rdrow_1_clock; // @[Math.scala 191:24:@28766.4]
  wire  x274_rdrow_1_reset; // @[Math.scala 191:24:@28766.4]
  wire [31:0] x274_rdrow_1_io_a; // @[Math.scala 191:24:@28766.4]
  wire [31:0] x274_rdrow_1_io_b; // @[Math.scala 191:24:@28766.4]
  wire  x274_rdrow_1_io_flow; // @[Math.scala 191:24:@28766.4]
  wire [31:0] x274_rdrow_1_io_result; // @[Math.scala 191:24:@28766.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@28792.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@28792.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@28792.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@28792.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@28792.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@28814.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@28814.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@28814.4]
  wire [31:0] RetimeWrapper_60_io_in; // @[package.scala 93:22:@28814.4]
  wire [31:0] RetimeWrapper_60_io_out; // @[package.scala 93:22:@28814.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@28840.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@28840.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@28840.4]
  wire [31:0] RetimeWrapper_61_io_in; // @[package.scala 93:22:@28840.4]
  wire [31:0] RetimeWrapper_61_io_out; // @[package.scala 93:22:@28840.4]
  wire  x454_sum_1_clock; // @[Math.scala 150:24:@28861.4]
  wire  x454_sum_1_reset; // @[Math.scala 150:24:@28861.4]
  wire [31:0] x454_sum_1_io_a; // @[Math.scala 150:24:@28861.4]
  wire [31:0] x454_sum_1_io_b; // @[Math.scala 150:24:@28861.4]
  wire  x454_sum_1_io_flow; // @[Math.scala 150:24:@28861.4]
  wire [31:0] x454_sum_1_io_result; // @[Math.scala 150:24:@28861.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@28871.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@28871.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@28871.4]
  wire [31:0] RetimeWrapper_62_io_in; // @[package.scala 93:22:@28871.4]
  wire [31:0] RetimeWrapper_62_io_out; // @[package.scala 93:22:@28871.4]
  wire  x282_sum_1_clock; // @[Math.scala 150:24:@28880.4]
  wire  x282_sum_1_reset; // @[Math.scala 150:24:@28880.4]
  wire [31:0] x282_sum_1_io_a; // @[Math.scala 150:24:@28880.4]
  wire [31:0] x282_sum_1_io_b; // @[Math.scala 150:24:@28880.4]
  wire  x282_sum_1_io_flow; // @[Math.scala 150:24:@28880.4]
  wire [31:0] x282_sum_1_io_result; // @[Math.scala 150:24:@28880.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@28890.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@28890.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@28890.4]
  wire [31:0] RetimeWrapper_63_io_in; // @[package.scala 93:22:@28890.4]
  wire [31:0] RetimeWrapper_63_io_out; // @[package.scala 93:22:@28890.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@28899.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@28899.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@28899.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@28899.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@28899.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@28908.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@28908.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@28908.4]
  wire [31:0] RetimeWrapper_65_io_in; // @[package.scala 93:22:@28908.4]
  wire [31:0] RetimeWrapper_65_io_out; // @[package.scala 93:22:@28908.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@28920.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@28920.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@28920.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@28920.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@28920.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@28947.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@28947.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@28947.4]
  wire [31:0] RetimeWrapper_67_io_in; // @[package.scala 93:22:@28947.4]
  wire [31:0] RetimeWrapper_67_io_out; // @[package.scala 93:22:@28947.4]
  wire  x287_sum_1_clock; // @[Math.scala 150:24:@28956.4]
  wire  x287_sum_1_reset; // @[Math.scala 150:24:@28956.4]
  wire [31:0] x287_sum_1_io_a; // @[Math.scala 150:24:@28956.4]
  wire [31:0] x287_sum_1_io_b; // @[Math.scala 150:24:@28956.4]
  wire  x287_sum_1_io_flow; // @[Math.scala 150:24:@28956.4]
  wire [31:0] x287_sum_1_io_result; // @[Math.scala 150:24:@28956.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@28966.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@28966.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@28966.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@28966.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@28966.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@28978.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@28978.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@28978.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@28978.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@28978.4]
  wire  x292_sum_1_clock; // @[Math.scala 150:24:@29005.4]
  wire  x292_sum_1_reset; // @[Math.scala 150:24:@29005.4]
  wire [31:0] x292_sum_1_io_a; // @[Math.scala 150:24:@29005.4]
  wire [31:0] x292_sum_1_io_b; // @[Math.scala 150:24:@29005.4]
  wire  x292_sum_1_io_flow; // @[Math.scala 150:24:@29005.4]
  wire [31:0] x292_sum_1_io_result; // @[Math.scala 150:24:@29005.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@29015.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@29015.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@29015.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@29015.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@29015.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@29027.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@29027.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@29027.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@29027.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@29027.4]
  wire  x295_1_clock; // @[Math.scala 262:24:@29050.4]
  wire [31:0] x295_1_io_a; // @[Math.scala 262:24:@29050.4]
  wire [31:0] x295_1_io_b; // @[Math.scala 262:24:@29050.4]
  wire  x295_1_io_flow; // @[Math.scala 262:24:@29050.4]
  wire [31:0] x295_1_io_result; // @[Math.scala 262:24:@29050.4]
  wire  x296_1_clock; // @[Math.scala 262:24:@29062.4]
  wire [31:0] x296_1_io_a; // @[Math.scala 262:24:@29062.4]
  wire [31:0] x296_1_io_b; // @[Math.scala 262:24:@29062.4]
  wire  x296_1_io_flow; // @[Math.scala 262:24:@29062.4]
  wire [31:0] x296_1_io_result; // @[Math.scala 262:24:@29062.4]
  wire  x297_1_clock; // @[Math.scala 262:24:@29074.4]
  wire [31:0] x297_1_io_a; // @[Math.scala 262:24:@29074.4]
  wire [31:0] x297_1_io_b; // @[Math.scala 262:24:@29074.4]
  wire  x297_1_io_flow; // @[Math.scala 262:24:@29074.4]
  wire [31:0] x297_1_io_result; // @[Math.scala 262:24:@29074.4]
  wire  x298_1_clock; // @[Math.scala 262:24:@29086.4]
  wire [31:0] x298_1_io_a; // @[Math.scala 262:24:@29086.4]
  wire [31:0] x298_1_io_b; // @[Math.scala 262:24:@29086.4]
  wire  x298_1_io_flow; // @[Math.scala 262:24:@29086.4]
  wire [31:0] x298_1_io_result; // @[Math.scala 262:24:@29086.4]
  wire  x299_1_clock; // @[Math.scala 262:24:@29098.4]
  wire [31:0] x299_1_io_a; // @[Math.scala 262:24:@29098.4]
  wire [31:0] x299_1_io_b; // @[Math.scala 262:24:@29098.4]
  wire  x299_1_io_flow; // @[Math.scala 262:24:@29098.4]
  wire [31:0] x299_1_io_result; // @[Math.scala 262:24:@29098.4]
  wire  x300_1_clock; // @[Math.scala 262:24:@29112.4]
  wire [31:0] x300_1_io_a; // @[Math.scala 262:24:@29112.4]
  wire [31:0] x300_1_io_b; // @[Math.scala 262:24:@29112.4]
  wire  x300_1_io_flow; // @[Math.scala 262:24:@29112.4]
  wire [31:0] x300_1_io_result; // @[Math.scala 262:24:@29112.4]
  wire  x301_1_clock; // @[Math.scala 262:24:@29124.4]
  wire [31:0] x301_1_io_a; // @[Math.scala 262:24:@29124.4]
  wire [31:0] x301_1_io_b; // @[Math.scala 262:24:@29124.4]
  wire  x301_1_io_flow; // @[Math.scala 262:24:@29124.4]
  wire [31:0] x301_1_io_result; // @[Math.scala 262:24:@29124.4]
  wire  x302_1_clock; // @[Math.scala 262:24:@29136.4]
  wire [31:0] x302_1_io_a; // @[Math.scala 262:24:@29136.4]
  wire [31:0] x302_1_io_b; // @[Math.scala 262:24:@29136.4]
  wire  x302_1_io_flow; // @[Math.scala 262:24:@29136.4]
  wire [31:0] x302_1_io_result; // @[Math.scala 262:24:@29136.4]
  wire  x303_1_clock; // @[Math.scala 262:24:@29148.4]
  wire [31:0] x303_1_io_a; // @[Math.scala 262:24:@29148.4]
  wire [31:0] x303_1_io_b; // @[Math.scala 262:24:@29148.4]
  wire  x303_1_io_flow; // @[Math.scala 262:24:@29148.4]
  wire [31:0] x303_1_io_result; // @[Math.scala 262:24:@29148.4]
  wire  x304_x3_1_clock; // @[Math.scala 150:24:@29158.4]
  wire  x304_x3_1_reset; // @[Math.scala 150:24:@29158.4]
  wire [31:0] x304_x3_1_io_a; // @[Math.scala 150:24:@29158.4]
  wire [31:0] x304_x3_1_io_b; // @[Math.scala 150:24:@29158.4]
  wire  x304_x3_1_io_flow; // @[Math.scala 150:24:@29158.4]
  wire [31:0] x304_x3_1_io_result; // @[Math.scala 150:24:@29158.4]
  wire  x305_x4_1_clock; // @[Math.scala 150:24:@29168.4]
  wire  x305_x4_1_reset; // @[Math.scala 150:24:@29168.4]
  wire [31:0] x305_x4_1_io_a; // @[Math.scala 150:24:@29168.4]
  wire [31:0] x305_x4_1_io_b; // @[Math.scala 150:24:@29168.4]
  wire  x305_x4_1_io_flow; // @[Math.scala 150:24:@29168.4]
  wire [31:0] x305_x4_1_io_result; // @[Math.scala 150:24:@29168.4]
  wire  x306_x3_1_clock; // @[Math.scala 150:24:@29178.4]
  wire  x306_x3_1_reset; // @[Math.scala 150:24:@29178.4]
  wire [31:0] x306_x3_1_io_a; // @[Math.scala 150:24:@29178.4]
  wire [31:0] x306_x3_1_io_b; // @[Math.scala 150:24:@29178.4]
  wire  x306_x3_1_io_flow; // @[Math.scala 150:24:@29178.4]
  wire [31:0] x306_x3_1_io_result; // @[Math.scala 150:24:@29178.4]
  wire  x307_x4_1_clock; // @[Math.scala 150:24:@29188.4]
  wire  x307_x4_1_reset; // @[Math.scala 150:24:@29188.4]
  wire [31:0] x307_x4_1_io_a; // @[Math.scala 150:24:@29188.4]
  wire [31:0] x307_x4_1_io_b; // @[Math.scala 150:24:@29188.4]
  wire  x307_x4_1_io_flow; // @[Math.scala 150:24:@29188.4]
  wire [31:0] x307_x4_1_io_result; // @[Math.scala 150:24:@29188.4]
  wire  x308_x3_1_clock; // @[Math.scala 150:24:@29198.4]
  wire  x308_x3_1_reset; // @[Math.scala 150:24:@29198.4]
  wire [31:0] x308_x3_1_io_a; // @[Math.scala 150:24:@29198.4]
  wire [31:0] x308_x3_1_io_b; // @[Math.scala 150:24:@29198.4]
  wire  x308_x3_1_io_flow; // @[Math.scala 150:24:@29198.4]
  wire [31:0] x308_x3_1_io_result; // @[Math.scala 150:24:@29198.4]
  wire  x309_x4_1_clock; // @[Math.scala 150:24:@29208.4]
  wire  x309_x4_1_reset; // @[Math.scala 150:24:@29208.4]
  wire [31:0] x309_x4_1_io_a; // @[Math.scala 150:24:@29208.4]
  wire [31:0] x309_x4_1_io_b; // @[Math.scala 150:24:@29208.4]
  wire  x309_x4_1_io_flow; // @[Math.scala 150:24:@29208.4]
  wire [31:0] x309_x4_1_io_result; // @[Math.scala 150:24:@29208.4]
  wire  x310_x3_1_clock; // @[Math.scala 150:24:@29218.4]
  wire  x310_x3_1_reset; // @[Math.scala 150:24:@29218.4]
  wire [31:0] x310_x3_1_io_a; // @[Math.scala 150:24:@29218.4]
  wire [31:0] x310_x3_1_io_b; // @[Math.scala 150:24:@29218.4]
  wire  x310_x3_1_io_flow; // @[Math.scala 150:24:@29218.4]
  wire [31:0] x310_x3_1_io_result; // @[Math.scala 150:24:@29218.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@29228.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@29228.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@29228.4]
  wire [31:0] RetimeWrapper_72_io_in; // @[package.scala 93:22:@29228.4]
  wire [31:0] RetimeWrapper_72_io_out; // @[package.scala 93:22:@29228.4]
  wire  x311_sum_1_clock; // @[Math.scala 150:24:@29237.4]
  wire  x311_sum_1_reset; // @[Math.scala 150:24:@29237.4]
  wire [31:0] x311_sum_1_io_a; // @[Math.scala 150:24:@29237.4]
  wire [31:0] x311_sum_1_io_b; // @[Math.scala 150:24:@29237.4]
  wire  x311_sum_1_io_flow; // @[Math.scala 150:24:@29237.4]
  wire [31:0] x311_sum_1_io_result; // @[Math.scala 150:24:@29237.4]
  wire [31:0] x312_1_io_b; // @[Math.scala 720:24:@29247.4]
  wire [31:0] x312_1_io_result; // @[Math.scala 720:24:@29247.4]
  wire  x313_mul_1_clock; // @[Math.scala 262:24:@29258.4]
  wire [31:0] x313_mul_1_io_a; // @[Math.scala 262:24:@29258.4]
  wire  x313_mul_1_io_flow; // @[Math.scala 262:24:@29258.4]
  wire [31:0] x313_mul_1_io_result; // @[Math.scala 262:24:@29258.4]
  wire [31:0] x314_1_io_b; // @[Math.scala 720:24:@29268.4]
  wire [31:0] x314_1_io_result; // @[Math.scala 720:24:@29268.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@29281.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@29281.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@29281.4]
  wire [31:0] RetimeWrapper_73_io_in; // @[package.scala 93:22:@29281.4]
  wire [31:0] RetimeWrapper_73_io_out; // @[package.scala 93:22:@29281.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@29290.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@29290.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@29290.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@29290.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@29290.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@29299.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@29299.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@29299.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@29299.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@29299.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@29308.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@29308.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@29308.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@29308.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@29308.4]
  wire  b213; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 62:18:@26966.4]
  wire  b214; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 63:18:@26967.4]
  wire  _T_205; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 67:30:@26969.4]
  wire  _T_206; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 67:37:@26970.4]
  wire  _T_210; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 69:76:@26975.4]
  wire  _T_211; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 69:62:@26976.4]
  wire  _T_213; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 69:101:@26977.4]
  wire [31:0] b211_number; // @[Math.scala 723:22:@26951.4 Math.scala 724:14:@26952.4]
  wire [31:0] _T_241; // @[Math.scala 406:49:@27067.4]
  wire [31:0] _T_243; // @[Math.scala 406:56:@27069.4]
  wire [31:0] _T_244; // @[Math.scala 406:56:@27070.4]
  wire [31:0] x374_number; // @[implicits.scala 133:21:@27071.4]
  wire [31:0] _T_254; // @[Math.scala 406:49:@27080.4]
  wire [31:0] _T_256; // @[Math.scala 406:56:@27082.4]
  wire [31:0] _T_257; // @[Math.scala 406:56:@27083.4]
  wire [31:0] b212_number; // @[Math.scala 723:22:@26963.4 Math.scala 724:14:@26964.4]
  wire  _T_261; // @[FixedPoint.scala 50:25:@27089.4]
  wire [15:0] _T_265; // @[Bitwise.scala 72:12:@27091.4]
  wire [15:0] _T_266; // @[FixedPoint.scala 18:52:@27092.4]
  wire  _T_272; // @[Math.scala 451:55:@27094.4]
  wire [15:0] _T_273; // @[FixedPoint.scala 18:52:@27095.4]
  wire  _T_279; // @[Math.scala 451:110:@27097.4]
  wire  _T_280; // @[Math.scala 451:94:@27098.4]
  wire [31:0] _T_282; // @[Cat.scala 30:58:@27100.4]
  wire [31:0] _T_292; // @[Math.scala 406:49:@27108.4]
  wire [31:0] _T_294; // @[Math.scala 406:56:@27110.4]
  wire [31:0] _T_295; // @[Math.scala 406:56:@27111.4]
  wire [31:0] x378_sum_number; // @[Math.scala 154:22:@27122.4 Math.scala 155:14:@27123.4]
  wire  _T_302; // @[FixedPoint.scala 50:25:@27127.4]
  wire [7:0] _T_306; // @[Bitwise.scala 72:12:@27129.4]
  wire [23:0] _T_307; // @[FixedPoint.scala 18:52:@27130.4]
  wire  _T_313; // @[Math.scala 451:55:@27132.4]
  wire [7:0] _T_314; // @[FixedPoint.scala 18:52:@27133.4]
  wire  _T_320; // @[Math.scala 451:110:@27135.4]
  wire  _T_321; // @[Math.scala 451:94:@27136.4]
  wire [31:0] _T_323; // @[Cat.scala 30:58:@27138.4]
  wire [31:0] _T_333; // @[Math.scala 406:49:@27146.4]
  wire [31:0] _T_335; // @[Math.scala 406:56:@27148.4]
  wire [31:0] _T_336; // @[Math.scala 406:56:@27149.4]
  wire [31:0] x381_sum_number; // @[Math.scala 154:22:@27160.4 Math.scala 155:14:@27161.4]
  wire  _T_343; // @[FixedPoint.scala 50:25:@27165.4]
  wire [3:0] _T_347; // @[Bitwise.scala 72:12:@27167.4]
  wire [27:0] _T_348; // @[FixedPoint.scala 18:52:@27168.4]
  wire  _T_354; // @[Math.scala 451:55:@27170.4]
  wire [3:0] _T_355; // @[FixedPoint.scala 18:52:@27171.4]
  wire  _T_361; // @[Math.scala 451:110:@27173.4]
  wire  _T_362; // @[Math.scala 451:94:@27174.4]
  wire [31:0] _T_364; // @[Cat.scala 30:58:@27176.4]
  wire [31:0] _T_374; // @[Math.scala 406:49:@27184.4]
  wire [31:0] _T_376; // @[Math.scala 406:56:@27186.4]
  wire [31:0] _T_377; // @[Math.scala 406:56:@27187.4]
  wire [31:0] x384_sum_number; // @[Math.scala 154:22:@27198.4 Math.scala 155:14:@27199.4]
  wire  _T_384; // @[FixedPoint.scala 50:25:@27203.4]
  wire [1:0] _T_388; // @[Bitwise.scala 72:12:@27205.4]
  wire [29:0] _T_389; // @[FixedPoint.scala 18:52:@27206.4]
  wire  _T_395; // @[Math.scala 451:55:@27208.4]
  wire [1:0] _T_396; // @[FixedPoint.scala 18:52:@27209.4]
  wire  _T_402; // @[Math.scala 451:110:@27211.4]
  wire  _T_403; // @[Math.scala 451:94:@27212.4]
  wire [31:0] _T_405; // @[Cat.scala 30:58:@27214.4]
  wire [31:0] _T_415; // @[Math.scala 406:49:@27222.4]
  wire [31:0] _T_417; // @[Math.scala 406:56:@27224.4]
  wire [31:0] _T_418; // @[Math.scala 406:56:@27225.4]
  wire [31:0] x387_sum_number; // @[Math.scala 154:22:@27236.4 Math.scala 155:14:@27237.4]
  wire  _T_425; // @[FixedPoint.scala 50:25:@27241.4]
  wire [1:0] _T_429; // @[Bitwise.scala 72:12:@27243.4]
  wire [29:0] _T_430; // @[FixedPoint.scala 18:52:@27244.4]
  wire  _T_436; // @[Math.scala 451:55:@27246.4]
  wire [1:0] _T_437; // @[FixedPoint.scala 18:52:@27247.4]
  wire  _T_443; // @[Math.scala 451:110:@27249.4]
  wire  _T_444; // @[Math.scala 451:94:@27250.4]
  wire [31:0] _T_448; // @[package.scala 96:25:@27258.4 package.scala 96:25:@27259.4]
  wire [31:0] _T_458; // @[Math.scala 406:49:@27267.4]
  wire [31:0] _T_460; // @[Math.scala 406:56:@27269.4]
  wire [31:0] _T_461; // @[Math.scala 406:56:@27270.4]
  wire [31:0] _T_465; // @[package.scala 96:25:@27278.4]
  wire [31:0] x390_sum_number; // @[Math.scala 154:22:@27290.4 Math.scala 155:14:@27291.4]
  wire  _T_472; // @[FixedPoint.scala 50:25:@27295.4]
  wire [1:0] _T_476; // @[Bitwise.scala 72:12:@27297.4]
  wire [29:0] _T_477; // @[FixedPoint.scala 18:52:@27298.4]
  wire  _T_483; // @[Math.scala 451:55:@27300.4]
  wire [1:0] _T_484; // @[FixedPoint.scala 18:52:@27301.4]
  wire  _T_490; // @[Math.scala 451:110:@27303.4]
  wire  _T_491; // @[Math.scala 451:94:@27304.4]
  wire [31:0] _T_493; // @[Cat.scala 30:58:@27306.4]
  wire [31:0] _T_503; // @[Math.scala 406:49:@27314.4]
  wire [31:0] _T_505; // @[Math.scala 406:56:@27316.4]
  wire [31:0] _T_506; // @[Math.scala 406:56:@27317.4]
  wire [31:0] x393_sum_number; // @[Math.scala 154:22:@27328.4 Math.scala 155:14:@27329.4]
  wire [31:0] _T_516; // @[Math.scala 476:37:@27334.4]
  wire  x462_x394_D1; // @[package.scala 96:25:@27372.4 package.scala 96:25:@27373.4]
  wire [31:0] x463_x393_sum_D1_number; // @[package.scala 96:25:@27381.4 package.scala 96:25:@27382.4]
  wire [31:0] x396_sub_number; // @[Math.scala 195:22:@27354.4 Math.scala 196:14:@27355.4]
  wire  _T_547; // @[FixedPoint.scala 50:25:@27389.4]
  wire [1:0] _T_551; // @[Bitwise.scala 72:12:@27391.4]
  wire [29:0] _T_552; // @[FixedPoint.scala 18:52:@27392.4]
  wire  _T_558; // @[Math.scala 451:55:@27394.4]
  wire [1:0] _T_559; // @[FixedPoint.scala 18:52:@27395.4]
  wire  _T_565; // @[Math.scala 451:110:@27397.4]
  wire  _T_566; // @[Math.scala 451:94:@27398.4]
  wire [31:0] _T_568; // @[Cat.scala 30:58:@27400.4]
  wire [31:0] x223_1_number; // @[Math.scala 454:20:@27401.4]
  wire [40:0] _GEN_0; // @[Math.scala 461:32:@27406.4]
  wire [40:0] _T_573; // @[Math.scala 461:32:@27406.4]
  wire [38:0] _GEN_1; // @[Math.scala 461:32:@27411.4]
  wire [38:0] _T_576; // @[Math.scala 461:32:@27411.4]
  wire  _T_609; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 163:101:@27500.4]
  wire  _T_613; // @[package.scala 96:25:@27508.4 package.scala 96:25:@27509.4]
  wire  _T_615; // @[implicits.scala 55:10:@27510.4]
  wire  _T_616; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 163:118:@27511.4]
  wire  _T_618; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 163:207:@27513.4]
  wire  _T_619; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 163:226:@27514.4]
  wire  x468_b213_D21; // @[package.scala 96:25:@27488.4 package.scala 96:25:@27489.4]
  wire  _T_620; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 163:252:@27515.4]
  wire  x469_b214_D21; // @[package.scala 96:25:@27497.4 package.scala 96:25:@27498.4]
  wire [31:0] x470_b211_D23_number; // @[package.scala 96:25:@27529.4 package.scala 96:25:@27530.4]
  wire [31:0] _T_630; // @[Math.scala 476:37:@27535.4]
  wire [31:0] x471_b212_D23_number; // @[package.scala 96:25:@27552.4 package.scala 96:25:@27553.4]
  wire [31:0] _T_645; // @[Math.scala 476:37:@27560.4]
  wire  x229; // @[package.scala 96:25:@27543.4 package.scala 96:25:@27544.4]
  wire  x230; // @[package.scala 96:25:@27568.4 package.scala 96:25:@27569.4]
  wire  x231; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 182:59:@27572.4]
  wire  _T_683; // @[package.scala 96:25:@27640.4 package.scala 96:25:@27641.4]
  wire  _T_685; // @[implicits.scala 55:10:@27642.4]
  wire  _T_686; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 201:194:@27643.4]
  wire  x477_x232_D21; // @[package.scala 96:25:@27628.4 package.scala 96:25:@27629.4]
  wire  _T_687; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 201:283:@27644.4]
  wire  x474_b213_D45; // @[package.scala 96:25:@27601.4 package.scala 96:25:@27602.4]
  wire  _T_688; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 201:291:@27645.4]
  wire  x476_b214_D45; // @[package.scala 96:25:@27619.4 package.scala 96:25:@27620.4]
  wire [31:0] x235_rdcol_number; // @[Math.scala 195:22:@27664.4 Math.scala 196:14:@27665.4]
  wire [31:0] _T_703; // @[Math.scala 476:37:@27670.4]
  wire  x478_x229_D1; // @[package.scala 96:25:@27687.4 package.scala 96:25:@27688.4]
  wire  x236; // @[package.scala 96:25:@27678.4 package.scala 96:25:@27679.4]
  wire  x237; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 211:24:@27691.4]
  wire  _T_717; // @[FixedPoint.scala 50:25:@27698.4]
  wire [15:0] _T_721; // @[Bitwise.scala 72:12:@27700.4]
  wire [15:0] _T_722; // @[FixedPoint.scala 18:52:@27701.4]
  wire  _T_728; // @[Math.scala 451:55:@27703.4]
  wire [15:0] _T_729; // @[FixedPoint.scala 18:52:@27704.4]
  wire  _T_735; // @[Math.scala 451:110:@27706.4]
  wire  _T_736; // @[Math.scala 451:94:@27707.4]
  wire [31:0] _T_738; // @[Cat.scala 30:58:@27709.4]
  wire [31:0] _T_750; // @[Math.scala 406:56:@27719.4]
  wire [31:0] _T_751; // @[Math.scala 406:56:@27720.4]
  wire [31:0] x403_sum_number; // @[Math.scala 154:22:@27731.4 Math.scala 155:14:@27732.4]
  wire  _T_758; // @[FixedPoint.scala 50:25:@27736.4]
  wire [7:0] _T_762; // @[Bitwise.scala 72:12:@27738.4]
  wire [23:0] _T_763; // @[FixedPoint.scala 18:52:@27739.4]
  wire  _T_769; // @[Math.scala 451:55:@27741.4]
  wire [7:0] _T_770; // @[FixedPoint.scala 18:52:@27742.4]
  wire  _T_776; // @[Math.scala 451:110:@27744.4]
  wire  _T_777; // @[Math.scala 451:94:@27745.4]
  wire [31:0] _T_781; // @[package.scala 96:25:@27753.4 package.scala 96:25:@27754.4]
  wire [31:0] _T_791; // @[Math.scala 406:49:@27762.4]
  wire [31:0] _T_793; // @[Math.scala 406:56:@27764.4]
  wire [31:0] _T_794; // @[Math.scala 406:56:@27765.4]
  wire [31:0] _T_798; // @[package.scala 96:25:@27773.4]
  wire [31:0] x406_sum_number; // @[Math.scala 154:22:@27785.4 Math.scala 155:14:@27786.4]
  wire  _T_805; // @[FixedPoint.scala 50:25:@27790.4]
  wire [3:0] _T_809; // @[Bitwise.scala 72:12:@27792.4]
  wire [27:0] _T_810; // @[FixedPoint.scala 18:52:@27793.4]
  wire  _T_816; // @[Math.scala 451:55:@27795.4]
  wire [3:0] _T_817; // @[FixedPoint.scala 18:52:@27796.4]
  wire  _T_823; // @[Math.scala 451:110:@27798.4]
  wire  _T_824; // @[Math.scala 451:94:@27799.4]
  wire [31:0] _T_826; // @[Cat.scala 30:58:@27801.4]
  wire [31:0] _T_836; // @[Math.scala 406:49:@27809.4]
  wire [31:0] _T_838; // @[Math.scala 406:56:@27811.4]
  wire [31:0] _T_839; // @[Math.scala 406:56:@27812.4]
  wire [31:0] x409_sum_number; // @[Math.scala 154:22:@27823.4 Math.scala 155:14:@27824.4]
  wire  _T_846; // @[FixedPoint.scala 50:25:@27828.4]
  wire [1:0] _T_850; // @[Bitwise.scala 72:12:@27830.4]
  wire [29:0] _T_851; // @[FixedPoint.scala 18:52:@27831.4]
  wire  _T_857; // @[Math.scala 451:55:@27833.4]
  wire [1:0] _T_858; // @[FixedPoint.scala 18:52:@27834.4]
  wire  _T_864; // @[Math.scala 451:110:@27836.4]
  wire  _T_865; // @[Math.scala 451:94:@27837.4]
  wire [31:0] _T_867; // @[Cat.scala 30:58:@27839.4]
  wire [31:0] _T_877; // @[Math.scala 406:49:@27847.4]
  wire [31:0] _T_879; // @[Math.scala 406:56:@27849.4]
  wire [31:0] _T_880; // @[Math.scala 406:56:@27850.4]
  wire [31:0] x412_sum_number; // @[Math.scala 154:22:@27861.4 Math.scala 155:14:@27862.4]
  wire  _T_887; // @[FixedPoint.scala 50:25:@27866.4]
  wire [1:0] _T_891; // @[Bitwise.scala 72:12:@27868.4]
  wire [29:0] _T_892; // @[FixedPoint.scala 18:52:@27869.4]
  wire  _T_898; // @[Math.scala 451:55:@27871.4]
  wire [1:0] _T_899; // @[FixedPoint.scala 18:52:@27872.4]
  wire  _T_905; // @[Math.scala 451:110:@27874.4]
  wire  _T_906; // @[Math.scala 451:94:@27875.4]
  wire [31:0] _T_908; // @[Cat.scala 30:58:@27877.4]
  wire [31:0] _T_918; // @[Math.scala 406:49:@27885.4]
  wire [31:0] _T_920; // @[Math.scala 406:56:@27887.4]
  wire [31:0] _T_921; // @[Math.scala 406:56:@27888.4]
  wire [31:0] x415_sum_number; // @[Math.scala 154:22:@27899.4 Math.scala 155:14:@27900.4]
  wire  _T_928; // @[FixedPoint.scala 50:25:@27904.4]
  wire [1:0] _T_932; // @[Bitwise.scala 72:12:@27906.4]
  wire [29:0] _T_933; // @[FixedPoint.scala 18:52:@27907.4]
  wire  _T_939; // @[Math.scala 451:55:@27909.4]
  wire [1:0] _T_940; // @[FixedPoint.scala 18:52:@27910.4]
  wire  _T_946; // @[Math.scala 451:110:@27912.4]
  wire  _T_947; // @[Math.scala 451:94:@27913.4]
  wire [31:0] _T_949; // @[Cat.scala 30:58:@27915.4]
  wire [31:0] _T_959; // @[Math.scala 406:49:@27923.4]
  wire [31:0] _T_961; // @[Math.scala 406:56:@27925.4]
  wire [31:0] _T_962; // @[Math.scala 406:56:@27926.4]
  wire [31:0] x418_sum_number; // @[Math.scala 154:22:@27937.4 Math.scala 155:14:@27938.4]
  wire [31:0] _T_972; // @[Math.scala 476:37:@27943.4]
  wire  x419; // @[package.scala 96:25:@27951.4 package.scala 96:25:@27952.4]
  wire [31:0] x479_x418_sum_D1_number; // @[package.scala 96:25:@27986.4 package.scala 96:25:@27987.4]
  wire [31:0] x421_sub_number; // @[Math.scala 195:22:@27977.4 Math.scala 196:14:@27978.4]
  wire  _T_1029; // @[package.scala 96:25:@28050.4 package.scala 96:25:@28051.4]
  wire  _T_1031; // @[implicits.scala 55:10:@28052.4]
  wire  _T_1032; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 274:194:@28053.4]
  wire  x481_x238_D20; // @[package.scala 96:25:@28029.4 package.scala 96:25:@28030.4]
  wire  _T_1033; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 274:283:@28054.4]
  wire  _T_1034; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 274:291:@28055.4]
  wire [31:0] x244_rdcol_number; // @[Math.scala 195:22:@28074.4 Math.scala 196:14:@28075.4]
  wire [31:0] _T_1049; // @[Math.scala 476:37:@28080.4]
  wire  x245; // @[package.scala 96:25:@28088.4 package.scala 96:25:@28089.4]
  wire  x246; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 288:59:@28092.4]
  wire  _T_1062; // @[FixedPoint.scala 50:25:@28101.4]
  wire [15:0] _T_1066; // @[Bitwise.scala 72:12:@28103.4]
  wire [15:0] _T_1067; // @[FixedPoint.scala 18:52:@28104.4]
  wire  _T_1073; // @[Math.scala 451:55:@28106.4]
  wire [15:0] _T_1074; // @[FixedPoint.scala 18:52:@28107.4]
  wire  _T_1080; // @[Math.scala 451:110:@28109.4]
  wire  _T_1081; // @[Math.scala 451:94:@28110.4]
  wire [31:0] _T_1083; // @[Cat.scala 30:58:@28112.4]
  wire [31:0] _T_1095; // @[Math.scala 406:56:@28122.4]
  wire [31:0] _T_1096; // @[Math.scala 406:56:@28123.4]
  wire [31:0] x425_sum_number; // @[Math.scala 154:22:@28134.4 Math.scala 155:14:@28135.4]
  wire  _T_1103; // @[FixedPoint.scala 50:25:@28139.4]
  wire [7:0] _T_1107; // @[Bitwise.scala 72:12:@28141.4]
  wire [23:0] _T_1108; // @[FixedPoint.scala 18:52:@28142.4]
  wire  _T_1114; // @[Math.scala 451:55:@28144.4]
  wire [7:0] _T_1115; // @[FixedPoint.scala 18:52:@28145.4]
  wire  _T_1121; // @[Math.scala 451:110:@28147.4]
  wire  _T_1122; // @[Math.scala 451:94:@28148.4]
  wire [31:0] _T_1126; // @[package.scala 96:25:@28156.4 package.scala 96:25:@28157.4]
  wire [31:0] _T_1136; // @[Math.scala 406:49:@28165.4]
  wire [31:0] _T_1138; // @[Math.scala 406:56:@28167.4]
  wire [31:0] _T_1139; // @[Math.scala 406:56:@28168.4]
  wire [31:0] _T_1143; // @[package.scala 96:25:@28176.4]
  wire [31:0] x428_sum_number; // @[Math.scala 154:22:@28188.4 Math.scala 155:14:@28189.4]
  wire  _T_1150; // @[FixedPoint.scala 50:25:@28193.4]
  wire [3:0] _T_1154; // @[Bitwise.scala 72:12:@28195.4]
  wire [27:0] _T_1155; // @[FixedPoint.scala 18:52:@28196.4]
  wire  _T_1161; // @[Math.scala 451:55:@28198.4]
  wire [3:0] _T_1162; // @[FixedPoint.scala 18:52:@28199.4]
  wire  _T_1168; // @[Math.scala 451:110:@28201.4]
  wire  _T_1169; // @[Math.scala 451:94:@28202.4]
  wire [31:0] _T_1171; // @[Cat.scala 30:58:@28204.4]
  wire [31:0] _T_1181; // @[Math.scala 406:49:@28212.4]
  wire [31:0] _T_1183; // @[Math.scala 406:56:@28214.4]
  wire [31:0] _T_1184; // @[Math.scala 406:56:@28215.4]
  wire [31:0] x431_sum_number; // @[Math.scala 154:22:@28226.4 Math.scala 155:14:@28227.4]
  wire  _T_1191; // @[FixedPoint.scala 50:25:@28231.4]
  wire [1:0] _T_1195; // @[Bitwise.scala 72:12:@28233.4]
  wire [29:0] _T_1196; // @[FixedPoint.scala 18:52:@28234.4]
  wire  _T_1202; // @[Math.scala 451:55:@28236.4]
  wire [1:0] _T_1203; // @[FixedPoint.scala 18:52:@28237.4]
  wire  _T_1209; // @[Math.scala 451:110:@28239.4]
  wire  _T_1210; // @[Math.scala 451:94:@28240.4]
  wire [31:0] _T_1212; // @[Cat.scala 30:58:@28242.4]
  wire [31:0] _T_1222; // @[Math.scala 406:49:@28250.4]
  wire [31:0] _T_1224; // @[Math.scala 406:56:@28252.4]
  wire [31:0] _T_1225; // @[Math.scala 406:56:@28253.4]
  wire [31:0] x434_sum_number; // @[Math.scala 154:22:@28264.4 Math.scala 155:14:@28265.4]
  wire  _T_1232; // @[FixedPoint.scala 50:25:@28269.4]
  wire [1:0] _T_1236; // @[Bitwise.scala 72:12:@28271.4]
  wire [29:0] _T_1237; // @[FixedPoint.scala 18:52:@28272.4]
  wire  _T_1243; // @[Math.scala 451:55:@28274.4]
  wire [1:0] _T_1244; // @[FixedPoint.scala 18:52:@28275.4]
  wire  _T_1250; // @[Math.scala 451:110:@28277.4]
  wire  _T_1251; // @[Math.scala 451:94:@28278.4]
  wire [31:0] _T_1253; // @[Cat.scala 30:58:@28280.4]
  wire [31:0] _T_1263; // @[Math.scala 406:49:@28288.4]
  wire [31:0] _T_1265; // @[Math.scala 406:56:@28290.4]
  wire [31:0] _T_1266; // @[Math.scala 406:56:@28291.4]
  wire [31:0] x437_sum_number; // @[Math.scala 154:22:@28302.4 Math.scala 155:14:@28303.4]
  wire  _T_1273; // @[FixedPoint.scala 50:25:@28307.4]
  wire [1:0] _T_1277; // @[Bitwise.scala 72:12:@28309.4]
  wire [29:0] _T_1278; // @[FixedPoint.scala 18:52:@28310.4]
  wire  _T_1284; // @[Math.scala 451:55:@28312.4]
  wire [1:0] _T_1285; // @[FixedPoint.scala 18:52:@28313.4]
  wire  _T_1291; // @[Math.scala 451:110:@28315.4]
  wire  _T_1292; // @[Math.scala 451:94:@28316.4]
  wire [31:0] _T_1294; // @[Cat.scala 30:58:@28318.4]
  wire [31:0] _T_1304; // @[Math.scala 406:49:@28326.4]
  wire [31:0] _T_1306; // @[Math.scala 406:56:@28328.4]
  wire [31:0] _T_1307; // @[Math.scala 406:56:@28329.4]
  wire [31:0] x440_sum_number; // @[Math.scala 154:22:@28340.4 Math.scala 155:14:@28341.4]
  wire [31:0] _T_1317; // @[Math.scala 476:37:@28346.4]
  wire  x441; // @[package.scala 96:25:@28354.4 package.scala 96:25:@28355.4]
  wire [31:0] x483_x440_sum_D1_number; // @[package.scala 96:25:@28389.4 package.scala 96:25:@28390.4]
  wire [31:0] x443_sub_number; // @[Math.scala 195:22:@28380.4 Math.scala 196:14:@28381.4]
  wire  _T_1371; // @[package.scala 96:25:@28444.4 package.scala 96:25:@28445.4]
  wire  _T_1373; // @[implicits.scala 55:10:@28446.4]
  wire  _T_1374; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 351:194:@28447.4]
  wire  x484_x247_D20; // @[package.scala 96:25:@28423.4 package.scala 96:25:@28424.4]
  wire  _T_1375; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 351:283:@28448.4]
  wire  _T_1376; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 351:291:@28449.4]
  wire [31:0] x253_rdrow_number; // @[Math.scala 195:22:@28468.4 Math.scala 196:14:@28469.4]
  wire [31:0] _T_1393; // @[Math.scala 406:49:@28475.4]
  wire [31:0] _T_1395; // @[Math.scala 406:56:@28477.4]
  wire [31:0] _T_1396; // @[Math.scala 406:56:@28478.4]
  wire [31:0] x445_number; // @[implicits.scala 133:21:@28479.4]
  wire  x255; // @[package.scala 96:25:@28493.4 package.scala 96:25:@28494.4]
  wire  x486_x230_D1; // @[package.scala 96:25:@28502.4 package.scala 96:25:@28503.4]
  wire  x256; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 363:24:@28506.4]
  wire [31:0] _T_1422; // @[Math.scala 406:49:@28515.4]
  wire [31:0] _T_1424; // @[Math.scala 406:56:@28517.4]
  wire [31:0] _T_1425; // @[Math.scala 406:56:@28518.4]
  wire [31:0] _T_1429; // @[package.scala 96:25:@28526.4]
  wire  _T_1433; // @[FixedPoint.scala 50:25:@28533.4]
  wire [1:0] _T_1437; // @[Bitwise.scala 72:12:@28535.4]
  wire [29:0] _T_1438; // @[FixedPoint.scala 18:52:@28536.4]
  wire  _T_1444; // @[Math.scala 451:55:@28538.4]
  wire [1:0] _T_1445; // @[FixedPoint.scala 18:52:@28539.4]
  wire  _T_1451; // @[Math.scala 451:110:@28541.4]
  wire  _T_1452; // @[Math.scala 451:94:@28542.4]
  wire [31:0] _T_1456; // @[package.scala 96:25:@28550.4 package.scala 96:25:@28551.4]
  wire [31:0] x259_1_number; // @[Math.scala 454:20:@28552.4]
  wire [40:0] _GEN_2; // @[Math.scala 461:32:@28557.4]
  wire [40:0] _T_1461; // @[Math.scala 461:32:@28557.4]
  wire [38:0] _GEN_3; // @[Math.scala 461:32:@28562.4]
  wire [38:0] _T_1464; // @[Math.scala 461:32:@28562.4]
  wire  _T_1497; // @[package.scala 96:25:@28639.4 package.scala 96:25:@28640.4]
  wire  _T_1499; // @[implicits.scala 55:10:@28641.4]
  wire  _T_1500; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 392:194:@28642.4]
  wire  x489_x257_D20; // @[package.scala 96:25:@28609.4 package.scala 96:25:@28610.4]
  wire  _T_1501; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 392:283:@28643.4]
  wire  _T_1502; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 392:291:@28644.4]
  wire  x264; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 402:59:@28655.4]
  wire  _T_1531; // @[package.scala 96:25:@28699.4 package.scala 96:25:@28700.4]
  wire  _T_1533; // @[implicits.scala 55:10:@28701.4]
  wire  _T_1534; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 417:194:@28702.4]
  wire  x493_x265_D20; // @[package.scala 96:25:@28687.4 package.scala 96:25:@28688.4]
  wire  _T_1535; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 417:283:@28703.4]
  wire  _T_1536; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 417:291:@28704.4]
  wire  x269; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 421:59:@28715.4]
  wire  _T_1560; // @[package.scala 96:25:@28748.4 package.scala 96:25:@28749.4]
  wire  _T_1562; // @[implicits.scala 55:10:@28750.4]
  wire  _T_1563; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 432:194:@28751.4]
  wire  x494_x270_D20; // @[package.scala 96:25:@28736.4 package.scala 96:25:@28737.4]
  wire  _T_1564; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 432:283:@28752.4]
  wire  _T_1565; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 432:291:@28753.4]
  wire [31:0] x274_rdrow_number; // @[Math.scala 195:22:@28772.4 Math.scala 196:14:@28773.4]
  wire [31:0] _T_1582; // @[Math.scala 406:49:@28779.4]
  wire [31:0] _T_1584; // @[Math.scala 406:56:@28781.4]
  wire [31:0] _T_1585; // @[Math.scala 406:56:@28782.4]
  wire [31:0] x450_number; // @[implicits.scala 133:21:@28783.4]
  wire  x276; // @[package.scala 96:25:@28797.4 package.scala 96:25:@28798.4]
  wire  x277; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 442:24:@28801.4]
  wire [31:0] _T_1608; // @[Math.scala 406:49:@28810.4]
  wire [31:0] _T_1610; // @[Math.scala 406:56:@28812.4]
  wire [31:0] _T_1611; // @[Math.scala 406:56:@28813.4]
  wire [31:0] _T_1615; // @[package.scala 96:25:@28821.4]
  wire  _T_1619; // @[FixedPoint.scala 50:25:@28828.4]
  wire [1:0] _T_1623; // @[Bitwise.scala 72:12:@28830.4]
  wire [29:0] _T_1624; // @[FixedPoint.scala 18:52:@28831.4]
  wire  _T_1630; // @[Math.scala 451:55:@28833.4]
  wire [1:0] _T_1631; // @[FixedPoint.scala 18:52:@28834.4]
  wire  _T_1637; // @[Math.scala 451:110:@28836.4]
  wire  _T_1638; // @[Math.scala 451:94:@28837.4]
  wire [31:0] _T_1642; // @[package.scala 96:25:@28845.4 package.scala 96:25:@28846.4]
  wire [31:0] x280_1_number; // @[Math.scala 454:20:@28847.4]
  wire [40:0] _GEN_4; // @[Math.scala 461:32:@28852.4]
  wire [40:0] _T_1647; // @[Math.scala 461:32:@28852.4]
  wire [38:0] _GEN_5; // @[Math.scala 461:32:@28857.4]
  wire [38:0] _T_1650; // @[Math.scala 461:32:@28857.4]
  wire  _T_1680; // @[package.scala 96:25:@28925.4 package.scala 96:25:@28926.4]
  wire  _T_1682; // @[implicits.scala 55:10:@28927.4]
  wire  _T_1683; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 469:194:@28928.4]
  wire  x497_x278_D20; // @[package.scala 96:25:@28904.4 package.scala 96:25:@28905.4]
  wire  _T_1684; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 469:283:@28929.4]
  wire  _T_1685; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 469:291:@28930.4]
  wire  x285; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 473:24:@28941.4]
  wire  _T_1712; // @[package.scala 96:25:@28983.4 package.scala 96:25:@28984.4]
  wire  _T_1714; // @[implicits.scala 55:10:@28985.4]
  wire  _T_1715; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 486:194:@28986.4]
  wire  x500_x286_D20; // @[package.scala 96:25:@28971.4 package.scala 96:25:@28972.4]
  wire  _T_1716; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 486:283:@28987.4]
  wire  _T_1717; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 486:291:@28988.4]
  wire  x290; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 490:24:@28999.4]
  wire  _T_1741; // @[package.scala 96:25:@29032.4 package.scala 96:25:@29033.4]
  wire  _T_1743; // @[implicits.scala 55:10:@29034.4]
  wire  _T_1744; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 501:194:@29035.4]
  wire  x501_x291_D20; // @[package.scala 96:25:@29020.4 package.scala 96:25:@29021.4]
  wire  _T_1745; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 501:283:@29036.4]
  wire  _T_1746; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 501:291:@29037.4]
  wire  _T_1873; // @[package.scala 96:25:@29313.4 package.scala 96:25:@29314.4]
  wire  _T_1875; // @[implicits.scala 55:10:@29315.4]
  wire  x504_b213_D66; // @[package.scala 96:25:@29304.4 package.scala 96:25:@29305.4]
  wire  _T_1876; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 563:117:@29316.4]
  wire  x503_b214_D66; // @[package.scala 96:25:@29295.4 package.scala 96:25:@29296.4]
  wire  _T_1877; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 563:123:@29317.4]
  wire [31:0] x226_sum_number; // @[Math.scala 154:22:@27452.4 Math.scala 155:14:@27453.4]
  wire [31:0] x465_x397_D13_number; // @[package.scala 96:25:@27461.4 package.scala 96:25:@27462.4]
  wire [31:0] x467_x375_D21_number; // @[package.scala 96:25:@27479.4 package.scala 96:25:@27480.4]
  wire [31:0] x472_x397_D37_number; // @[package.scala 96:25:@27583.4 package.scala 96:25:@27584.4]
  wire [31:0] x473_x375_D45_number; // @[package.scala 96:25:@27592.4 package.scala 96:25:@27593.4]
  wire [31:0] x475_x226_sum_D24_number; // @[package.scala 96:25:@27610.4 package.scala 96:25:@27611.4]
  wire [31:0] x241_sum_number; // @[Math.scala 154:22:@28020.4 Math.scala 155:14:@28021.4]
  wire [31:0] x482_x422_D13_number; // @[package.scala 96:25:@28038.4 package.scala 96:25:@28039.4]
  wire [31:0] x250_sum_number; // @[Math.scala 154:22:@28414.4 Math.scala 155:14:@28415.4]
  wire [31:0] x485_x444_D13_number; // @[package.scala 96:25:@28432.4 package.scala 96:25:@28433.4]
  wire [31:0] x490_x261_sum_D1_number; // @[package.scala 96:25:@28618.4 package.scala 96:25:@28619.4]
  wire [31:0] x491_x446_D20_number; // @[package.scala 96:25:@28627.4 package.scala 96:25:@28628.4]
  wire [31:0] x266_sum_number; // @[Math.scala 154:22:@28678.4 Math.scala 155:14:@28679.4]
  wire [31:0] x271_sum_number; // @[Math.scala 154:22:@28727.4 Math.scala 155:14:@28728.4]
  wire [31:0] x496_x451_D20_number; // @[package.scala 96:25:@28895.4 package.scala 96:25:@28896.4]
  wire [31:0] x498_x282_sum_D1_number; // @[package.scala 96:25:@28913.4 package.scala 96:25:@28914.4]
  wire [31:0] x287_sum_number; // @[Math.scala 154:22:@28962.4 Math.scala 155:14:@28963.4]
  wire [31:0] x292_sum_number; // @[Math.scala 154:22:@29011.4 Math.scala 155:14:@29012.4]
  _ _ ( // @[Math.scala 720:24:@26946.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@26958.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@26981.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x217_lb_0 x217_lb_0 ( // @[m_x217_lb_0.scala 35:17:@26991.4]
    .clock(x217_lb_0_clock),
    .reset(x217_lb_0_reset),
    .io_rPort_8_banks_1(x217_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x217_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x217_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x217_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x217_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x217_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x217_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x217_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x217_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x217_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x217_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x217_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x217_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x217_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x217_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x217_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x217_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x217_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x217_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x217_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x217_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x217_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x217_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x217_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x217_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x217_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x217_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x217_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x217_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x217_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x217_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x217_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x217_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x217_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x217_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x217_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x217_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x217_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x217_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x217_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x217_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x217_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x217_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x217_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x217_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x217_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x217_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x217_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x217_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x217_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x217_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x217_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x217_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x217_lb_0_io_rPort_0_output_0),
    .io_wPort_0_banks_1(x217_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x217_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x217_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x217_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x217_lb_0_io_wPort_0_en_0)
  );
  x198_sum x378_sum_1 ( // @[Math.scala 150:24:@27116.4]
    .clock(x378_sum_1_clock),
    .reset(x378_sum_1_reset),
    .io_a(x378_sum_1_io_a),
    .io_b(x378_sum_1_io_b),
    .io_flow(x378_sum_1_io_flow),
    .io_result(x378_sum_1_io_result)
  );
  x198_sum x381_sum_1 ( // @[Math.scala 150:24:@27154.4]
    .clock(x381_sum_1_clock),
    .reset(x381_sum_1_reset),
    .io_a(x381_sum_1_io_a),
    .io_b(x381_sum_1_io_b),
    .io_flow(x381_sum_1_io_flow),
    .io_result(x381_sum_1_io_result)
  );
  x198_sum x384_sum_1 ( // @[Math.scala 150:24:@27192.4]
    .clock(x384_sum_1_clock),
    .reset(x384_sum_1_reset),
    .io_a(x384_sum_1_io_a),
    .io_b(x384_sum_1_io_b),
    .io_flow(x384_sum_1_io_flow),
    .io_result(x384_sum_1_io_result)
  );
  x198_sum x387_sum_1 ( // @[Math.scala 150:24:@27230.4]
    .clock(x387_sum_1_clock),
    .reset(x387_sum_1_reset),
    .io_a(x387_sum_1_io_a),
    .io_b(x387_sum_1_io_b),
    .io_flow(x387_sum_1_io_flow),
    .io_result(x387_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_1 ( // @[package.scala 93:22:@27253.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_2 ( // @[package.scala 93:22:@27271.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x198_sum x390_sum_1 ( // @[Math.scala 150:24:@27284.4]
    .clock(x390_sum_1_clock),
    .reset(x390_sum_1_reset),
    .io_a(x390_sum_1_io_a),
    .io_b(x390_sum_1_io_b),
    .io_flow(x390_sum_1_io_flow),
    .io_result(x390_sum_1_io_result)
  );
  x198_sum x393_sum_1 ( // @[Math.scala 150:24:@27322.4]
    .clock(x393_sum_1_clock),
    .reset(x393_sum_1_reset),
    .io_a(x393_sum_1_io_a),
    .io_b(x393_sum_1_io_b),
    .io_flow(x393_sum_1_io_flow),
    .io_result(x393_sum_1_io_result)
  );
  x370_sub x396_sub_1 ( // @[Math.scala 191:24:@27348.4]
    .clock(x396_sub_1_clock),
    .reset(x396_sub_1_reset),
    .io_a(x396_sub_1_io_a),
    .io_b(x396_sub_1_io_b),
    .io_flow(x396_sub_1_io_flow),
    .io_result(x396_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@27358.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@27367.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_5 ( // @[package.scala 93:22:@27376.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  x198_sum x400_sum_1 ( // @[Math.scala 150:24:@27415.4]
    .clock(x400_sum_1_clock),
    .reset(x400_sum_1_reset),
    .io_a(x400_sum_1_io_a),
    .io_b(x400_sum_1_io_b),
    .io_flow(x400_sum_1_io_flow),
    .io_result(x400_sum_1_io_result)
  );
  x225_div x225_div_1 ( // @[Math.scala 327:24:@27427.4]
    .clock(x225_div_1_clock),
    .io_a(x225_div_1_io_a),
    .io_flow(x225_div_1_io_flow),
    .io_result(x225_div_1_io_result)
  );
  RetimeWrapper_184 RetimeWrapper_6 ( // @[package.scala 93:22:@27437.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x198_sum x226_sum_1 ( // @[Math.scala 150:24:@27446.4]
    .clock(x226_sum_1_clock),
    .reset(x226_sum_1_reset),
    .io_a(x226_sum_1_io_a),
    .io_b(x226_sum_1_io_b),
    .io_flow(x226_sum_1_io_flow),
    .io_result(x226_sum_1_io_result)
  );
  RetimeWrapper_186 RetimeWrapper_7 ( // @[package.scala 93:22:@27456.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_187 RetimeWrapper_8 ( // @[package.scala 93:22:@27465.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_188 RetimeWrapper_9 ( // @[package.scala 93:22:@27474.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_189 RetimeWrapper_10 ( // @[package.scala 93:22:@27483.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_189 RetimeWrapper_11 ( // @[package.scala 93:22:@27492.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_189 RetimeWrapper_12 ( // @[package.scala 93:22:@27503.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_192 RetimeWrapper_13 ( // @[package.scala 93:22:@27524.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper RetimeWrapper_14 ( // @[package.scala 93:22:@27538.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_192 RetimeWrapper_15 ( // @[package.scala 93:22:@27547.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper RetimeWrapper_16 ( // @[package.scala 93:22:@27563.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_196 RetimeWrapper_17 ( // @[package.scala 93:22:@27578.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_197 RetimeWrapper_18 ( // @[package.scala 93:22:@27587.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_198 RetimeWrapper_19 ( // @[package.scala 93:22:@27596.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_199 RetimeWrapper_20 ( // @[package.scala 93:22:@27605.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_198 RetimeWrapper_21 ( // @[package.scala 93:22:@27614.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_189 RetimeWrapper_22 ( // @[package.scala 93:22:@27623.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_198 RetimeWrapper_23 ( // @[package.scala 93:22:@27635.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  x370_sub x235_rdcol_1 ( // @[Math.scala 191:24:@27658.4]
    .clock(x235_rdcol_1_clock),
    .reset(x235_rdcol_1_reset),
    .io_a(x235_rdcol_1_io_a),
    .io_b(x235_rdcol_1_io_b),
    .io_flow(x235_rdcol_1_io_flow),
    .io_result(x235_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_24 ( // @[package.scala 93:22:@27673.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper RetimeWrapper_25 ( // @[package.scala 93:22:@27682.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  x198_sum x403_sum_1 ( // @[Math.scala 150:24:@27725.4]
    .clock(x403_sum_1_clock),
    .reset(x403_sum_1_reset),
    .io_a(x403_sum_1_io_a),
    .io_b(x403_sum_1_io_b),
    .io_flow(x403_sum_1_io_flow),
    .io_result(x403_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_26 ( // @[package.scala 93:22:@27748.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_27 ( // @[package.scala 93:22:@27766.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  x198_sum x406_sum_1 ( // @[Math.scala 150:24:@27779.4]
    .clock(x406_sum_1_clock),
    .reset(x406_sum_1_reset),
    .io_a(x406_sum_1_io_a),
    .io_b(x406_sum_1_io_b),
    .io_flow(x406_sum_1_io_flow),
    .io_result(x406_sum_1_io_result)
  );
  x198_sum x409_sum_1 ( // @[Math.scala 150:24:@27817.4]
    .clock(x409_sum_1_clock),
    .reset(x409_sum_1_reset),
    .io_a(x409_sum_1_io_a),
    .io_b(x409_sum_1_io_b),
    .io_flow(x409_sum_1_io_flow),
    .io_result(x409_sum_1_io_result)
  );
  x198_sum x412_sum_1 ( // @[Math.scala 150:24:@27855.4]
    .clock(x412_sum_1_clock),
    .reset(x412_sum_1_reset),
    .io_a(x412_sum_1_io_a),
    .io_b(x412_sum_1_io_b),
    .io_flow(x412_sum_1_io_flow),
    .io_result(x412_sum_1_io_result)
  );
  x198_sum x415_sum_1 ( // @[Math.scala 150:24:@27893.4]
    .clock(x415_sum_1_clock),
    .reset(x415_sum_1_reset),
    .io_a(x415_sum_1_io_a),
    .io_b(x415_sum_1_io_b),
    .io_flow(x415_sum_1_io_flow),
    .io_result(x415_sum_1_io_result)
  );
  x198_sum x418_sum_1 ( // @[Math.scala 150:24:@27931.4]
    .clock(x418_sum_1_clock),
    .reset(x418_sum_1_reset),
    .io_a(x418_sum_1_io_a),
    .io_b(x418_sum_1_io_b),
    .io_flow(x418_sum_1_io_flow),
    .io_result(x418_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_28 ( // @[package.scala 93:22:@27946.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper RetimeWrapper_29 ( // @[package.scala 93:22:@27960.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  x370_sub x421_sub_1 ( // @[Math.scala 191:24:@27971.4]
    .clock(x421_sub_1_clock),
    .reset(x421_sub_1_reset),
    .io_a(x421_sub_1_io_a),
    .io_b(x421_sub_1_io_b),
    .io_flow(x421_sub_1_io_flow),
    .io_result(x421_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_30 ( // @[package.scala 93:22:@27981.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  x225_div x240_div_1 ( // @[Math.scala 327:24:@27995.4]
    .clock(x240_div_1_clock),
    .io_a(x240_div_1_io_a),
    .io_flow(x240_div_1_io_flow),
    .io_result(x240_div_1_io_result)
  );
  RetimeWrapper_218 RetimeWrapper_31 ( // @[package.scala 93:22:@28005.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  x198_sum x241_sum_1 ( // @[Math.scala 150:24:@28014.4]
    .clock(x241_sum_1_clock),
    .reset(x241_sum_1_reset),
    .io_a(x241_sum_1_io_a),
    .io_b(x241_sum_1_io_b),
    .io_flow(x241_sum_1_io_flow),
    .io_result(x241_sum_1_io_result)
  );
  RetimeWrapper_220 RetimeWrapper_32 ( // @[package.scala 93:22:@28024.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_33 ( // @[package.scala 93:22:@28033.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_198 RetimeWrapper_34 ( // @[package.scala 93:22:@28045.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  x370_sub x244_rdcol_1 ( // @[Math.scala 191:24:@28068.4]
    .clock(x244_rdcol_1_clock),
    .reset(x244_rdcol_1_reset),
    .io_a(x244_rdcol_1_io_a),
    .io_b(x244_rdcol_1_io_b),
    .io_flow(x244_rdcol_1_io_flow),
    .io_result(x244_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_35 ( // @[package.scala 93:22:@28083.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  x198_sum x425_sum_1 ( // @[Math.scala 150:24:@28128.4]
    .clock(x425_sum_1_clock),
    .reset(x425_sum_1_reset),
    .io_a(x425_sum_1_io_a),
    .io_b(x425_sum_1_io_b),
    .io_flow(x425_sum_1_io_flow),
    .io_result(x425_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_36 ( // @[package.scala 93:22:@28151.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_37 ( // @[package.scala 93:22:@28169.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  x198_sum x428_sum_1 ( // @[Math.scala 150:24:@28182.4]
    .clock(x428_sum_1_clock),
    .reset(x428_sum_1_reset),
    .io_a(x428_sum_1_io_a),
    .io_b(x428_sum_1_io_b),
    .io_flow(x428_sum_1_io_flow),
    .io_result(x428_sum_1_io_result)
  );
  x198_sum x431_sum_1 ( // @[Math.scala 150:24:@28220.4]
    .clock(x431_sum_1_clock),
    .reset(x431_sum_1_reset),
    .io_a(x431_sum_1_io_a),
    .io_b(x431_sum_1_io_b),
    .io_flow(x431_sum_1_io_flow),
    .io_result(x431_sum_1_io_result)
  );
  x198_sum x434_sum_1 ( // @[Math.scala 150:24:@28258.4]
    .clock(x434_sum_1_clock),
    .reset(x434_sum_1_reset),
    .io_a(x434_sum_1_io_a),
    .io_b(x434_sum_1_io_b),
    .io_flow(x434_sum_1_io_flow),
    .io_result(x434_sum_1_io_result)
  );
  x198_sum x437_sum_1 ( // @[Math.scala 150:24:@28296.4]
    .clock(x437_sum_1_clock),
    .reset(x437_sum_1_reset),
    .io_a(x437_sum_1_io_a),
    .io_b(x437_sum_1_io_b),
    .io_flow(x437_sum_1_io_flow),
    .io_result(x437_sum_1_io_result)
  );
  x198_sum x440_sum_1 ( // @[Math.scala 150:24:@28334.4]
    .clock(x440_sum_1_clock),
    .reset(x440_sum_1_reset),
    .io_a(x440_sum_1_io_a),
    .io_b(x440_sum_1_io_b),
    .io_flow(x440_sum_1_io_flow),
    .io_result(x440_sum_1_io_result)
  );
  RetimeWrapper RetimeWrapper_38 ( // @[package.scala 93:22:@28349.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper RetimeWrapper_39 ( // @[package.scala 93:22:@28363.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  x370_sub x443_sub_1 ( // @[Math.scala 191:24:@28374.4]
    .clock(x443_sub_1_clock),
    .reset(x443_sub_1_reset),
    .io_a(x443_sub_1_io_a),
    .io_b(x443_sub_1_io_b),
    .io_flow(x443_sub_1_io_flow),
    .io_result(x443_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_40 ( // @[package.scala 93:22:@28384.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  x225_div x249_div_1 ( // @[Math.scala 327:24:@28398.4]
    .clock(x249_div_1_clock),
    .io_a(x249_div_1_io_a),
    .io_flow(x249_div_1_io_flow),
    .io_result(x249_div_1_io_result)
  );
  x198_sum x250_sum_1 ( // @[Math.scala 150:24:@28408.4]
    .clock(x250_sum_1_clock),
    .reset(x250_sum_1_reset),
    .io_a(x250_sum_1_io_a),
    .io_b(x250_sum_1_io_b),
    .io_flow(x250_sum_1_io_flow),
    .io_result(x250_sum_1_io_result)
  );
  RetimeWrapper_220 RetimeWrapper_41 ( // @[package.scala 93:22:@28418.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_42 ( // @[package.scala 93:22:@28427.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_198 RetimeWrapper_43 ( // @[package.scala 93:22:@28439.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  x370_sub x253_rdrow_1 ( // @[Math.scala 191:24:@28462.4]
    .clock(x253_rdrow_1_clock),
    .reset(x253_rdrow_1_reset),
    .io_a(x253_rdrow_1_io_a),
    .io_b(x253_rdrow_1_io_b),
    .io_flow(x253_rdrow_1_io_flow),
    .io_result(x253_rdrow_1_io_result)
  );
  RetimeWrapper RetimeWrapper_44 ( // @[package.scala 93:22:@28488.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper RetimeWrapper_45 ( // @[package.scala 93:22:@28497.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_46 ( // @[package.scala 93:22:@28519.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_47 ( // @[package.scala 93:22:@28545.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  x198_sum x449_sum_1 ( // @[Math.scala 150:24:@28566.4]
    .clock(x449_sum_1_clock),
    .reset(x449_sum_1_reset),
    .io_a(x449_sum_1_io_a),
    .io_b(x449_sum_1_io_b),
    .io_flow(x449_sum_1_io_flow),
    .io_result(x449_sum_1_io_result)
  );
  RetimeWrapper_192 RetimeWrapper_48 ( // @[package.scala 93:22:@28576.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_248 RetimeWrapper_49 ( // @[package.scala 93:22:@28585.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  x198_sum x261_sum_1 ( // @[Math.scala 150:24:@28594.4]
    .clock(x261_sum_1_clock),
    .reset(x261_sum_1_reset),
    .io_a(x261_sum_1_io_a),
    .io_b(x261_sum_1_io_b),
    .io_flow(x261_sum_1_io_flow),
    .io_result(x261_sum_1_io_result)
  );
  RetimeWrapper_220 RetimeWrapper_50 ( // @[package.scala 93:22:@28604.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_51 ( // @[package.scala 93:22:@28613.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_187 RetimeWrapper_52 ( // @[package.scala 93:22:@28622.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_198 RetimeWrapper_53 ( // @[package.scala 93:22:@28634.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_254 RetimeWrapper_54 ( // @[package.scala 93:22:@28661.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  x198_sum x266_sum_1 ( // @[Math.scala 150:24:@28672.4]
    .clock(x266_sum_1_clock),
    .reset(x266_sum_1_reset),
    .io_a(x266_sum_1_io_a),
    .io_b(x266_sum_1_io_b),
    .io_flow(x266_sum_1_io_flow),
    .io_result(x266_sum_1_io_result)
  );
  RetimeWrapper_220 RetimeWrapper_55 ( // @[package.scala 93:22:@28682.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_198 RetimeWrapper_56 ( // @[package.scala 93:22:@28694.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  x198_sum x271_sum_1 ( // @[Math.scala 150:24:@28721.4]
    .clock(x271_sum_1_clock),
    .reset(x271_sum_1_reset),
    .io_a(x271_sum_1_io_a),
    .io_b(x271_sum_1_io_b),
    .io_flow(x271_sum_1_io_flow),
    .io_result(x271_sum_1_io_result)
  );
  RetimeWrapper_220 RetimeWrapper_57 ( // @[package.scala 93:22:@28731.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_198 RetimeWrapper_58 ( // @[package.scala 93:22:@28743.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  x370_sub x274_rdrow_1 ( // @[Math.scala 191:24:@28766.4]
    .clock(x274_rdrow_1_clock),
    .reset(x274_rdrow_1_reset),
    .io_a(x274_rdrow_1_io_a),
    .io_b(x274_rdrow_1_io_b),
    .io_flow(x274_rdrow_1_io_flow),
    .io_result(x274_rdrow_1_io_result)
  );
  RetimeWrapper RetimeWrapper_59 ( // @[package.scala 93:22:@28792.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_60 ( // @[package.scala 93:22:@28814.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_61 ( // @[package.scala 93:22:@28840.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  x198_sum x454_sum_1 ( // @[Math.scala 150:24:@28861.4]
    .clock(x454_sum_1_clock),
    .reset(x454_sum_1_reset),
    .io_a(x454_sum_1_io_a),
    .io_b(x454_sum_1_io_b),
    .io_flow(x454_sum_1_io_flow),
    .io_result(x454_sum_1_io_result)
  );
  RetimeWrapper_248 RetimeWrapper_62 ( // @[package.scala 93:22:@28871.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  x198_sum x282_sum_1 ( // @[Math.scala 150:24:@28880.4]
    .clock(x282_sum_1_clock),
    .reset(x282_sum_1_reset),
    .io_a(x282_sum_1_io_a),
    .io_b(x282_sum_1_io_b),
    .io_flow(x282_sum_1_io_flow),
    .io_result(x282_sum_1_io_result)
  );
  RetimeWrapper_187 RetimeWrapper_63 ( // @[package.scala 93:22:@28890.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_220 RetimeWrapper_64 ( // @[package.scala 93:22:@28899.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_65 ( // @[package.scala 93:22:@28908.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_198 RetimeWrapper_66 ( // @[package.scala 93:22:@28920.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_254 RetimeWrapper_67 ( // @[package.scala 93:22:@28947.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  x198_sum x287_sum_1 ( // @[Math.scala 150:24:@28956.4]
    .clock(x287_sum_1_clock),
    .reset(x287_sum_1_reset),
    .io_a(x287_sum_1_io_a),
    .io_b(x287_sum_1_io_b),
    .io_flow(x287_sum_1_io_flow),
    .io_result(x287_sum_1_io_result)
  );
  RetimeWrapper_220 RetimeWrapper_68 ( // @[package.scala 93:22:@28966.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_198 RetimeWrapper_69 ( // @[package.scala 93:22:@28978.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  x198_sum x292_sum_1 ( // @[Math.scala 150:24:@29005.4]
    .clock(x292_sum_1_clock),
    .reset(x292_sum_1_reset),
    .io_a(x292_sum_1_io_a),
    .io_b(x292_sum_1_io_b),
    .io_flow(x292_sum_1_io_flow),
    .io_result(x292_sum_1_io_result)
  );
  RetimeWrapper_220 RetimeWrapper_70 ( // @[package.scala 93:22:@29015.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_198 RetimeWrapper_71 ( // @[package.scala 93:22:@29027.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  x295 x295_1 ( // @[Math.scala 262:24:@29050.4]
    .clock(x295_1_clock),
    .io_a(x295_1_io_a),
    .io_b(x295_1_io_b),
    .io_flow(x295_1_io_flow),
    .io_result(x295_1_io_result)
  );
  x295 x296_1 ( // @[Math.scala 262:24:@29062.4]
    .clock(x296_1_clock),
    .io_a(x296_1_io_a),
    .io_b(x296_1_io_b),
    .io_flow(x296_1_io_flow),
    .io_result(x296_1_io_result)
  );
  x295 x297_1 ( // @[Math.scala 262:24:@29074.4]
    .clock(x297_1_clock),
    .io_a(x297_1_io_a),
    .io_b(x297_1_io_b),
    .io_flow(x297_1_io_flow),
    .io_result(x297_1_io_result)
  );
  x295 x298_1 ( // @[Math.scala 262:24:@29086.4]
    .clock(x298_1_clock),
    .io_a(x298_1_io_a),
    .io_b(x298_1_io_b),
    .io_flow(x298_1_io_flow),
    .io_result(x298_1_io_result)
  );
  x295 x299_1 ( // @[Math.scala 262:24:@29098.4]
    .clock(x299_1_clock),
    .io_a(x299_1_io_a),
    .io_b(x299_1_io_b),
    .io_flow(x299_1_io_flow),
    .io_result(x299_1_io_result)
  );
  x295 x300_1 ( // @[Math.scala 262:24:@29112.4]
    .clock(x300_1_clock),
    .io_a(x300_1_io_a),
    .io_b(x300_1_io_b),
    .io_flow(x300_1_io_flow),
    .io_result(x300_1_io_result)
  );
  x295 x301_1 ( // @[Math.scala 262:24:@29124.4]
    .clock(x301_1_clock),
    .io_a(x301_1_io_a),
    .io_b(x301_1_io_b),
    .io_flow(x301_1_io_flow),
    .io_result(x301_1_io_result)
  );
  x295 x302_1 ( // @[Math.scala 262:24:@29136.4]
    .clock(x302_1_clock),
    .io_a(x302_1_io_a),
    .io_b(x302_1_io_b),
    .io_flow(x302_1_io_flow),
    .io_result(x302_1_io_result)
  );
  x295 x303_1 ( // @[Math.scala 262:24:@29148.4]
    .clock(x303_1_clock),
    .io_a(x303_1_io_a),
    .io_b(x303_1_io_b),
    .io_flow(x303_1_io_flow),
    .io_result(x303_1_io_result)
  );
  x304_x3 x304_x3_1 ( // @[Math.scala 150:24:@29158.4]
    .clock(x304_x3_1_clock),
    .reset(x304_x3_1_reset),
    .io_a(x304_x3_1_io_a),
    .io_b(x304_x3_1_io_b),
    .io_flow(x304_x3_1_io_flow),
    .io_result(x304_x3_1_io_result)
  );
  x304_x3 x305_x4_1 ( // @[Math.scala 150:24:@29168.4]
    .clock(x305_x4_1_clock),
    .reset(x305_x4_1_reset),
    .io_a(x305_x4_1_io_a),
    .io_b(x305_x4_1_io_b),
    .io_flow(x305_x4_1_io_flow),
    .io_result(x305_x4_1_io_result)
  );
  x304_x3 x306_x3_1 ( // @[Math.scala 150:24:@29178.4]
    .clock(x306_x3_1_clock),
    .reset(x306_x3_1_reset),
    .io_a(x306_x3_1_io_a),
    .io_b(x306_x3_1_io_b),
    .io_flow(x306_x3_1_io_flow),
    .io_result(x306_x3_1_io_result)
  );
  x304_x3 x307_x4_1 ( // @[Math.scala 150:24:@29188.4]
    .clock(x307_x4_1_clock),
    .reset(x307_x4_1_reset),
    .io_a(x307_x4_1_io_a),
    .io_b(x307_x4_1_io_b),
    .io_flow(x307_x4_1_io_flow),
    .io_result(x307_x4_1_io_result)
  );
  x304_x3 x308_x3_1 ( // @[Math.scala 150:24:@29198.4]
    .clock(x308_x3_1_clock),
    .reset(x308_x3_1_reset),
    .io_a(x308_x3_1_io_a),
    .io_b(x308_x3_1_io_b),
    .io_flow(x308_x3_1_io_flow),
    .io_result(x308_x3_1_io_result)
  );
  x304_x3 x309_x4_1 ( // @[Math.scala 150:24:@29208.4]
    .clock(x309_x4_1_clock),
    .reset(x309_x4_1_reset),
    .io_a(x309_x4_1_io_a),
    .io_b(x309_x4_1_io_b),
    .io_flow(x309_x4_1_io_flow),
    .io_result(x309_x4_1_io_result)
  );
  x304_x3 x310_x3_1 ( // @[Math.scala 150:24:@29218.4]
    .clock(x310_x3_1_clock),
    .reset(x310_x3_1_reset),
    .io_a(x310_x3_1_io_a),
    .io_b(x310_x3_1_io_b),
    .io_flow(x310_x3_1_io_flow),
    .io_result(x310_x3_1_io_result)
  );
  RetimeWrapper_286 RetimeWrapper_72 ( // @[package.scala 93:22:@29228.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  x304_x3 x311_sum_1 ( // @[Math.scala 150:24:@29237.4]
    .clock(x311_sum_1_clock),
    .reset(x311_sum_1_reset),
    .io_a(x311_sum_1_io_a),
    .io_b(x311_sum_1_io_b),
    .io_flow(x311_sum_1_io_flow),
    .io_result(x311_sum_1_io_result)
  );
  x312 x312_1 ( // @[Math.scala 720:24:@29247.4]
    .io_b(x312_1_io_b),
    .io_result(x312_1_io_result)
  );
  x313_mul x313_mul_1 ( // @[Math.scala 262:24:@29258.4]
    .clock(x313_mul_1_clock),
    .io_a(x313_mul_1_io_a),
    .io_flow(x313_mul_1_io_flow),
    .io_result(x313_mul_1_io_result)
  );
  x314 x314_1 ( // @[Math.scala 720:24:@29268.4]
    .io_b(x314_1_io_b),
    .io_result(x314_1_io_result)
  );
  RetimeWrapper_286 RetimeWrapper_73 ( // @[package.scala 93:22:@29281.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_46 RetimeWrapper_74 ( // @[package.scala 93:22:@29290.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_46 RetimeWrapper_75 ( // @[package.scala 93:22:@29299.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_46 RetimeWrapper_76 ( // @[package.scala 93:22:@29308.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  assign b213 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 62:18:@26966.4]
  assign b214 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 63:18:@26967.4]
  assign _T_205 = b213 & b214; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 67:30:@26969.4]
  assign _T_206 = _T_205 & io_sigsIn_datapathEn; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 67:37:@26970.4]
  assign _T_210 = io_in_x184_TID == 8'h0; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 69:76:@26975.4]
  assign _T_211 = _T_206 & _T_210; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 69:62:@26976.4]
  assign _T_213 = io_in_x184_TDEST == 8'h0; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 69:101:@26977.4]
  assign b211_number = __io_result; // @[Math.scala 723:22:@26951.4 Math.scala 724:14:@26952.4]
  assign _T_241 = $signed(b211_number); // @[Math.scala 406:49:@27067.4]
  assign _T_243 = $signed(_T_241) & $signed(32'sh3); // @[Math.scala 406:56:@27069.4]
  assign _T_244 = $signed(_T_243); // @[Math.scala 406:56:@27070.4]
  assign x374_number = $unsigned(_T_244); // @[implicits.scala 133:21:@27071.4]
  assign _T_254 = $signed(x374_number); // @[Math.scala 406:49:@27080.4]
  assign _T_256 = $signed(_T_254) & $signed(32'sh3); // @[Math.scala 406:56:@27082.4]
  assign _T_257 = $signed(_T_256); // @[Math.scala 406:56:@27083.4]
  assign b212_number = __1_io_result; // @[Math.scala 723:22:@26963.4 Math.scala 724:14:@26964.4]
  assign _T_261 = b212_number[31]; // @[FixedPoint.scala 50:25:@27089.4]
  assign _T_265 = _T_261 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@27091.4]
  assign _T_266 = b212_number[31:16]; // @[FixedPoint.scala 18:52:@27092.4]
  assign _T_272 = _T_266 == 16'hffff; // @[Math.scala 451:55:@27094.4]
  assign _T_273 = b212_number[15:0]; // @[FixedPoint.scala 18:52:@27095.4]
  assign _T_279 = _T_273 != 16'h0; // @[Math.scala 451:110:@27097.4]
  assign _T_280 = _T_272 & _T_279; // @[Math.scala 451:94:@27098.4]
  assign _T_282 = {_T_265,_T_266}; // @[Cat.scala 30:58:@27100.4]
  assign _T_292 = $signed(b212_number); // @[Math.scala 406:49:@27108.4]
  assign _T_294 = $signed(_T_292) & $signed(32'shffff); // @[Math.scala 406:56:@27110.4]
  assign _T_295 = $signed(_T_294); // @[Math.scala 406:56:@27111.4]
  assign x378_sum_number = x378_sum_1_io_result; // @[Math.scala 154:22:@27122.4 Math.scala 155:14:@27123.4]
  assign _T_302 = x378_sum_number[31]; // @[FixedPoint.scala 50:25:@27127.4]
  assign _T_306 = _T_302 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@27129.4]
  assign _T_307 = x378_sum_number[31:8]; // @[FixedPoint.scala 18:52:@27130.4]
  assign _T_313 = _T_307 == 24'hffffff; // @[Math.scala 451:55:@27132.4]
  assign _T_314 = x378_sum_number[7:0]; // @[FixedPoint.scala 18:52:@27133.4]
  assign _T_320 = _T_314 != 8'h0; // @[Math.scala 451:110:@27135.4]
  assign _T_321 = _T_313 & _T_320; // @[Math.scala 451:94:@27136.4]
  assign _T_323 = {_T_306,_T_307}; // @[Cat.scala 30:58:@27138.4]
  assign _T_333 = $signed(x378_sum_number); // @[Math.scala 406:49:@27146.4]
  assign _T_335 = $signed(_T_333) & $signed(32'shff); // @[Math.scala 406:56:@27148.4]
  assign _T_336 = $signed(_T_335); // @[Math.scala 406:56:@27149.4]
  assign x381_sum_number = x381_sum_1_io_result; // @[Math.scala 154:22:@27160.4 Math.scala 155:14:@27161.4]
  assign _T_343 = x381_sum_number[31]; // @[FixedPoint.scala 50:25:@27165.4]
  assign _T_347 = _T_343 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@27167.4]
  assign _T_348 = x381_sum_number[31:4]; // @[FixedPoint.scala 18:52:@27168.4]
  assign _T_354 = _T_348 == 28'hfffffff; // @[Math.scala 451:55:@27170.4]
  assign _T_355 = x381_sum_number[3:0]; // @[FixedPoint.scala 18:52:@27171.4]
  assign _T_361 = _T_355 != 4'h0; // @[Math.scala 451:110:@27173.4]
  assign _T_362 = _T_354 & _T_361; // @[Math.scala 451:94:@27174.4]
  assign _T_364 = {_T_347,_T_348}; // @[Cat.scala 30:58:@27176.4]
  assign _T_374 = $signed(x381_sum_number); // @[Math.scala 406:49:@27184.4]
  assign _T_376 = $signed(_T_374) & $signed(32'shf); // @[Math.scala 406:56:@27186.4]
  assign _T_377 = $signed(_T_376); // @[Math.scala 406:56:@27187.4]
  assign x384_sum_number = x384_sum_1_io_result; // @[Math.scala 154:22:@27198.4 Math.scala 155:14:@27199.4]
  assign _T_384 = x384_sum_number[31]; // @[FixedPoint.scala 50:25:@27203.4]
  assign _T_388 = _T_384 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27205.4]
  assign _T_389 = x384_sum_number[31:2]; // @[FixedPoint.scala 18:52:@27206.4]
  assign _T_395 = _T_389 == 30'h3fffffff; // @[Math.scala 451:55:@27208.4]
  assign _T_396 = x384_sum_number[1:0]; // @[FixedPoint.scala 18:52:@27209.4]
  assign _T_402 = _T_396 != 2'h0; // @[Math.scala 451:110:@27211.4]
  assign _T_403 = _T_395 & _T_402; // @[Math.scala 451:94:@27212.4]
  assign _T_405 = {_T_388,_T_389}; // @[Cat.scala 30:58:@27214.4]
  assign _T_415 = $signed(x384_sum_number); // @[Math.scala 406:49:@27222.4]
  assign _T_417 = $signed(_T_415) & $signed(32'sh3); // @[Math.scala 406:56:@27224.4]
  assign _T_418 = $signed(_T_417); // @[Math.scala 406:56:@27225.4]
  assign x387_sum_number = x387_sum_1_io_result; // @[Math.scala 154:22:@27236.4 Math.scala 155:14:@27237.4]
  assign _T_425 = x387_sum_number[31]; // @[FixedPoint.scala 50:25:@27241.4]
  assign _T_429 = _T_425 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27243.4]
  assign _T_430 = x387_sum_number[31:2]; // @[FixedPoint.scala 18:52:@27244.4]
  assign _T_436 = _T_430 == 30'h3fffffff; // @[Math.scala 451:55:@27246.4]
  assign _T_437 = x387_sum_number[1:0]; // @[FixedPoint.scala 18:52:@27247.4]
  assign _T_443 = _T_437 != 2'h0; // @[Math.scala 451:110:@27249.4]
  assign _T_444 = _T_436 & _T_443; // @[Math.scala 451:94:@27250.4]
  assign _T_448 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@27258.4 package.scala 96:25:@27259.4]
  assign _T_458 = $signed(x387_sum_number); // @[Math.scala 406:49:@27267.4]
  assign _T_460 = $signed(_T_458) & $signed(32'sh3); // @[Math.scala 406:56:@27269.4]
  assign _T_461 = $signed(_T_460); // @[Math.scala 406:56:@27270.4]
  assign _T_465 = $signed(RetimeWrapper_2_io_out); // @[package.scala 96:25:@27278.4]
  assign x390_sum_number = x390_sum_1_io_result; // @[Math.scala 154:22:@27290.4 Math.scala 155:14:@27291.4]
  assign _T_472 = x390_sum_number[31]; // @[FixedPoint.scala 50:25:@27295.4]
  assign _T_476 = _T_472 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27297.4]
  assign _T_477 = x390_sum_number[31:2]; // @[FixedPoint.scala 18:52:@27298.4]
  assign _T_483 = _T_477 == 30'h3fffffff; // @[Math.scala 451:55:@27300.4]
  assign _T_484 = x390_sum_number[1:0]; // @[FixedPoint.scala 18:52:@27301.4]
  assign _T_490 = _T_484 != 2'h0; // @[Math.scala 451:110:@27303.4]
  assign _T_491 = _T_483 & _T_490; // @[Math.scala 451:94:@27304.4]
  assign _T_493 = {_T_476,_T_477}; // @[Cat.scala 30:58:@27306.4]
  assign _T_503 = $signed(x390_sum_number); // @[Math.scala 406:49:@27314.4]
  assign _T_505 = $signed(_T_503) & $signed(32'sh3); // @[Math.scala 406:56:@27316.4]
  assign _T_506 = $signed(_T_505); // @[Math.scala 406:56:@27317.4]
  assign x393_sum_number = x393_sum_1_io_result; // @[Math.scala 154:22:@27328.4 Math.scala 155:14:@27329.4]
  assign _T_516 = $signed(x393_sum_number); // @[Math.scala 476:37:@27334.4]
  assign x462_x394_D1 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@27372.4 package.scala 96:25:@27373.4]
  assign x463_x393_sum_D1_number = RetimeWrapper_5_io_out; // @[package.scala 96:25:@27381.4 package.scala 96:25:@27382.4]
  assign x396_sub_number = x396_sub_1_io_result; // @[Math.scala 195:22:@27354.4 Math.scala 196:14:@27355.4]
  assign _T_547 = x374_number[31]; // @[FixedPoint.scala 50:25:@27389.4]
  assign _T_551 = _T_547 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27391.4]
  assign _T_552 = x374_number[31:2]; // @[FixedPoint.scala 18:52:@27392.4]
  assign _T_558 = _T_552 == 30'h3fffffff; // @[Math.scala 451:55:@27394.4]
  assign _T_559 = x374_number[1:0]; // @[FixedPoint.scala 18:52:@27395.4]
  assign _T_565 = _T_559 != 2'h0; // @[Math.scala 451:110:@27397.4]
  assign _T_566 = _T_558 & _T_565; // @[Math.scala 451:94:@27398.4]
  assign _T_568 = {_T_551,_T_552}; // @[Cat.scala 30:58:@27400.4]
  assign x223_1_number = _T_566 ? 32'h0 : _T_568; // @[Math.scala 454:20:@27401.4]
  assign _GEN_0 = {{9'd0}, x223_1_number}; // @[Math.scala 461:32:@27406.4]
  assign _T_573 = _GEN_0 << 9; // @[Math.scala 461:32:@27406.4]
  assign _GEN_1 = {{7'd0}, x223_1_number}; // @[Math.scala 461:32:@27411.4]
  assign _T_576 = _GEN_1 << 7; // @[Math.scala 461:32:@27411.4]
  assign _T_609 = ~ io_sigsIn_break; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 163:101:@27500.4]
  assign _T_613 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@27508.4 package.scala 96:25:@27509.4]
  assign _T_615 = io_rr ? _T_613 : 1'h0; // @[implicits.scala 55:10:@27510.4]
  assign _T_616 = _T_609 & _T_615; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 163:118:@27511.4]
  assign _T_618 = _T_616 & _T_609; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 163:207:@27513.4]
  assign _T_619 = _T_618 & io_sigsIn_backpressure; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 163:226:@27514.4]
  assign x468_b213_D21 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@27488.4 package.scala 96:25:@27489.4]
  assign _T_620 = _T_619 & x468_b213_D21; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 163:252:@27515.4]
  assign x469_b214_D21 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@27497.4 package.scala 96:25:@27498.4]
  assign x470_b211_D23_number = RetimeWrapper_13_io_out; // @[package.scala 96:25:@27529.4 package.scala 96:25:@27530.4]
  assign _T_630 = $signed(x470_b211_D23_number); // @[Math.scala 476:37:@27535.4]
  assign x471_b212_D23_number = RetimeWrapper_15_io_out; // @[package.scala 96:25:@27552.4 package.scala 96:25:@27553.4]
  assign _T_645 = $signed(x471_b212_D23_number); // @[Math.scala 476:37:@27560.4]
  assign x229 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@27543.4 package.scala 96:25:@27544.4]
  assign x230 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@27568.4 package.scala 96:25:@27569.4]
  assign x231 = x229 | x230; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 182:59:@27572.4]
  assign _T_683 = RetimeWrapper_23_io_out; // @[package.scala 96:25:@27640.4 package.scala 96:25:@27641.4]
  assign _T_685 = io_rr ? _T_683 : 1'h0; // @[implicits.scala 55:10:@27642.4]
  assign _T_686 = _T_609 & _T_685; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 201:194:@27643.4]
  assign x477_x232_D21 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@27628.4 package.scala 96:25:@27629.4]
  assign _T_687 = _T_686 & x477_x232_D21; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 201:283:@27644.4]
  assign x474_b213_D45 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@27601.4 package.scala 96:25:@27602.4]
  assign _T_688 = _T_687 & x474_b213_D45; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 201:291:@27645.4]
  assign x476_b214_D45 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@27619.4 package.scala 96:25:@27620.4]
  assign x235_rdcol_number = x235_rdcol_1_io_result; // @[Math.scala 195:22:@27664.4 Math.scala 196:14:@27665.4]
  assign _T_703 = $signed(x235_rdcol_number); // @[Math.scala 476:37:@27670.4]
  assign x478_x229_D1 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@27687.4 package.scala 96:25:@27688.4]
  assign x236 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@27678.4 package.scala 96:25:@27679.4]
  assign x237 = x478_x229_D1 | x236; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 211:24:@27691.4]
  assign _T_717 = x235_rdcol_number[31]; // @[FixedPoint.scala 50:25:@27698.4]
  assign _T_721 = _T_717 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@27700.4]
  assign _T_722 = x235_rdcol_number[31:16]; // @[FixedPoint.scala 18:52:@27701.4]
  assign _T_728 = _T_722 == 16'hffff; // @[Math.scala 451:55:@27703.4]
  assign _T_729 = x235_rdcol_number[15:0]; // @[FixedPoint.scala 18:52:@27704.4]
  assign _T_735 = _T_729 != 16'h0; // @[Math.scala 451:110:@27706.4]
  assign _T_736 = _T_728 & _T_735; // @[Math.scala 451:94:@27707.4]
  assign _T_738 = {_T_721,_T_722}; // @[Cat.scala 30:58:@27709.4]
  assign _T_750 = $signed(_T_703) & $signed(32'shffff); // @[Math.scala 406:56:@27719.4]
  assign _T_751 = $signed(_T_750); // @[Math.scala 406:56:@27720.4]
  assign x403_sum_number = x403_sum_1_io_result; // @[Math.scala 154:22:@27731.4 Math.scala 155:14:@27732.4]
  assign _T_758 = x403_sum_number[31]; // @[FixedPoint.scala 50:25:@27736.4]
  assign _T_762 = _T_758 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@27738.4]
  assign _T_763 = x403_sum_number[31:8]; // @[FixedPoint.scala 18:52:@27739.4]
  assign _T_769 = _T_763 == 24'hffffff; // @[Math.scala 451:55:@27741.4]
  assign _T_770 = x403_sum_number[7:0]; // @[FixedPoint.scala 18:52:@27742.4]
  assign _T_776 = _T_770 != 8'h0; // @[Math.scala 451:110:@27744.4]
  assign _T_777 = _T_769 & _T_776; // @[Math.scala 451:94:@27745.4]
  assign _T_781 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@27753.4 package.scala 96:25:@27754.4]
  assign _T_791 = $signed(x403_sum_number); // @[Math.scala 406:49:@27762.4]
  assign _T_793 = $signed(_T_791) & $signed(32'shff); // @[Math.scala 406:56:@27764.4]
  assign _T_794 = $signed(_T_793); // @[Math.scala 406:56:@27765.4]
  assign _T_798 = $signed(RetimeWrapper_27_io_out); // @[package.scala 96:25:@27773.4]
  assign x406_sum_number = x406_sum_1_io_result; // @[Math.scala 154:22:@27785.4 Math.scala 155:14:@27786.4]
  assign _T_805 = x406_sum_number[31]; // @[FixedPoint.scala 50:25:@27790.4]
  assign _T_809 = _T_805 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@27792.4]
  assign _T_810 = x406_sum_number[31:4]; // @[FixedPoint.scala 18:52:@27793.4]
  assign _T_816 = _T_810 == 28'hfffffff; // @[Math.scala 451:55:@27795.4]
  assign _T_817 = x406_sum_number[3:0]; // @[FixedPoint.scala 18:52:@27796.4]
  assign _T_823 = _T_817 != 4'h0; // @[Math.scala 451:110:@27798.4]
  assign _T_824 = _T_816 & _T_823; // @[Math.scala 451:94:@27799.4]
  assign _T_826 = {_T_809,_T_810}; // @[Cat.scala 30:58:@27801.4]
  assign _T_836 = $signed(x406_sum_number); // @[Math.scala 406:49:@27809.4]
  assign _T_838 = $signed(_T_836) & $signed(32'shf); // @[Math.scala 406:56:@27811.4]
  assign _T_839 = $signed(_T_838); // @[Math.scala 406:56:@27812.4]
  assign x409_sum_number = x409_sum_1_io_result; // @[Math.scala 154:22:@27823.4 Math.scala 155:14:@27824.4]
  assign _T_846 = x409_sum_number[31]; // @[FixedPoint.scala 50:25:@27828.4]
  assign _T_850 = _T_846 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27830.4]
  assign _T_851 = x409_sum_number[31:2]; // @[FixedPoint.scala 18:52:@27831.4]
  assign _T_857 = _T_851 == 30'h3fffffff; // @[Math.scala 451:55:@27833.4]
  assign _T_858 = x409_sum_number[1:0]; // @[FixedPoint.scala 18:52:@27834.4]
  assign _T_864 = _T_858 != 2'h0; // @[Math.scala 451:110:@27836.4]
  assign _T_865 = _T_857 & _T_864; // @[Math.scala 451:94:@27837.4]
  assign _T_867 = {_T_850,_T_851}; // @[Cat.scala 30:58:@27839.4]
  assign _T_877 = $signed(x409_sum_number); // @[Math.scala 406:49:@27847.4]
  assign _T_879 = $signed(_T_877) & $signed(32'sh3); // @[Math.scala 406:56:@27849.4]
  assign _T_880 = $signed(_T_879); // @[Math.scala 406:56:@27850.4]
  assign x412_sum_number = x412_sum_1_io_result; // @[Math.scala 154:22:@27861.4 Math.scala 155:14:@27862.4]
  assign _T_887 = x412_sum_number[31]; // @[FixedPoint.scala 50:25:@27866.4]
  assign _T_891 = _T_887 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27868.4]
  assign _T_892 = x412_sum_number[31:2]; // @[FixedPoint.scala 18:52:@27869.4]
  assign _T_898 = _T_892 == 30'h3fffffff; // @[Math.scala 451:55:@27871.4]
  assign _T_899 = x412_sum_number[1:0]; // @[FixedPoint.scala 18:52:@27872.4]
  assign _T_905 = _T_899 != 2'h0; // @[Math.scala 451:110:@27874.4]
  assign _T_906 = _T_898 & _T_905; // @[Math.scala 451:94:@27875.4]
  assign _T_908 = {_T_891,_T_892}; // @[Cat.scala 30:58:@27877.4]
  assign _T_918 = $signed(x412_sum_number); // @[Math.scala 406:49:@27885.4]
  assign _T_920 = $signed(_T_918) & $signed(32'sh3); // @[Math.scala 406:56:@27887.4]
  assign _T_921 = $signed(_T_920); // @[Math.scala 406:56:@27888.4]
  assign x415_sum_number = x415_sum_1_io_result; // @[Math.scala 154:22:@27899.4 Math.scala 155:14:@27900.4]
  assign _T_928 = x415_sum_number[31]; // @[FixedPoint.scala 50:25:@27904.4]
  assign _T_932 = _T_928 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27906.4]
  assign _T_933 = x415_sum_number[31:2]; // @[FixedPoint.scala 18:52:@27907.4]
  assign _T_939 = _T_933 == 30'h3fffffff; // @[Math.scala 451:55:@27909.4]
  assign _T_940 = x415_sum_number[1:0]; // @[FixedPoint.scala 18:52:@27910.4]
  assign _T_946 = _T_940 != 2'h0; // @[Math.scala 451:110:@27912.4]
  assign _T_947 = _T_939 & _T_946; // @[Math.scala 451:94:@27913.4]
  assign _T_949 = {_T_932,_T_933}; // @[Cat.scala 30:58:@27915.4]
  assign _T_959 = $signed(x415_sum_number); // @[Math.scala 406:49:@27923.4]
  assign _T_961 = $signed(_T_959) & $signed(32'sh3); // @[Math.scala 406:56:@27925.4]
  assign _T_962 = $signed(_T_961); // @[Math.scala 406:56:@27926.4]
  assign x418_sum_number = x418_sum_1_io_result; // @[Math.scala 154:22:@27937.4 Math.scala 155:14:@27938.4]
  assign _T_972 = $signed(x418_sum_number); // @[Math.scala 476:37:@27943.4]
  assign x419 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@27951.4 package.scala 96:25:@27952.4]
  assign x479_x418_sum_D1_number = RetimeWrapper_30_io_out; // @[package.scala 96:25:@27986.4 package.scala 96:25:@27987.4]
  assign x421_sub_number = x421_sub_1_io_result; // @[Math.scala 195:22:@27977.4 Math.scala 196:14:@27978.4]
  assign _T_1029 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@28050.4 package.scala 96:25:@28051.4]
  assign _T_1031 = io_rr ? _T_1029 : 1'h0; // @[implicits.scala 55:10:@28052.4]
  assign _T_1032 = _T_609 & _T_1031; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 274:194:@28053.4]
  assign x481_x238_D20 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@28029.4 package.scala 96:25:@28030.4]
  assign _T_1033 = _T_1032 & x481_x238_D20; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 274:283:@28054.4]
  assign _T_1034 = _T_1033 & x474_b213_D45; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 274:291:@28055.4]
  assign x244_rdcol_number = x244_rdcol_1_io_result; // @[Math.scala 195:22:@28074.4 Math.scala 196:14:@28075.4]
  assign _T_1049 = $signed(x244_rdcol_number); // @[Math.scala 476:37:@28080.4]
  assign x245 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@28088.4 package.scala 96:25:@28089.4]
  assign x246 = x478_x229_D1 | x245; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 288:59:@28092.4]
  assign _T_1062 = x244_rdcol_number[31]; // @[FixedPoint.scala 50:25:@28101.4]
  assign _T_1066 = _T_1062 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@28103.4]
  assign _T_1067 = x244_rdcol_number[31:16]; // @[FixedPoint.scala 18:52:@28104.4]
  assign _T_1073 = _T_1067 == 16'hffff; // @[Math.scala 451:55:@28106.4]
  assign _T_1074 = x244_rdcol_number[15:0]; // @[FixedPoint.scala 18:52:@28107.4]
  assign _T_1080 = _T_1074 != 16'h0; // @[Math.scala 451:110:@28109.4]
  assign _T_1081 = _T_1073 & _T_1080; // @[Math.scala 451:94:@28110.4]
  assign _T_1083 = {_T_1066,_T_1067}; // @[Cat.scala 30:58:@28112.4]
  assign _T_1095 = $signed(_T_1049) & $signed(32'shffff); // @[Math.scala 406:56:@28122.4]
  assign _T_1096 = $signed(_T_1095); // @[Math.scala 406:56:@28123.4]
  assign x425_sum_number = x425_sum_1_io_result; // @[Math.scala 154:22:@28134.4 Math.scala 155:14:@28135.4]
  assign _T_1103 = x425_sum_number[31]; // @[FixedPoint.scala 50:25:@28139.4]
  assign _T_1107 = _T_1103 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@28141.4]
  assign _T_1108 = x425_sum_number[31:8]; // @[FixedPoint.scala 18:52:@28142.4]
  assign _T_1114 = _T_1108 == 24'hffffff; // @[Math.scala 451:55:@28144.4]
  assign _T_1115 = x425_sum_number[7:0]; // @[FixedPoint.scala 18:52:@28145.4]
  assign _T_1121 = _T_1115 != 8'h0; // @[Math.scala 451:110:@28147.4]
  assign _T_1122 = _T_1114 & _T_1121; // @[Math.scala 451:94:@28148.4]
  assign _T_1126 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@28156.4 package.scala 96:25:@28157.4]
  assign _T_1136 = $signed(x425_sum_number); // @[Math.scala 406:49:@28165.4]
  assign _T_1138 = $signed(_T_1136) & $signed(32'shff); // @[Math.scala 406:56:@28167.4]
  assign _T_1139 = $signed(_T_1138); // @[Math.scala 406:56:@28168.4]
  assign _T_1143 = $signed(RetimeWrapper_37_io_out); // @[package.scala 96:25:@28176.4]
  assign x428_sum_number = x428_sum_1_io_result; // @[Math.scala 154:22:@28188.4 Math.scala 155:14:@28189.4]
  assign _T_1150 = x428_sum_number[31]; // @[FixedPoint.scala 50:25:@28193.4]
  assign _T_1154 = _T_1150 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@28195.4]
  assign _T_1155 = x428_sum_number[31:4]; // @[FixedPoint.scala 18:52:@28196.4]
  assign _T_1161 = _T_1155 == 28'hfffffff; // @[Math.scala 451:55:@28198.4]
  assign _T_1162 = x428_sum_number[3:0]; // @[FixedPoint.scala 18:52:@28199.4]
  assign _T_1168 = _T_1162 != 4'h0; // @[Math.scala 451:110:@28201.4]
  assign _T_1169 = _T_1161 & _T_1168; // @[Math.scala 451:94:@28202.4]
  assign _T_1171 = {_T_1154,_T_1155}; // @[Cat.scala 30:58:@28204.4]
  assign _T_1181 = $signed(x428_sum_number); // @[Math.scala 406:49:@28212.4]
  assign _T_1183 = $signed(_T_1181) & $signed(32'shf); // @[Math.scala 406:56:@28214.4]
  assign _T_1184 = $signed(_T_1183); // @[Math.scala 406:56:@28215.4]
  assign x431_sum_number = x431_sum_1_io_result; // @[Math.scala 154:22:@28226.4 Math.scala 155:14:@28227.4]
  assign _T_1191 = x431_sum_number[31]; // @[FixedPoint.scala 50:25:@28231.4]
  assign _T_1195 = _T_1191 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28233.4]
  assign _T_1196 = x431_sum_number[31:2]; // @[FixedPoint.scala 18:52:@28234.4]
  assign _T_1202 = _T_1196 == 30'h3fffffff; // @[Math.scala 451:55:@28236.4]
  assign _T_1203 = x431_sum_number[1:0]; // @[FixedPoint.scala 18:52:@28237.4]
  assign _T_1209 = _T_1203 != 2'h0; // @[Math.scala 451:110:@28239.4]
  assign _T_1210 = _T_1202 & _T_1209; // @[Math.scala 451:94:@28240.4]
  assign _T_1212 = {_T_1195,_T_1196}; // @[Cat.scala 30:58:@28242.4]
  assign _T_1222 = $signed(x431_sum_number); // @[Math.scala 406:49:@28250.4]
  assign _T_1224 = $signed(_T_1222) & $signed(32'sh3); // @[Math.scala 406:56:@28252.4]
  assign _T_1225 = $signed(_T_1224); // @[Math.scala 406:56:@28253.4]
  assign x434_sum_number = x434_sum_1_io_result; // @[Math.scala 154:22:@28264.4 Math.scala 155:14:@28265.4]
  assign _T_1232 = x434_sum_number[31]; // @[FixedPoint.scala 50:25:@28269.4]
  assign _T_1236 = _T_1232 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28271.4]
  assign _T_1237 = x434_sum_number[31:2]; // @[FixedPoint.scala 18:52:@28272.4]
  assign _T_1243 = _T_1237 == 30'h3fffffff; // @[Math.scala 451:55:@28274.4]
  assign _T_1244 = x434_sum_number[1:0]; // @[FixedPoint.scala 18:52:@28275.4]
  assign _T_1250 = _T_1244 != 2'h0; // @[Math.scala 451:110:@28277.4]
  assign _T_1251 = _T_1243 & _T_1250; // @[Math.scala 451:94:@28278.4]
  assign _T_1253 = {_T_1236,_T_1237}; // @[Cat.scala 30:58:@28280.4]
  assign _T_1263 = $signed(x434_sum_number); // @[Math.scala 406:49:@28288.4]
  assign _T_1265 = $signed(_T_1263) & $signed(32'sh3); // @[Math.scala 406:56:@28290.4]
  assign _T_1266 = $signed(_T_1265); // @[Math.scala 406:56:@28291.4]
  assign x437_sum_number = x437_sum_1_io_result; // @[Math.scala 154:22:@28302.4 Math.scala 155:14:@28303.4]
  assign _T_1273 = x437_sum_number[31]; // @[FixedPoint.scala 50:25:@28307.4]
  assign _T_1277 = _T_1273 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28309.4]
  assign _T_1278 = x437_sum_number[31:2]; // @[FixedPoint.scala 18:52:@28310.4]
  assign _T_1284 = _T_1278 == 30'h3fffffff; // @[Math.scala 451:55:@28312.4]
  assign _T_1285 = x437_sum_number[1:0]; // @[FixedPoint.scala 18:52:@28313.4]
  assign _T_1291 = _T_1285 != 2'h0; // @[Math.scala 451:110:@28315.4]
  assign _T_1292 = _T_1284 & _T_1291; // @[Math.scala 451:94:@28316.4]
  assign _T_1294 = {_T_1277,_T_1278}; // @[Cat.scala 30:58:@28318.4]
  assign _T_1304 = $signed(x437_sum_number); // @[Math.scala 406:49:@28326.4]
  assign _T_1306 = $signed(_T_1304) & $signed(32'sh3); // @[Math.scala 406:56:@28328.4]
  assign _T_1307 = $signed(_T_1306); // @[Math.scala 406:56:@28329.4]
  assign x440_sum_number = x440_sum_1_io_result; // @[Math.scala 154:22:@28340.4 Math.scala 155:14:@28341.4]
  assign _T_1317 = $signed(x440_sum_number); // @[Math.scala 476:37:@28346.4]
  assign x441 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@28354.4 package.scala 96:25:@28355.4]
  assign x483_x440_sum_D1_number = RetimeWrapper_40_io_out; // @[package.scala 96:25:@28389.4 package.scala 96:25:@28390.4]
  assign x443_sub_number = x443_sub_1_io_result; // @[Math.scala 195:22:@28380.4 Math.scala 196:14:@28381.4]
  assign _T_1371 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@28444.4 package.scala 96:25:@28445.4]
  assign _T_1373 = io_rr ? _T_1371 : 1'h0; // @[implicits.scala 55:10:@28446.4]
  assign _T_1374 = _T_609 & _T_1373; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 351:194:@28447.4]
  assign x484_x247_D20 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@28423.4 package.scala 96:25:@28424.4]
  assign _T_1375 = _T_1374 & x484_x247_D20; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 351:283:@28448.4]
  assign _T_1376 = _T_1375 & x474_b213_D45; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 351:291:@28449.4]
  assign x253_rdrow_number = x253_rdrow_1_io_result; // @[Math.scala 195:22:@28468.4 Math.scala 196:14:@28469.4]
  assign _T_1393 = $signed(x253_rdrow_number); // @[Math.scala 406:49:@28475.4]
  assign _T_1395 = $signed(_T_1393) & $signed(32'sh3); // @[Math.scala 406:56:@28477.4]
  assign _T_1396 = $signed(_T_1395); // @[Math.scala 406:56:@28478.4]
  assign x445_number = $unsigned(_T_1396); // @[implicits.scala 133:21:@28479.4]
  assign x255 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@28493.4 package.scala 96:25:@28494.4]
  assign x486_x230_D1 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@28502.4 package.scala 96:25:@28503.4]
  assign x256 = x255 | x486_x230_D1; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 363:24:@28506.4]
  assign _T_1422 = $signed(x445_number); // @[Math.scala 406:49:@28515.4]
  assign _T_1424 = $signed(_T_1422) & $signed(32'sh3); // @[Math.scala 406:56:@28517.4]
  assign _T_1425 = $signed(_T_1424); // @[Math.scala 406:56:@28518.4]
  assign _T_1429 = $signed(RetimeWrapper_46_io_out); // @[package.scala 96:25:@28526.4]
  assign _T_1433 = x445_number[31]; // @[FixedPoint.scala 50:25:@28533.4]
  assign _T_1437 = _T_1433 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28535.4]
  assign _T_1438 = x445_number[31:2]; // @[FixedPoint.scala 18:52:@28536.4]
  assign _T_1444 = _T_1438 == 30'h3fffffff; // @[Math.scala 451:55:@28538.4]
  assign _T_1445 = x445_number[1:0]; // @[FixedPoint.scala 18:52:@28539.4]
  assign _T_1451 = _T_1445 != 2'h0; // @[Math.scala 451:110:@28541.4]
  assign _T_1452 = _T_1444 & _T_1451; // @[Math.scala 451:94:@28542.4]
  assign _T_1456 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@28550.4 package.scala 96:25:@28551.4]
  assign x259_1_number = _T_1452 ? 32'h0 : _T_1456; // @[Math.scala 454:20:@28552.4]
  assign _GEN_2 = {{9'd0}, x259_1_number}; // @[Math.scala 461:32:@28557.4]
  assign _T_1461 = _GEN_2 << 9; // @[Math.scala 461:32:@28557.4]
  assign _GEN_3 = {{7'd0}, x259_1_number}; // @[Math.scala 461:32:@28562.4]
  assign _T_1464 = _GEN_3 << 7; // @[Math.scala 461:32:@28562.4]
  assign _T_1497 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@28639.4 package.scala 96:25:@28640.4]
  assign _T_1499 = io_rr ? _T_1497 : 1'h0; // @[implicits.scala 55:10:@28641.4]
  assign _T_1500 = _T_609 & _T_1499; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 392:194:@28642.4]
  assign x489_x257_D20 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@28609.4 package.scala 96:25:@28610.4]
  assign _T_1501 = _T_1500 & x489_x257_D20; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 392:283:@28643.4]
  assign _T_1502 = _T_1501 & x474_b213_D45; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 392:291:@28644.4]
  assign x264 = x255 | x236; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 402:59:@28655.4]
  assign _T_1531 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@28699.4 package.scala 96:25:@28700.4]
  assign _T_1533 = io_rr ? _T_1531 : 1'h0; // @[implicits.scala 55:10:@28701.4]
  assign _T_1534 = _T_609 & _T_1533; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 417:194:@28702.4]
  assign x493_x265_D20 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@28687.4 package.scala 96:25:@28688.4]
  assign _T_1535 = _T_1534 & x493_x265_D20; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 417:283:@28703.4]
  assign _T_1536 = _T_1535 & x474_b213_D45; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 417:291:@28704.4]
  assign x269 = x255 | x245; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 421:59:@28715.4]
  assign _T_1560 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@28748.4 package.scala 96:25:@28749.4]
  assign _T_1562 = io_rr ? _T_1560 : 1'h0; // @[implicits.scala 55:10:@28750.4]
  assign _T_1563 = _T_609 & _T_1562; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 432:194:@28751.4]
  assign x494_x270_D20 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@28736.4 package.scala 96:25:@28737.4]
  assign _T_1564 = _T_1563 & x494_x270_D20; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 432:283:@28752.4]
  assign _T_1565 = _T_1564 & x474_b213_D45; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 432:291:@28753.4]
  assign x274_rdrow_number = x274_rdrow_1_io_result; // @[Math.scala 195:22:@28772.4 Math.scala 196:14:@28773.4]
  assign _T_1582 = $signed(x274_rdrow_number); // @[Math.scala 406:49:@28779.4]
  assign _T_1584 = $signed(_T_1582) & $signed(32'sh3); // @[Math.scala 406:56:@28781.4]
  assign _T_1585 = $signed(_T_1584); // @[Math.scala 406:56:@28782.4]
  assign x450_number = $unsigned(_T_1585); // @[implicits.scala 133:21:@28783.4]
  assign x276 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@28797.4 package.scala 96:25:@28798.4]
  assign x277 = x276 | x486_x230_D1; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 442:24:@28801.4]
  assign _T_1608 = $signed(x450_number); // @[Math.scala 406:49:@28810.4]
  assign _T_1610 = $signed(_T_1608) & $signed(32'sh3); // @[Math.scala 406:56:@28812.4]
  assign _T_1611 = $signed(_T_1610); // @[Math.scala 406:56:@28813.4]
  assign _T_1615 = $signed(RetimeWrapper_60_io_out); // @[package.scala 96:25:@28821.4]
  assign _T_1619 = x450_number[31]; // @[FixedPoint.scala 50:25:@28828.4]
  assign _T_1623 = _T_1619 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28830.4]
  assign _T_1624 = x450_number[31:2]; // @[FixedPoint.scala 18:52:@28831.4]
  assign _T_1630 = _T_1624 == 30'h3fffffff; // @[Math.scala 451:55:@28833.4]
  assign _T_1631 = x450_number[1:0]; // @[FixedPoint.scala 18:52:@28834.4]
  assign _T_1637 = _T_1631 != 2'h0; // @[Math.scala 451:110:@28836.4]
  assign _T_1638 = _T_1630 & _T_1637; // @[Math.scala 451:94:@28837.4]
  assign _T_1642 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@28845.4 package.scala 96:25:@28846.4]
  assign x280_1_number = _T_1638 ? 32'h0 : _T_1642; // @[Math.scala 454:20:@28847.4]
  assign _GEN_4 = {{9'd0}, x280_1_number}; // @[Math.scala 461:32:@28852.4]
  assign _T_1647 = _GEN_4 << 9; // @[Math.scala 461:32:@28852.4]
  assign _GEN_5 = {{7'd0}, x280_1_number}; // @[Math.scala 461:32:@28857.4]
  assign _T_1650 = _GEN_5 << 7; // @[Math.scala 461:32:@28857.4]
  assign _T_1680 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@28925.4 package.scala 96:25:@28926.4]
  assign _T_1682 = io_rr ? _T_1680 : 1'h0; // @[implicits.scala 55:10:@28927.4]
  assign _T_1683 = _T_609 & _T_1682; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 469:194:@28928.4]
  assign x497_x278_D20 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@28904.4 package.scala 96:25:@28905.4]
  assign _T_1684 = _T_1683 & x497_x278_D20; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 469:283:@28929.4]
  assign _T_1685 = _T_1684 & x474_b213_D45; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 469:291:@28930.4]
  assign x285 = x276 | x236; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 473:24:@28941.4]
  assign _T_1712 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@28983.4 package.scala 96:25:@28984.4]
  assign _T_1714 = io_rr ? _T_1712 : 1'h0; // @[implicits.scala 55:10:@28985.4]
  assign _T_1715 = _T_609 & _T_1714; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 486:194:@28986.4]
  assign x500_x286_D20 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@28971.4 package.scala 96:25:@28972.4]
  assign _T_1716 = _T_1715 & x500_x286_D20; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 486:283:@28987.4]
  assign _T_1717 = _T_1716 & x474_b213_D45; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 486:291:@28988.4]
  assign x290 = x276 | x245; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 490:24:@28999.4]
  assign _T_1741 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@29032.4 package.scala 96:25:@29033.4]
  assign _T_1743 = io_rr ? _T_1741 : 1'h0; // @[implicits.scala 55:10:@29034.4]
  assign _T_1744 = _T_609 & _T_1743; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 501:194:@29035.4]
  assign x501_x291_D20 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@29020.4 package.scala 96:25:@29021.4]
  assign _T_1745 = _T_1744 & x501_x291_D20; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 501:283:@29036.4]
  assign _T_1746 = _T_1745 & x474_b213_D45; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 501:291:@29037.4]
  assign _T_1873 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@29313.4 package.scala 96:25:@29314.4]
  assign _T_1875 = io_rr ? _T_1873 : 1'h0; // @[implicits.scala 55:10:@29315.4]
  assign x504_b213_D66 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@29304.4 package.scala 96:25:@29305.4]
  assign _T_1876 = _T_1875 & x504_b213_D66; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 563:117:@29316.4]
  assign x503_b214_D66 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@29295.4 package.scala 96:25:@29296.4]
  assign _T_1877 = _T_1876 & x503_b214_D66; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 563:123:@29317.4]
  assign x226_sum_number = x226_sum_1_io_result; // @[Math.scala 154:22:@27452.4 Math.scala 155:14:@27453.4]
  assign x465_x397_D13_number = RetimeWrapper_7_io_out; // @[package.scala 96:25:@27461.4 package.scala 96:25:@27462.4]
  assign x467_x375_D21_number = RetimeWrapper_9_io_out; // @[package.scala 96:25:@27479.4 package.scala 96:25:@27480.4]
  assign x472_x397_D37_number = RetimeWrapper_17_io_out; // @[package.scala 96:25:@27583.4 package.scala 96:25:@27584.4]
  assign x473_x375_D45_number = RetimeWrapper_18_io_out; // @[package.scala 96:25:@27592.4 package.scala 96:25:@27593.4]
  assign x475_x226_sum_D24_number = RetimeWrapper_20_io_out; // @[package.scala 96:25:@27610.4 package.scala 96:25:@27611.4]
  assign x241_sum_number = x241_sum_1_io_result; // @[Math.scala 154:22:@28020.4 Math.scala 155:14:@28021.4]
  assign x482_x422_D13_number = RetimeWrapper_33_io_out; // @[package.scala 96:25:@28038.4 package.scala 96:25:@28039.4]
  assign x250_sum_number = x250_sum_1_io_result; // @[Math.scala 154:22:@28414.4 Math.scala 155:14:@28415.4]
  assign x485_x444_D13_number = RetimeWrapper_42_io_out; // @[package.scala 96:25:@28432.4 package.scala 96:25:@28433.4]
  assign x490_x261_sum_D1_number = RetimeWrapper_51_io_out; // @[package.scala 96:25:@28618.4 package.scala 96:25:@28619.4]
  assign x491_x446_D20_number = RetimeWrapper_52_io_out; // @[package.scala 96:25:@28627.4 package.scala 96:25:@28628.4]
  assign x266_sum_number = x266_sum_1_io_result; // @[Math.scala 154:22:@28678.4 Math.scala 155:14:@28679.4]
  assign x271_sum_number = x271_sum_1_io_result; // @[Math.scala 154:22:@28727.4 Math.scala 155:14:@28728.4]
  assign x496_x451_D20_number = RetimeWrapper_63_io_out; // @[package.scala 96:25:@28895.4 package.scala 96:25:@28896.4]
  assign x498_x282_sum_D1_number = RetimeWrapper_65_io_out; // @[package.scala 96:25:@28913.4 package.scala 96:25:@28914.4]
  assign x287_sum_number = x287_sum_1_io_result; // @[Math.scala 154:22:@28962.4 Math.scala 155:14:@28963.4]
  assign x292_sum_number = x292_sum_1_io_result; // @[Math.scala 154:22:@29011.4 Math.scala 155:14:@29012.4]
  assign io_in_x185_TVALID = _T_1877 & io_sigsIn_backpressure; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 563:22:@29319.4]
  assign io_in_x185_TDATA = {{224'd0}, RetimeWrapper_73_io_out}; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 564:24:@29320.4]
  assign io_in_x184_TREADY = _T_211 & _T_213; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 67:22:@26971.4 sm_x319_inr_Foreach_SAMPLER_BOX.scala 69:22:@26979.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@26949.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@26961.4]
  assign RetimeWrapper_clock = clock; // @[:@26982.4]
  assign RetimeWrapper_reset = reset; // @[:@26983.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26985.4]
  assign RetimeWrapper_io_in = io_in_x184_TDATA[31:0]; // @[package.scala 94:16:@26984.4]
  assign x217_lb_0_clock = clock; // @[:@26992.4]
  assign x217_lb_0_reset = reset; // @[:@26993.4]
  assign x217_lb_0_io_rPort_8_banks_1 = x472_x397_D37_number[1:0]; // @[MemInterfaceType.scala 106:58:@28933.4]
  assign x217_lb_0_io_rPort_8_banks_0 = x496_x451_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@28932.4]
  assign x217_lb_0_io_rPort_8_ofs_0 = x498_x282_sum_D1_number[9:0]; // @[MemInterfaceType.scala 107:54:@28934.4]
  assign x217_lb_0_io_rPort_8_en_0 = _T_1685 & x476_b214_D45; // @[MemInterfaceType.scala 110:79:@28936.4]
  assign x217_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28935.4]
  assign x217_lb_0_io_rPort_7_banks_1 = x482_x422_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@28058.4]
  assign x217_lb_0_io_rPort_7_banks_0 = x473_x375_D45_number[2:0]; // @[MemInterfaceType.scala 106:58:@28057.4]
  assign x217_lb_0_io_rPort_7_ofs_0 = x241_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@28059.4]
  assign x217_lb_0_io_rPort_7_en_0 = _T_1034 & x476_b214_D45; // @[MemInterfaceType.scala 110:79:@28061.4]
  assign x217_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28060.4]
  assign x217_lb_0_io_rPort_6_banks_1 = x472_x397_D37_number[1:0]; // @[MemInterfaceType.scala 106:58:@28647.4]
  assign x217_lb_0_io_rPort_6_banks_0 = x491_x446_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@28646.4]
  assign x217_lb_0_io_rPort_6_ofs_0 = x490_x261_sum_D1_number[9:0]; // @[MemInterfaceType.scala 107:54:@28648.4]
  assign x217_lb_0_io_rPort_6_en_0 = _T_1502 & x476_b214_D45; // @[MemInterfaceType.scala 110:79:@28650.4]
  assign x217_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28649.4]
  assign x217_lb_0_io_rPort_5_banks_1 = x485_x444_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@28756.4]
  assign x217_lb_0_io_rPort_5_banks_0 = x491_x446_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@28755.4]
  assign x217_lb_0_io_rPort_5_ofs_0 = x271_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@28757.4]
  assign x217_lb_0_io_rPort_5_en_0 = _T_1565 & x476_b214_D45; // @[MemInterfaceType.scala 110:79:@28759.4]
  assign x217_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28758.4]
  assign x217_lb_0_io_rPort_4_banks_1 = x482_x422_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@28707.4]
  assign x217_lb_0_io_rPort_4_banks_0 = x491_x446_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@28706.4]
  assign x217_lb_0_io_rPort_4_ofs_0 = x266_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@28708.4]
  assign x217_lb_0_io_rPort_4_en_0 = _T_1536 & x476_b214_D45; // @[MemInterfaceType.scala 110:79:@28710.4]
  assign x217_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28709.4]
  assign x217_lb_0_io_rPort_3_banks_1 = x485_x444_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@28452.4]
  assign x217_lb_0_io_rPort_3_banks_0 = x473_x375_D45_number[2:0]; // @[MemInterfaceType.scala 106:58:@28451.4]
  assign x217_lb_0_io_rPort_3_ofs_0 = x250_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@28453.4]
  assign x217_lb_0_io_rPort_3_en_0 = _T_1376 & x476_b214_D45; // @[MemInterfaceType.scala 110:79:@28455.4]
  assign x217_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28454.4]
  assign x217_lb_0_io_rPort_2_banks_1 = x472_x397_D37_number[1:0]; // @[MemInterfaceType.scala 106:58:@27648.4]
  assign x217_lb_0_io_rPort_2_banks_0 = x473_x375_D45_number[2:0]; // @[MemInterfaceType.scala 106:58:@27647.4]
  assign x217_lb_0_io_rPort_2_ofs_0 = x475_x226_sum_D24_number[9:0]; // @[MemInterfaceType.scala 107:54:@27649.4]
  assign x217_lb_0_io_rPort_2_en_0 = _T_688 & x476_b214_D45; // @[MemInterfaceType.scala 110:79:@27651.4]
  assign x217_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27650.4]
  assign x217_lb_0_io_rPort_1_banks_1 = x485_x444_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@29040.4]
  assign x217_lb_0_io_rPort_1_banks_0 = x496_x451_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@29039.4]
  assign x217_lb_0_io_rPort_1_ofs_0 = x292_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@29041.4]
  assign x217_lb_0_io_rPort_1_en_0 = _T_1746 & x476_b214_D45; // @[MemInterfaceType.scala 110:79:@29043.4]
  assign x217_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@29042.4]
  assign x217_lb_0_io_rPort_0_banks_1 = x482_x422_D13_number[1:0]; // @[MemInterfaceType.scala 106:58:@28991.4]
  assign x217_lb_0_io_rPort_0_banks_0 = x496_x451_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@28990.4]
  assign x217_lb_0_io_rPort_0_ofs_0 = x287_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@28992.4]
  assign x217_lb_0_io_rPort_0_en_0 = _T_1717 & x476_b214_D45; // @[MemInterfaceType.scala 110:79:@28994.4]
  assign x217_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28993.4]
  assign x217_lb_0_io_wPort_0_banks_1 = x465_x397_D13_number[1:0]; // @[MemInterfaceType.scala 88:58:@27518.4]
  assign x217_lb_0_io_wPort_0_banks_0 = x467_x375_D21_number[2:0]; // @[MemInterfaceType.scala 88:58:@27517.4]
  assign x217_lb_0_io_wPort_0_ofs_0 = x226_sum_number[9:0]; // @[MemInterfaceType.scala 89:54:@27519.4]
  assign x217_lb_0_io_wPort_0_data_0 = RetimeWrapper_8_io_out; // @[MemInterfaceType.scala 90:56:@27520.4]
  assign x217_lb_0_io_wPort_0_en_0 = _T_620 & x469_b214_D21; // @[MemInterfaceType.scala 93:57:@27522.4]
  assign x378_sum_1_clock = clock; // @[:@27117.4]
  assign x378_sum_1_reset = reset; // @[:@27118.4]
  assign x378_sum_1_io_a = _T_280 ? 32'h0 : _T_282; // @[Math.scala 151:17:@27119.4]
  assign x378_sum_1_io_b = $unsigned(_T_295); // @[Math.scala 152:17:@27120.4]
  assign x378_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@27121.4]
  assign x381_sum_1_clock = clock; // @[:@27155.4]
  assign x381_sum_1_reset = reset; // @[:@27156.4]
  assign x381_sum_1_io_a = _T_321 ? 32'h0 : _T_323; // @[Math.scala 151:17:@27157.4]
  assign x381_sum_1_io_b = $unsigned(_T_336); // @[Math.scala 152:17:@27158.4]
  assign x381_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@27159.4]
  assign x384_sum_1_clock = clock; // @[:@27193.4]
  assign x384_sum_1_reset = reset; // @[:@27194.4]
  assign x384_sum_1_io_a = _T_362 ? 32'h0 : _T_364; // @[Math.scala 151:17:@27195.4]
  assign x384_sum_1_io_b = $unsigned(_T_377); // @[Math.scala 152:17:@27196.4]
  assign x384_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@27197.4]
  assign x387_sum_1_clock = clock; // @[:@27231.4]
  assign x387_sum_1_reset = reset; // @[:@27232.4]
  assign x387_sum_1_io_a = _T_403 ? 32'h0 : _T_405; // @[Math.scala 151:17:@27233.4]
  assign x387_sum_1_io_b = $unsigned(_T_418); // @[Math.scala 152:17:@27234.4]
  assign x387_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@27235.4]
  assign RetimeWrapper_1_clock = clock; // @[:@27254.4]
  assign RetimeWrapper_1_reset = reset; // @[:@27255.4]
  assign RetimeWrapper_1_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@27257.4]
  assign RetimeWrapper_1_io_in = {_T_429,_T_430}; // @[package.scala 94:16:@27256.4]
  assign RetimeWrapper_2_clock = clock; // @[:@27272.4]
  assign RetimeWrapper_2_reset = reset; // @[:@27273.4]
  assign RetimeWrapper_2_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@27276.4]
  assign RetimeWrapper_2_io_in = $unsigned(_T_461); // @[package.scala 94:16:@27275.4]
  assign x390_sum_1_clock = clock; // @[:@27285.4]
  assign x390_sum_1_reset = reset; // @[:@27286.4]
  assign x390_sum_1_io_a = _T_444 ? 32'h0 : _T_448; // @[Math.scala 151:17:@27287.4]
  assign x390_sum_1_io_b = $unsigned(_T_465); // @[Math.scala 152:17:@27288.4]
  assign x390_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@27289.4]
  assign x393_sum_1_clock = clock; // @[:@27323.4]
  assign x393_sum_1_reset = reset; // @[:@27324.4]
  assign x393_sum_1_io_a = _T_491 ? 32'h0 : _T_493; // @[Math.scala 151:17:@27325.4]
  assign x393_sum_1_io_b = $unsigned(_T_506); // @[Math.scala 152:17:@27326.4]
  assign x393_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@27327.4]
  assign x396_sub_1_clock = clock; // @[:@27349.4]
  assign x396_sub_1_reset = reset; // @[:@27350.4]
  assign x396_sub_1_io_a = x393_sum_1_io_result; // @[Math.scala 192:17:@27351.4]
  assign x396_sub_1_io_b = 32'h3; // @[Math.scala 193:17:@27352.4]
  assign x396_sub_1_io_flow = io_in_x185_TREADY; // @[Math.scala 194:20:@27353.4]
  assign RetimeWrapper_3_clock = clock; // @[:@27359.4]
  assign RetimeWrapper_3_reset = reset; // @[:@27360.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27362.4]
  assign RetimeWrapper_3_io_in = $signed(_T_516) < $signed(32'sh6); // @[package.scala 94:16:@27361.4]
  assign RetimeWrapper_4_clock = clock; // @[:@27368.4]
  assign RetimeWrapper_4_reset = reset; // @[:@27369.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27371.4]
  assign RetimeWrapper_4_io_in = $signed(_T_516) < $signed(32'sh3); // @[package.scala 94:16:@27370.4]
  assign RetimeWrapper_5_clock = clock; // @[:@27377.4]
  assign RetimeWrapper_5_reset = reset; // @[:@27378.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27380.4]
  assign RetimeWrapper_5_io_in = x393_sum_1_io_result; // @[package.scala 94:16:@27379.4]
  assign x400_sum_1_clock = clock; // @[:@27416.4]
  assign x400_sum_1_reset = reset; // @[:@27417.4]
  assign x400_sum_1_io_a = _T_573[31:0]; // @[Math.scala 151:17:@27418.4]
  assign x400_sum_1_io_b = _T_576[31:0]; // @[Math.scala 152:17:@27419.4]
  assign x400_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@27420.4]
  assign x225_div_1_clock = clock; // @[:@27428.4]
  assign x225_div_1_io_a = __1_io_result; // @[Math.scala 328:17:@27430.4]
  assign x225_div_1_io_flow = io_in_x185_TREADY; // @[Math.scala 330:20:@27432.4]
  assign RetimeWrapper_6_clock = clock; // @[:@27438.4]
  assign RetimeWrapper_6_reset = reset; // @[:@27439.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27441.4]
  assign RetimeWrapper_6_io_in = x400_sum_1_io_result; // @[package.scala 94:16:@27440.4]
  assign x226_sum_1_clock = clock; // @[:@27447.4]
  assign x226_sum_1_reset = reset; // @[:@27448.4]
  assign x226_sum_1_io_a = RetimeWrapper_6_io_out; // @[Math.scala 151:17:@27449.4]
  assign x226_sum_1_io_b = x225_div_1_io_result; // @[Math.scala 152:17:@27450.4]
  assign x226_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@27451.4]
  assign RetimeWrapper_7_clock = clock; // @[:@27457.4]
  assign RetimeWrapper_7_reset = reset; // @[:@27458.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27460.4]
  assign RetimeWrapper_7_io_in = x462_x394_D1 ? x463_x393_sum_D1_number : x396_sub_number; // @[package.scala 94:16:@27459.4]
  assign RetimeWrapper_8_clock = clock; // @[:@27466.4]
  assign RetimeWrapper_8_reset = reset; // @[:@27467.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27469.4]
  assign RetimeWrapper_8_io_in = RetimeWrapper_io_out; // @[package.scala 94:16:@27468.4]
  assign RetimeWrapper_9_clock = clock; // @[:@27475.4]
  assign RetimeWrapper_9_reset = reset; // @[:@27476.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27478.4]
  assign RetimeWrapper_9_io_in = $unsigned(_T_257); // @[package.scala 94:16:@27477.4]
  assign RetimeWrapper_10_clock = clock; // @[:@27484.4]
  assign RetimeWrapper_10_reset = reset; // @[:@27485.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27487.4]
  assign RetimeWrapper_10_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@27486.4]
  assign RetimeWrapper_11_clock = clock; // @[:@27493.4]
  assign RetimeWrapper_11_reset = reset; // @[:@27494.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27496.4]
  assign RetimeWrapper_11_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@27495.4]
  assign RetimeWrapper_12_clock = clock; // @[:@27504.4]
  assign RetimeWrapper_12_reset = reset; // @[:@27505.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27507.4]
  assign RetimeWrapper_12_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27506.4]
  assign RetimeWrapper_13_clock = clock; // @[:@27525.4]
  assign RetimeWrapper_13_reset = reset; // @[:@27526.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27528.4]
  assign RetimeWrapper_13_io_in = __io_result; // @[package.scala 94:16:@27527.4]
  assign RetimeWrapper_14_clock = clock; // @[:@27539.4]
  assign RetimeWrapper_14_reset = reset; // @[:@27540.4]
  assign RetimeWrapper_14_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@27542.4]
  assign RetimeWrapper_14_io_in = $signed(_T_630) < $signed(32'sh0); // @[package.scala 94:16:@27541.4]
  assign RetimeWrapper_15_clock = clock; // @[:@27548.4]
  assign RetimeWrapper_15_reset = reset; // @[:@27549.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27551.4]
  assign RetimeWrapper_15_io_in = __1_io_result; // @[package.scala 94:16:@27550.4]
  assign RetimeWrapper_16_clock = clock; // @[:@27564.4]
  assign RetimeWrapper_16_reset = reset; // @[:@27565.4]
  assign RetimeWrapper_16_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@27567.4]
  assign RetimeWrapper_16_io_in = $signed(_T_645) < $signed(32'sh0); // @[package.scala 94:16:@27566.4]
  assign RetimeWrapper_17_clock = clock; // @[:@27579.4]
  assign RetimeWrapper_17_reset = reset; // @[:@27580.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27582.4]
  assign RetimeWrapper_17_io_in = x462_x394_D1 ? x463_x393_sum_D1_number : x396_sub_number; // @[package.scala 94:16:@27581.4]
  assign RetimeWrapper_18_clock = clock; // @[:@27588.4]
  assign RetimeWrapper_18_reset = reset; // @[:@27589.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27591.4]
  assign RetimeWrapper_18_io_in = $unsigned(_T_257); // @[package.scala 94:16:@27590.4]
  assign RetimeWrapper_19_clock = clock; // @[:@27597.4]
  assign RetimeWrapper_19_reset = reset; // @[:@27598.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27600.4]
  assign RetimeWrapper_19_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@27599.4]
  assign RetimeWrapper_20_clock = clock; // @[:@27606.4]
  assign RetimeWrapper_20_reset = reset; // @[:@27607.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27609.4]
  assign RetimeWrapper_20_io_in = x226_sum_1_io_result; // @[package.scala 94:16:@27608.4]
  assign RetimeWrapper_21_clock = clock; // @[:@27615.4]
  assign RetimeWrapper_21_reset = reset; // @[:@27616.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27618.4]
  assign RetimeWrapper_21_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@27617.4]
  assign RetimeWrapper_22_clock = clock; // @[:@27624.4]
  assign RetimeWrapper_22_reset = reset; // @[:@27625.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27627.4]
  assign RetimeWrapper_22_io_in = ~ x231; // @[package.scala 94:16:@27626.4]
  assign RetimeWrapper_23_clock = clock; // @[:@27636.4]
  assign RetimeWrapper_23_reset = reset; // @[:@27637.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27639.4]
  assign RetimeWrapper_23_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27638.4]
  assign x235_rdcol_1_clock = clock; // @[:@27659.4]
  assign x235_rdcol_1_reset = reset; // @[:@27660.4]
  assign x235_rdcol_1_io_a = RetimeWrapper_15_io_out; // @[Math.scala 192:17:@27661.4]
  assign x235_rdcol_1_io_b = 32'h1; // @[Math.scala 193:17:@27662.4]
  assign x235_rdcol_1_io_flow = io_in_x185_TREADY; // @[Math.scala 194:20:@27663.4]
  assign RetimeWrapper_24_clock = clock; // @[:@27674.4]
  assign RetimeWrapper_24_reset = reset; // @[:@27675.4]
  assign RetimeWrapper_24_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@27677.4]
  assign RetimeWrapper_24_io_in = $signed(_T_703) < $signed(32'sh0); // @[package.scala 94:16:@27676.4]
  assign RetimeWrapper_25_clock = clock; // @[:@27683.4]
  assign RetimeWrapper_25_reset = reset; // @[:@27684.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27686.4]
  assign RetimeWrapper_25_io_in = RetimeWrapper_14_io_out; // @[package.scala 94:16:@27685.4]
  assign x403_sum_1_clock = clock; // @[:@27726.4]
  assign x403_sum_1_reset = reset; // @[:@27727.4]
  assign x403_sum_1_io_a = _T_736 ? 32'h0 : _T_738; // @[Math.scala 151:17:@27728.4]
  assign x403_sum_1_io_b = $unsigned(_T_751); // @[Math.scala 152:17:@27729.4]
  assign x403_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@27730.4]
  assign RetimeWrapper_26_clock = clock; // @[:@27749.4]
  assign RetimeWrapper_26_reset = reset; // @[:@27750.4]
  assign RetimeWrapper_26_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@27752.4]
  assign RetimeWrapper_26_io_in = {_T_762,_T_763}; // @[package.scala 94:16:@27751.4]
  assign RetimeWrapper_27_clock = clock; // @[:@27767.4]
  assign RetimeWrapper_27_reset = reset; // @[:@27768.4]
  assign RetimeWrapper_27_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@27771.4]
  assign RetimeWrapper_27_io_in = $unsigned(_T_794); // @[package.scala 94:16:@27770.4]
  assign x406_sum_1_clock = clock; // @[:@27780.4]
  assign x406_sum_1_reset = reset; // @[:@27781.4]
  assign x406_sum_1_io_a = _T_777 ? 32'h0 : _T_781; // @[Math.scala 151:17:@27782.4]
  assign x406_sum_1_io_b = $unsigned(_T_798); // @[Math.scala 152:17:@27783.4]
  assign x406_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@27784.4]
  assign x409_sum_1_clock = clock; // @[:@27818.4]
  assign x409_sum_1_reset = reset; // @[:@27819.4]
  assign x409_sum_1_io_a = _T_824 ? 32'h0 : _T_826; // @[Math.scala 151:17:@27820.4]
  assign x409_sum_1_io_b = $unsigned(_T_839); // @[Math.scala 152:17:@27821.4]
  assign x409_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@27822.4]
  assign x412_sum_1_clock = clock; // @[:@27856.4]
  assign x412_sum_1_reset = reset; // @[:@27857.4]
  assign x412_sum_1_io_a = _T_865 ? 32'h0 : _T_867; // @[Math.scala 151:17:@27858.4]
  assign x412_sum_1_io_b = $unsigned(_T_880); // @[Math.scala 152:17:@27859.4]
  assign x412_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@27860.4]
  assign x415_sum_1_clock = clock; // @[:@27894.4]
  assign x415_sum_1_reset = reset; // @[:@27895.4]
  assign x415_sum_1_io_a = _T_906 ? 32'h0 : _T_908; // @[Math.scala 151:17:@27896.4]
  assign x415_sum_1_io_b = $unsigned(_T_921); // @[Math.scala 152:17:@27897.4]
  assign x415_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@27898.4]
  assign x418_sum_1_clock = clock; // @[:@27932.4]
  assign x418_sum_1_reset = reset; // @[:@27933.4]
  assign x418_sum_1_io_a = _T_947 ? 32'h0 : _T_949; // @[Math.scala 151:17:@27934.4]
  assign x418_sum_1_io_b = $unsigned(_T_962); // @[Math.scala 152:17:@27935.4]
  assign x418_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@27936.4]
  assign RetimeWrapper_28_clock = clock; // @[:@27947.4]
  assign RetimeWrapper_28_reset = reset; // @[:@27948.4]
  assign RetimeWrapper_28_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@27950.4]
  assign RetimeWrapper_28_io_in = $signed(_T_972) < $signed(32'sh3); // @[package.scala 94:16:@27949.4]
  assign RetimeWrapper_29_clock = clock; // @[:@27961.4]
  assign RetimeWrapper_29_reset = reset; // @[:@27962.4]
  assign RetimeWrapper_29_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@27964.4]
  assign RetimeWrapper_29_io_in = $signed(_T_972) < $signed(32'sh6); // @[package.scala 94:16:@27963.4]
  assign x421_sub_1_clock = clock; // @[:@27972.4]
  assign x421_sub_1_reset = reset; // @[:@27973.4]
  assign x421_sub_1_io_a = x418_sum_1_io_result; // @[Math.scala 192:17:@27974.4]
  assign x421_sub_1_io_b = 32'h3; // @[Math.scala 193:17:@27975.4]
  assign x421_sub_1_io_flow = io_in_x185_TREADY; // @[Math.scala 194:20:@27976.4]
  assign RetimeWrapper_30_clock = clock; // @[:@27982.4]
  assign RetimeWrapper_30_reset = reset; // @[:@27983.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27985.4]
  assign RetimeWrapper_30_io_in = x418_sum_1_io_result; // @[package.scala 94:16:@27984.4]
  assign x240_div_1_clock = clock; // @[:@27996.4]
  assign x240_div_1_io_a = x235_rdcol_1_io_result; // @[Math.scala 328:17:@27998.4]
  assign x240_div_1_io_flow = io_in_x185_TREADY; // @[Math.scala 330:20:@28000.4]
  assign RetimeWrapper_31_clock = clock; // @[:@28006.4]
  assign RetimeWrapper_31_reset = reset; // @[:@28007.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28009.4]
  assign RetimeWrapper_31_io_in = x400_sum_1_io_result; // @[package.scala 94:16:@28008.4]
  assign x241_sum_1_clock = clock; // @[:@28015.4]
  assign x241_sum_1_reset = reset; // @[:@28016.4]
  assign x241_sum_1_io_a = RetimeWrapper_31_io_out; // @[Math.scala 151:17:@28017.4]
  assign x241_sum_1_io_b = x240_div_1_io_result; // @[Math.scala 152:17:@28018.4]
  assign x241_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@28019.4]
  assign RetimeWrapper_32_clock = clock; // @[:@28025.4]
  assign RetimeWrapper_32_reset = reset; // @[:@28026.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28028.4]
  assign RetimeWrapper_32_io_in = ~ x237; // @[package.scala 94:16:@28027.4]
  assign RetimeWrapper_33_clock = clock; // @[:@28034.4]
  assign RetimeWrapper_33_reset = reset; // @[:@28035.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28037.4]
  assign RetimeWrapper_33_io_in = x419 ? x479_x418_sum_D1_number : x421_sub_number; // @[package.scala 94:16:@28036.4]
  assign RetimeWrapper_34_clock = clock; // @[:@28046.4]
  assign RetimeWrapper_34_reset = reset; // @[:@28047.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28049.4]
  assign RetimeWrapper_34_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28048.4]
  assign x244_rdcol_1_clock = clock; // @[:@28069.4]
  assign x244_rdcol_1_reset = reset; // @[:@28070.4]
  assign x244_rdcol_1_io_a = RetimeWrapper_15_io_out; // @[Math.scala 192:17:@28071.4]
  assign x244_rdcol_1_io_b = 32'h2; // @[Math.scala 193:17:@28072.4]
  assign x244_rdcol_1_io_flow = io_in_x185_TREADY; // @[Math.scala 194:20:@28073.4]
  assign RetimeWrapper_35_clock = clock; // @[:@28084.4]
  assign RetimeWrapper_35_reset = reset; // @[:@28085.4]
  assign RetimeWrapper_35_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@28087.4]
  assign RetimeWrapper_35_io_in = $signed(_T_1049) < $signed(32'sh0); // @[package.scala 94:16:@28086.4]
  assign x425_sum_1_clock = clock; // @[:@28129.4]
  assign x425_sum_1_reset = reset; // @[:@28130.4]
  assign x425_sum_1_io_a = _T_1081 ? 32'h0 : _T_1083; // @[Math.scala 151:17:@28131.4]
  assign x425_sum_1_io_b = $unsigned(_T_1096); // @[Math.scala 152:17:@28132.4]
  assign x425_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@28133.4]
  assign RetimeWrapper_36_clock = clock; // @[:@28152.4]
  assign RetimeWrapper_36_reset = reset; // @[:@28153.4]
  assign RetimeWrapper_36_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@28155.4]
  assign RetimeWrapper_36_io_in = {_T_1107,_T_1108}; // @[package.scala 94:16:@28154.4]
  assign RetimeWrapper_37_clock = clock; // @[:@28170.4]
  assign RetimeWrapper_37_reset = reset; // @[:@28171.4]
  assign RetimeWrapper_37_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@28174.4]
  assign RetimeWrapper_37_io_in = $unsigned(_T_1139); // @[package.scala 94:16:@28173.4]
  assign x428_sum_1_clock = clock; // @[:@28183.4]
  assign x428_sum_1_reset = reset; // @[:@28184.4]
  assign x428_sum_1_io_a = _T_1122 ? 32'h0 : _T_1126; // @[Math.scala 151:17:@28185.4]
  assign x428_sum_1_io_b = $unsigned(_T_1143); // @[Math.scala 152:17:@28186.4]
  assign x428_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@28187.4]
  assign x431_sum_1_clock = clock; // @[:@28221.4]
  assign x431_sum_1_reset = reset; // @[:@28222.4]
  assign x431_sum_1_io_a = _T_1169 ? 32'h0 : _T_1171; // @[Math.scala 151:17:@28223.4]
  assign x431_sum_1_io_b = $unsigned(_T_1184); // @[Math.scala 152:17:@28224.4]
  assign x431_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@28225.4]
  assign x434_sum_1_clock = clock; // @[:@28259.4]
  assign x434_sum_1_reset = reset; // @[:@28260.4]
  assign x434_sum_1_io_a = _T_1210 ? 32'h0 : _T_1212; // @[Math.scala 151:17:@28261.4]
  assign x434_sum_1_io_b = $unsigned(_T_1225); // @[Math.scala 152:17:@28262.4]
  assign x434_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@28263.4]
  assign x437_sum_1_clock = clock; // @[:@28297.4]
  assign x437_sum_1_reset = reset; // @[:@28298.4]
  assign x437_sum_1_io_a = _T_1251 ? 32'h0 : _T_1253; // @[Math.scala 151:17:@28299.4]
  assign x437_sum_1_io_b = $unsigned(_T_1266); // @[Math.scala 152:17:@28300.4]
  assign x437_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@28301.4]
  assign x440_sum_1_clock = clock; // @[:@28335.4]
  assign x440_sum_1_reset = reset; // @[:@28336.4]
  assign x440_sum_1_io_a = _T_1292 ? 32'h0 : _T_1294; // @[Math.scala 151:17:@28337.4]
  assign x440_sum_1_io_b = $unsigned(_T_1307); // @[Math.scala 152:17:@28338.4]
  assign x440_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@28339.4]
  assign RetimeWrapper_38_clock = clock; // @[:@28350.4]
  assign RetimeWrapper_38_reset = reset; // @[:@28351.4]
  assign RetimeWrapper_38_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@28353.4]
  assign RetimeWrapper_38_io_in = $signed(_T_1317) < $signed(32'sh3); // @[package.scala 94:16:@28352.4]
  assign RetimeWrapper_39_clock = clock; // @[:@28364.4]
  assign RetimeWrapper_39_reset = reset; // @[:@28365.4]
  assign RetimeWrapper_39_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@28367.4]
  assign RetimeWrapper_39_io_in = $signed(_T_1317) < $signed(32'sh6); // @[package.scala 94:16:@28366.4]
  assign x443_sub_1_clock = clock; // @[:@28375.4]
  assign x443_sub_1_reset = reset; // @[:@28376.4]
  assign x443_sub_1_io_a = x440_sum_1_io_result; // @[Math.scala 192:17:@28377.4]
  assign x443_sub_1_io_b = 32'h3; // @[Math.scala 193:17:@28378.4]
  assign x443_sub_1_io_flow = io_in_x185_TREADY; // @[Math.scala 194:20:@28379.4]
  assign RetimeWrapper_40_clock = clock; // @[:@28385.4]
  assign RetimeWrapper_40_reset = reset; // @[:@28386.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28388.4]
  assign RetimeWrapper_40_io_in = x440_sum_1_io_result; // @[package.scala 94:16:@28387.4]
  assign x249_div_1_clock = clock; // @[:@28399.4]
  assign x249_div_1_io_a = x244_rdcol_1_io_result; // @[Math.scala 328:17:@28401.4]
  assign x249_div_1_io_flow = io_in_x185_TREADY; // @[Math.scala 330:20:@28403.4]
  assign x250_sum_1_clock = clock; // @[:@28409.4]
  assign x250_sum_1_reset = reset; // @[:@28410.4]
  assign x250_sum_1_io_a = RetimeWrapper_31_io_out; // @[Math.scala 151:17:@28411.4]
  assign x250_sum_1_io_b = x249_div_1_io_result; // @[Math.scala 152:17:@28412.4]
  assign x250_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@28413.4]
  assign RetimeWrapper_41_clock = clock; // @[:@28419.4]
  assign RetimeWrapper_41_reset = reset; // @[:@28420.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28422.4]
  assign RetimeWrapper_41_io_in = ~ x246; // @[package.scala 94:16:@28421.4]
  assign RetimeWrapper_42_clock = clock; // @[:@28428.4]
  assign RetimeWrapper_42_reset = reset; // @[:@28429.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28431.4]
  assign RetimeWrapper_42_io_in = x441 ? x483_x440_sum_D1_number : x443_sub_number; // @[package.scala 94:16:@28430.4]
  assign RetimeWrapper_43_clock = clock; // @[:@28440.4]
  assign RetimeWrapper_43_reset = reset; // @[:@28441.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28443.4]
  assign RetimeWrapper_43_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28442.4]
  assign x253_rdrow_1_clock = clock; // @[:@28463.4]
  assign x253_rdrow_1_reset = reset; // @[:@28464.4]
  assign x253_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@28465.4]
  assign x253_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@28466.4]
  assign x253_rdrow_1_io_flow = io_in_x185_TREADY; // @[Math.scala 194:20:@28467.4]
  assign RetimeWrapper_44_clock = clock; // @[:@28489.4]
  assign RetimeWrapper_44_reset = reset; // @[:@28490.4]
  assign RetimeWrapper_44_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@28492.4]
  assign RetimeWrapper_44_io_in = $signed(_T_1393) < $signed(32'sh0); // @[package.scala 94:16:@28491.4]
  assign RetimeWrapper_45_clock = clock; // @[:@28498.4]
  assign RetimeWrapper_45_reset = reset; // @[:@28499.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28501.4]
  assign RetimeWrapper_45_io_in = RetimeWrapper_16_io_out; // @[package.scala 94:16:@28500.4]
  assign RetimeWrapper_46_clock = clock; // @[:@28520.4]
  assign RetimeWrapper_46_reset = reset; // @[:@28521.4]
  assign RetimeWrapper_46_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@28524.4]
  assign RetimeWrapper_46_io_in = $unsigned(_T_1425); // @[package.scala 94:16:@28523.4]
  assign RetimeWrapper_47_clock = clock; // @[:@28546.4]
  assign RetimeWrapper_47_reset = reset; // @[:@28547.4]
  assign RetimeWrapper_47_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@28549.4]
  assign RetimeWrapper_47_io_in = {_T_1437,_T_1438}; // @[package.scala 94:16:@28548.4]
  assign x449_sum_1_clock = clock; // @[:@28567.4]
  assign x449_sum_1_reset = reset; // @[:@28568.4]
  assign x449_sum_1_io_a = _T_1461[31:0]; // @[Math.scala 151:17:@28569.4]
  assign x449_sum_1_io_b = _T_1464[31:0]; // @[Math.scala 152:17:@28570.4]
  assign x449_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@28571.4]
  assign RetimeWrapper_48_clock = clock; // @[:@28577.4]
  assign RetimeWrapper_48_reset = reset; // @[:@28578.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28580.4]
  assign RetimeWrapper_48_io_in = x225_div_1_io_result; // @[package.scala 94:16:@28579.4]
  assign RetimeWrapper_49_clock = clock; // @[:@28586.4]
  assign RetimeWrapper_49_reset = reset; // @[:@28587.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28589.4]
  assign RetimeWrapper_49_io_in = x449_sum_1_io_result; // @[package.scala 94:16:@28588.4]
  assign x261_sum_1_clock = clock; // @[:@28595.4]
  assign x261_sum_1_reset = reset; // @[:@28596.4]
  assign x261_sum_1_io_a = RetimeWrapper_49_io_out; // @[Math.scala 151:17:@28597.4]
  assign x261_sum_1_io_b = RetimeWrapper_48_io_out; // @[Math.scala 152:17:@28598.4]
  assign x261_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@28599.4]
  assign RetimeWrapper_50_clock = clock; // @[:@28605.4]
  assign RetimeWrapper_50_reset = reset; // @[:@28606.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28608.4]
  assign RetimeWrapper_50_io_in = ~ x256; // @[package.scala 94:16:@28607.4]
  assign RetimeWrapper_51_clock = clock; // @[:@28614.4]
  assign RetimeWrapper_51_reset = reset; // @[:@28615.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28617.4]
  assign RetimeWrapper_51_io_in = x261_sum_1_io_result; // @[package.scala 94:16:@28616.4]
  assign RetimeWrapper_52_clock = clock; // @[:@28623.4]
  assign RetimeWrapper_52_reset = reset; // @[:@28624.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28626.4]
  assign RetimeWrapper_52_io_in = $unsigned(_T_1429); // @[package.scala 94:16:@28625.4]
  assign RetimeWrapper_53_clock = clock; // @[:@28635.4]
  assign RetimeWrapper_53_reset = reset; // @[:@28636.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28638.4]
  assign RetimeWrapper_53_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28637.4]
  assign RetimeWrapper_54_clock = clock; // @[:@28662.4]
  assign RetimeWrapper_54_reset = reset; // @[:@28663.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28665.4]
  assign RetimeWrapper_54_io_in = x449_sum_1_io_result; // @[package.scala 94:16:@28664.4]
  assign x266_sum_1_clock = clock; // @[:@28673.4]
  assign x266_sum_1_reset = reset; // @[:@28674.4]
  assign x266_sum_1_io_a = RetimeWrapper_54_io_out; // @[Math.scala 151:17:@28675.4]
  assign x266_sum_1_io_b = x240_div_1_io_result; // @[Math.scala 152:17:@28676.4]
  assign x266_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@28677.4]
  assign RetimeWrapper_55_clock = clock; // @[:@28683.4]
  assign RetimeWrapper_55_reset = reset; // @[:@28684.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28686.4]
  assign RetimeWrapper_55_io_in = ~ x264; // @[package.scala 94:16:@28685.4]
  assign RetimeWrapper_56_clock = clock; // @[:@28695.4]
  assign RetimeWrapper_56_reset = reset; // @[:@28696.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28698.4]
  assign RetimeWrapper_56_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28697.4]
  assign x271_sum_1_clock = clock; // @[:@28722.4]
  assign x271_sum_1_reset = reset; // @[:@28723.4]
  assign x271_sum_1_io_a = RetimeWrapper_54_io_out; // @[Math.scala 151:17:@28724.4]
  assign x271_sum_1_io_b = x249_div_1_io_result; // @[Math.scala 152:17:@28725.4]
  assign x271_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@28726.4]
  assign RetimeWrapper_57_clock = clock; // @[:@28732.4]
  assign RetimeWrapper_57_reset = reset; // @[:@28733.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28735.4]
  assign RetimeWrapper_57_io_in = ~ x269; // @[package.scala 94:16:@28734.4]
  assign RetimeWrapper_58_clock = clock; // @[:@28744.4]
  assign RetimeWrapper_58_reset = reset; // @[:@28745.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28747.4]
  assign RetimeWrapper_58_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28746.4]
  assign x274_rdrow_1_clock = clock; // @[:@28767.4]
  assign x274_rdrow_1_reset = reset; // @[:@28768.4]
  assign x274_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@28769.4]
  assign x274_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@28770.4]
  assign x274_rdrow_1_io_flow = io_in_x185_TREADY; // @[Math.scala 194:20:@28771.4]
  assign RetimeWrapper_59_clock = clock; // @[:@28793.4]
  assign RetimeWrapper_59_reset = reset; // @[:@28794.4]
  assign RetimeWrapper_59_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@28796.4]
  assign RetimeWrapper_59_io_in = $signed(_T_1582) < $signed(32'sh0); // @[package.scala 94:16:@28795.4]
  assign RetimeWrapper_60_clock = clock; // @[:@28815.4]
  assign RetimeWrapper_60_reset = reset; // @[:@28816.4]
  assign RetimeWrapper_60_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@28819.4]
  assign RetimeWrapper_60_io_in = $unsigned(_T_1611); // @[package.scala 94:16:@28818.4]
  assign RetimeWrapper_61_clock = clock; // @[:@28841.4]
  assign RetimeWrapper_61_reset = reset; // @[:@28842.4]
  assign RetimeWrapper_61_io_flow = io_in_x185_TREADY; // @[package.scala 95:18:@28844.4]
  assign RetimeWrapper_61_io_in = {_T_1623,_T_1624}; // @[package.scala 94:16:@28843.4]
  assign x454_sum_1_clock = clock; // @[:@28862.4]
  assign x454_sum_1_reset = reset; // @[:@28863.4]
  assign x454_sum_1_io_a = _T_1647[31:0]; // @[Math.scala 151:17:@28864.4]
  assign x454_sum_1_io_b = _T_1650[31:0]; // @[Math.scala 152:17:@28865.4]
  assign x454_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@28866.4]
  assign RetimeWrapper_62_clock = clock; // @[:@28872.4]
  assign RetimeWrapper_62_reset = reset; // @[:@28873.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28875.4]
  assign RetimeWrapper_62_io_in = x454_sum_1_io_result; // @[package.scala 94:16:@28874.4]
  assign x282_sum_1_clock = clock; // @[:@28881.4]
  assign x282_sum_1_reset = reset; // @[:@28882.4]
  assign x282_sum_1_io_a = RetimeWrapper_62_io_out; // @[Math.scala 151:17:@28883.4]
  assign x282_sum_1_io_b = RetimeWrapper_48_io_out; // @[Math.scala 152:17:@28884.4]
  assign x282_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@28885.4]
  assign RetimeWrapper_63_clock = clock; // @[:@28891.4]
  assign RetimeWrapper_63_reset = reset; // @[:@28892.4]
  assign RetimeWrapper_63_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28894.4]
  assign RetimeWrapper_63_io_in = $unsigned(_T_1615); // @[package.scala 94:16:@28893.4]
  assign RetimeWrapper_64_clock = clock; // @[:@28900.4]
  assign RetimeWrapper_64_reset = reset; // @[:@28901.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28903.4]
  assign RetimeWrapper_64_io_in = ~ x277; // @[package.scala 94:16:@28902.4]
  assign RetimeWrapper_65_clock = clock; // @[:@28909.4]
  assign RetimeWrapper_65_reset = reset; // @[:@28910.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28912.4]
  assign RetimeWrapper_65_io_in = x282_sum_1_io_result; // @[package.scala 94:16:@28911.4]
  assign RetimeWrapper_66_clock = clock; // @[:@28921.4]
  assign RetimeWrapper_66_reset = reset; // @[:@28922.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28924.4]
  assign RetimeWrapper_66_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28923.4]
  assign RetimeWrapper_67_clock = clock; // @[:@28948.4]
  assign RetimeWrapper_67_reset = reset; // @[:@28949.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28951.4]
  assign RetimeWrapper_67_io_in = x454_sum_1_io_result; // @[package.scala 94:16:@28950.4]
  assign x287_sum_1_clock = clock; // @[:@28957.4]
  assign x287_sum_1_reset = reset; // @[:@28958.4]
  assign x287_sum_1_io_a = RetimeWrapper_67_io_out; // @[Math.scala 151:17:@28959.4]
  assign x287_sum_1_io_b = x240_div_1_io_result; // @[Math.scala 152:17:@28960.4]
  assign x287_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@28961.4]
  assign RetimeWrapper_68_clock = clock; // @[:@28967.4]
  assign RetimeWrapper_68_reset = reset; // @[:@28968.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28970.4]
  assign RetimeWrapper_68_io_in = ~ x285; // @[package.scala 94:16:@28969.4]
  assign RetimeWrapper_69_clock = clock; // @[:@28979.4]
  assign RetimeWrapper_69_reset = reset; // @[:@28980.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28982.4]
  assign RetimeWrapper_69_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28981.4]
  assign x292_sum_1_clock = clock; // @[:@29006.4]
  assign x292_sum_1_reset = reset; // @[:@29007.4]
  assign x292_sum_1_io_a = RetimeWrapper_67_io_out; // @[Math.scala 151:17:@29008.4]
  assign x292_sum_1_io_b = x249_div_1_io_result; // @[Math.scala 152:17:@29009.4]
  assign x292_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@29010.4]
  assign RetimeWrapper_70_clock = clock; // @[:@29016.4]
  assign RetimeWrapper_70_reset = reset; // @[:@29017.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29019.4]
  assign RetimeWrapper_70_io_in = ~ x290; // @[package.scala 94:16:@29018.4]
  assign RetimeWrapper_71_clock = clock; // @[:@29028.4]
  assign RetimeWrapper_71_reset = reset; // @[:@29029.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29031.4]
  assign RetimeWrapper_71_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@29030.4]
  assign x295_1_clock = clock; // @[:@29051.4]
  assign x295_1_io_a = x217_lb_0_io_rPort_2_output_0; // @[Math.scala 263:17:@29053.4]
  assign x295_1_io_b = 32'h1; // @[Math.scala 264:17:@29054.4]
  assign x295_1_io_flow = io_in_x185_TREADY; // @[Math.scala 265:20:@29055.4]
  assign x296_1_clock = clock; // @[:@29063.4]
  assign x296_1_io_a = x217_lb_0_io_rPort_7_output_0; // @[Math.scala 263:17:@29065.4]
  assign x296_1_io_b = 32'h2; // @[Math.scala 264:17:@29066.4]
  assign x296_1_io_flow = io_in_x185_TREADY; // @[Math.scala 265:20:@29067.4]
  assign x297_1_clock = clock; // @[:@29075.4]
  assign x297_1_io_a = x217_lb_0_io_rPort_3_output_0; // @[Math.scala 263:17:@29077.4]
  assign x297_1_io_b = 32'h1; // @[Math.scala 264:17:@29078.4]
  assign x297_1_io_flow = io_in_x185_TREADY; // @[Math.scala 265:20:@29079.4]
  assign x298_1_clock = clock; // @[:@29087.4]
  assign x298_1_io_a = x217_lb_0_io_rPort_6_output_0; // @[Math.scala 263:17:@29089.4]
  assign x298_1_io_b = 32'h2; // @[Math.scala 264:17:@29090.4]
  assign x298_1_io_flow = io_in_x185_TREADY; // @[Math.scala 265:20:@29091.4]
  assign x299_1_clock = clock; // @[:@29099.4]
  assign x299_1_io_a = x217_lb_0_io_rPort_4_output_0; // @[Math.scala 263:17:@29101.4]
  assign x299_1_io_b = 32'h4; // @[Math.scala 264:17:@29102.4]
  assign x299_1_io_flow = io_in_x185_TREADY; // @[Math.scala 265:20:@29103.4]
  assign x300_1_clock = clock; // @[:@29113.4]
  assign x300_1_io_a = x217_lb_0_io_rPort_5_output_0; // @[Math.scala 263:17:@29115.4]
  assign x300_1_io_b = 32'h2; // @[Math.scala 264:17:@29116.4]
  assign x300_1_io_flow = io_in_x185_TREADY; // @[Math.scala 265:20:@29117.4]
  assign x301_1_clock = clock; // @[:@29125.4]
  assign x301_1_io_a = x217_lb_0_io_rPort_8_output_0; // @[Math.scala 263:17:@29127.4]
  assign x301_1_io_b = 32'h1; // @[Math.scala 264:17:@29128.4]
  assign x301_1_io_flow = io_in_x185_TREADY; // @[Math.scala 265:20:@29129.4]
  assign x302_1_clock = clock; // @[:@29137.4]
  assign x302_1_io_a = x217_lb_0_io_rPort_0_output_0; // @[Math.scala 263:17:@29139.4]
  assign x302_1_io_b = 32'h2; // @[Math.scala 264:17:@29140.4]
  assign x302_1_io_flow = io_in_x185_TREADY; // @[Math.scala 265:20:@29141.4]
  assign x303_1_clock = clock; // @[:@29149.4]
  assign x303_1_io_a = x217_lb_0_io_rPort_1_output_0; // @[Math.scala 263:17:@29151.4]
  assign x303_1_io_b = 32'h1; // @[Math.scala 264:17:@29152.4]
  assign x303_1_io_flow = io_in_x185_TREADY; // @[Math.scala 265:20:@29153.4]
  assign x304_x3_1_clock = clock; // @[:@29159.4]
  assign x304_x3_1_reset = reset; // @[:@29160.4]
  assign x304_x3_1_io_a = x295_1_io_result; // @[Math.scala 151:17:@29161.4]
  assign x304_x3_1_io_b = x296_1_io_result; // @[Math.scala 152:17:@29162.4]
  assign x304_x3_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@29163.4]
  assign x305_x4_1_clock = clock; // @[:@29169.4]
  assign x305_x4_1_reset = reset; // @[:@29170.4]
  assign x305_x4_1_io_a = x297_1_io_result; // @[Math.scala 151:17:@29171.4]
  assign x305_x4_1_io_b = x298_1_io_result; // @[Math.scala 152:17:@29172.4]
  assign x305_x4_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@29173.4]
  assign x306_x3_1_clock = clock; // @[:@29179.4]
  assign x306_x3_1_reset = reset; // @[:@29180.4]
  assign x306_x3_1_io_a = x299_1_io_result; // @[Math.scala 151:17:@29181.4]
  assign x306_x3_1_io_b = x300_1_io_result; // @[Math.scala 152:17:@29182.4]
  assign x306_x3_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@29183.4]
  assign x307_x4_1_clock = clock; // @[:@29189.4]
  assign x307_x4_1_reset = reset; // @[:@29190.4]
  assign x307_x4_1_io_a = x301_1_io_result; // @[Math.scala 151:17:@29191.4]
  assign x307_x4_1_io_b = x302_1_io_result; // @[Math.scala 152:17:@29192.4]
  assign x307_x4_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@29193.4]
  assign x308_x3_1_clock = clock; // @[:@29199.4]
  assign x308_x3_1_reset = reset; // @[:@29200.4]
  assign x308_x3_1_io_a = x304_x3_1_io_result; // @[Math.scala 151:17:@29201.4]
  assign x308_x3_1_io_b = x305_x4_1_io_result; // @[Math.scala 152:17:@29202.4]
  assign x308_x3_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@29203.4]
  assign x309_x4_1_clock = clock; // @[:@29209.4]
  assign x309_x4_1_reset = reset; // @[:@29210.4]
  assign x309_x4_1_io_a = x306_x3_1_io_result; // @[Math.scala 151:17:@29211.4]
  assign x309_x4_1_io_b = x307_x4_1_io_result; // @[Math.scala 152:17:@29212.4]
  assign x309_x4_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@29213.4]
  assign x310_x3_1_clock = clock; // @[:@29219.4]
  assign x310_x3_1_reset = reset; // @[:@29220.4]
  assign x310_x3_1_io_a = x308_x3_1_io_result; // @[Math.scala 151:17:@29221.4]
  assign x310_x3_1_io_b = x309_x4_1_io_result; // @[Math.scala 152:17:@29222.4]
  assign x310_x3_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@29223.4]
  assign RetimeWrapper_72_clock = clock; // @[:@29229.4]
  assign RetimeWrapper_72_reset = reset; // @[:@29230.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29232.4]
  assign RetimeWrapper_72_io_in = x303_1_io_result; // @[package.scala 94:16:@29231.4]
  assign x311_sum_1_clock = clock; // @[:@29238.4]
  assign x311_sum_1_reset = reset; // @[:@29239.4]
  assign x311_sum_1_io_a = x310_x3_1_io_result; // @[Math.scala 151:17:@29240.4]
  assign x311_sum_1_io_b = RetimeWrapper_72_io_out; // @[Math.scala 152:17:@29241.4]
  assign x311_sum_1_io_flow = io_in_x185_TREADY; // @[Math.scala 153:20:@29242.4]
  assign x312_1_io_b = x311_sum_1_io_result; // @[Math.scala 721:17:@29250.4]
  assign x313_mul_1_clock = clock; // @[:@29259.4]
  assign x313_mul_1_io_a = x312_1_io_result; // @[Math.scala 263:17:@29261.4]
  assign x313_mul_1_io_flow = io_in_x185_TREADY; // @[Math.scala 265:20:@29263.4]
  assign x314_1_io_b = x313_mul_1_io_result; // @[Math.scala 721:17:@29271.4]
  assign RetimeWrapper_73_clock = clock; // @[:@29282.4]
  assign RetimeWrapper_73_reset = reset; // @[:@29283.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29285.4]
  assign RetimeWrapper_73_io_in = x314_1_io_result; // @[package.scala 94:16:@29284.4]
  assign RetimeWrapper_74_clock = clock; // @[:@29291.4]
  assign RetimeWrapper_74_reset = reset; // @[:@29292.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29294.4]
  assign RetimeWrapper_74_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@29293.4]
  assign RetimeWrapper_75_clock = clock; // @[:@29300.4]
  assign RetimeWrapper_75_reset = reset; // @[:@29301.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29303.4]
  assign RetimeWrapper_75_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@29302.4]
  assign RetimeWrapper_76_clock = clock; // @[:@29309.4]
  assign RetimeWrapper_76_reset = reset; // @[:@29310.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29312.4]
  assign RetimeWrapper_76_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@29311.4]
endmodule
module x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1( // @[:@29330.2]
  input          clock, // @[:@29331.4]
  input          reset, // @[:@29332.4]
  output         io_in_x185_TVALID, // @[:@29333.4]
  input          io_in_x185_TREADY, // @[:@29333.4]
  output [255:0] io_in_x185_TDATA, // @[:@29333.4]
  input          io_in_x184_TVALID, // @[:@29333.4]
  output         io_in_x184_TREADY, // @[:@29333.4]
  input  [255:0] io_in_x184_TDATA, // @[:@29333.4]
  input  [7:0]   io_in_x184_TID, // @[:@29333.4]
  input  [7:0]   io_in_x184_TDEST, // @[:@29333.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@29333.4]
  input          io_sigsIn_smChildAcks_0, // @[:@29333.4]
  output         io_sigsOut_smDoneIn_0, // @[:@29333.4]
  input          io_rr // @[:@29333.4]
);
  wire  x210_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@29367.4]
  wire  x210_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@29367.4]
  wire  x210_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@29367.4]
  wire  x210_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@29367.4]
  wire [12:0] x210_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@29367.4]
  wire [12:0] x210_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@29367.4]
  wire  x210_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@29367.4]
  wire  x210_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@29367.4]
  wire  x210_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@29367.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 32:18:@29427.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 32:18:@29427.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 32:18:@29427.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 32:18:@29427.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 32:18:@29427.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 32:18:@29427.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 32:18:@29427.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 32:18:@29427.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 32:18:@29427.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 32:18:@29427.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 32:18:@29427.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 32:18:@29427.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@29455.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@29455.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@29455.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@29455.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@29455.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@29497.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@29497.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@29497.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@29497.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@29497.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@29505.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@29505.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@29505.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@29505.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@29505.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 576:24:@29539.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 576:24:@29539.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x185_TVALID; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 576:24:@29539.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x185_TREADY; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 576:24:@29539.4]
  wire [255:0] x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x185_TDATA; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 576:24:@29539.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x184_TREADY; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 576:24:@29539.4]
  wire [255:0] x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x184_TDATA; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 576:24:@29539.4]
  wire [7:0] x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x184_TID; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 576:24:@29539.4]
  wire [7:0] x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x184_TDEST; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 576:24:@29539.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 576:24:@29539.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 576:24:@29539.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 576:24:@29539.4]
  wire [31:0] x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 576:24:@29539.4]
  wire [31:0] x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 576:24:@29539.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 576:24:@29539.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 576:24:@29539.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 576:24:@29539.4]
  wire  _T_240; // @[package.scala 96:25:@29460.4 package.scala 96:25:@29461.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x320_outr_UnitPipe.scala 69:66:@29466.4]
  wire  _T_253; // @[package.scala 96:25:@29502.4 package.scala 96:25:@29503.4]
  wire  _T_259; // @[package.scala 96:25:@29510.4 package.scala 96:25:@29511.4]
  wire  _T_262; // @[SpatialBlocks.scala 138:93:@29513.4]
  wire  x319_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@29514.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:36:@29522.4]
  wire  _T_265; // @[SpatialBlocks.scala 157:78:@29523.4]
  wire  _T_272; // @[SpatialBlocks.scala 159:58:@29535.4]
  x192_ctrchain x210_ctrchain ( // @[SpatialBlocks.scala 37:22:@29367.4]
    .clock(x210_ctrchain_clock),
    .reset(x210_ctrchain_reset),
    .io_input_reset(x210_ctrchain_io_input_reset),
    .io_input_enable(x210_ctrchain_io_input_enable),
    .io_output_counts_1(x210_ctrchain_io_output_counts_1),
    .io_output_counts_0(x210_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x210_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x210_ctrchain_io_output_oobs_1),
    .io_output_done(x210_ctrchain_io_output_done)
  );
  x319_inr_Foreach_SAMPLER_BOX_sm x319_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 32:18:@29427.4]
    .clock(x319_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x319_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x319_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x319_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x319_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x319_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x319_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x319_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x319_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x319_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x319_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x319_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@29455.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@29497.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@29505.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1 x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 576:24:@29539.4]
    .clock(x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x185_TVALID(x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x185_TVALID),
    .io_in_x185_TREADY(x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x185_TREADY),
    .io_in_x185_TDATA(x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x185_TDATA),
    .io_in_x184_TREADY(x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x184_TREADY),
    .io_in_x184_TDATA(x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x184_TDATA),
    .io_in_x184_TID(x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x184_TID),
    .io_in_x184_TDEST(x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x184_TDEST),
    .io_sigsIn_backpressure(x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_240 = RetimeWrapper_io_out; // @[package.scala 96:25:@29460.4 package.scala 96:25:@29461.4]
  assign x319_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x184_TVALID | x319_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x320_outr_UnitPipe.scala 69:66:@29466.4]
  assign _T_253 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@29502.4 package.scala 96:25:@29503.4]
  assign _T_259 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@29510.4 package.scala 96:25:@29511.4]
  assign _T_262 = ~ _T_259; // @[SpatialBlocks.scala 138:93:@29513.4]
  assign x319_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_253 & _T_262; // @[SpatialBlocks.scala 138:90:@29514.4]
  assign _T_264 = x319_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@29522.4]
  assign _T_265 = ~ x319_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@29523.4]
  assign _T_272 = x319_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@29535.4]
  assign io_in_x185_TVALID = x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x185_TVALID; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 48:23:@29598.4]
  assign io_in_x185_TDATA = x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x185_TDATA; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 48:23:@29596.4]
  assign io_in_x184_TREADY = x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x184_TREADY; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 49:23:@29606.4]
  assign io_sigsOut_smDoneIn_0 = x319_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@29520.4]
  assign x210_ctrchain_clock = clock; // @[:@29368.4]
  assign x210_ctrchain_reset = reset; // @[:@29369.4]
  assign x210_ctrchain_io_input_reset = x319_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@29538.4]
  assign x210_ctrchain_io_input_enable = _T_272 & x319_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@29490.4 SpatialBlocks.scala 159:42:@29537.4]
  assign x319_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@29428.4]
  assign x319_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@29429.4]
  assign x319_inr_Foreach_SAMPLER_BOX_sm_io_enable = x319_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x319_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@29517.4]
  assign x319_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_240 : 1'h0; // @[sm_x320_outr_UnitPipe.scala 67:50:@29463.4]
  assign x319_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@29519.4]
  assign x319_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x185_TREADY | x319_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@29491.4]
  assign x319_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x320_outr_UnitPipe.scala 71:48:@29469.4]
  assign RetimeWrapper_clock = clock; // @[:@29456.4]
  assign RetimeWrapper_reset = reset; // @[:@29457.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@29459.4]
  assign RetimeWrapper_io_in = x210_ctrchain_io_output_done; // @[package.scala 94:16:@29458.4]
  assign RetimeWrapper_1_clock = clock; // @[:@29498.4]
  assign RetimeWrapper_1_reset = reset; // @[:@29499.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@29501.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@29500.4]
  assign RetimeWrapper_2_clock = clock; // @[:@29506.4]
  assign RetimeWrapper_2_reset = reset; // @[:@29507.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@29509.4]
  assign RetimeWrapper_2_io_in = x319_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@29508.4]
  assign x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@29540.4]
  assign x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@29541.4]
  assign x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x185_TREADY = io_in_x185_TREADY; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 48:23:@29597.4]
  assign x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x184_TDATA = io_in_x184_TDATA; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 49:23:@29605.4]
  assign x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x184_TID = io_in_x184_TID; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 49:23:@29601.4]
  assign x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x184_TDEST = io_in_x184_TDEST; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 49:23:@29600.4]
  assign x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x185_TREADY | x319_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 581:22:@29624.4]
  assign x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_264 & _T_265; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 581:22:@29622.4]
  assign x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x319_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 581:22:@29620.4]
  assign x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x210_ctrchain_io_output_counts_1[12]}},x210_ctrchain_io_output_counts_1}; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 581:22:@29615.4]
  assign x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x210_ctrchain_io_output_counts_0[12]}},x210_ctrchain_io_output_counts_0}; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 581:22:@29614.4]
  assign x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x210_ctrchain_io_output_oobs_0; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 581:22:@29612.4]
  assign x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x210_ctrchain_io_output_oobs_1; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 581:22:@29613.4]
  assign x319_inr_Foreach_SAMPLER_BOX_kernelx319_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x319_inr_Foreach_SAMPLER_BOX.scala 580:18:@29608.4]
endmodule
module x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1( // @[:@29638.2]
  input          clock, // @[:@29639.4]
  input          reset, // @[:@29640.4]
  output         io_in_x185_TVALID, // @[:@29641.4]
  input          io_in_x185_TREADY, // @[:@29641.4]
  output [255:0] io_in_x185_TDATA, // @[:@29641.4]
  input          io_in_x184_TVALID, // @[:@29641.4]
  output         io_in_x184_TREADY, // @[:@29641.4]
  input  [255:0] io_in_x184_TDATA, // @[:@29641.4]
  input  [7:0]   io_in_x184_TID, // @[:@29641.4]
  input  [7:0]   io_in_x184_TDEST, // @[:@29641.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@29641.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@29641.4]
  input          io_sigsIn_smChildAcks_0, // @[:@29641.4]
  input          io_sigsIn_smChildAcks_1, // @[:@29641.4]
  output         io_sigsOut_smDoneIn_0, // @[:@29641.4]
  output         io_sigsOut_smDoneIn_1, // @[:@29641.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@29641.4]
  output         io_sigsOut_smCtrCopyDone_1, // @[:@29641.4]
  input          io_rr // @[:@29641.4]
);
  wire  x187_fifoinraw_0_clock; // @[m_x187_fifoinraw_0.scala 27:17:@29655.4]
  wire  x187_fifoinraw_0_reset; // @[m_x187_fifoinraw_0.scala 27:17:@29655.4]
  wire  x188_fifoinpacked_0_clock; // @[m_x188_fifoinpacked_0.scala 27:17:@29679.4]
  wire  x188_fifoinpacked_0_reset; // @[m_x188_fifoinpacked_0.scala 27:17:@29679.4]
  wire  x188_fifoinpacked_0_io_wPort_0_en_0; // @[m_x188_fifoinpacked_0.scala 27:17:@29679.4]
  wire  x188_fifoinpacked_0_io_full; // @[m_x188_fifoinpacked_0.scala 27:17:@29679.4]
  wire  x188_fifoinpacked_0_io_active_0_in; // @[m_x188_fifoinpacked_0.scala 27:17:@29679.4]
  wire  x188_fifoinpacked_0_io_active_0_out; // @[m_x188_fifoinpacked_0.scala 27:17:@29679.4]
  wire  x189_fifooutraw_0_clock; // @[m_x189_fifooutraw_0.scala 27:17:@29703.4]
  wire  x189_fifooutraw_0_reset; // @[m_x189_fifooutraw_0.scala 27:17:@29703.4]
  wire  x192_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@29727.4]
  wire  x192_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@29727.4]
  wire  x192_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@29727.4]
  wire  x192_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@29727.4]
  wire [12:0] x192_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@29727.4]
  wire [12:0] x192_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@29727.4]
  wire  x192_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@29727.4]
  wire  x192_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@29727.4]
  wire  x192_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@29727.4]
  wire  x206_inr_Foreach_sm_clock; // @[sm_x206_inr_Foreach.scala 32:18:@29787.4]
  wire  x206_inr_Foreach_sm_reset; // @[sm_x206_inr_Foreach.scala 32:18:@29787.4]
  wire  x206_inr_Foreach_sm_io_enable; // @[sm_x206_inr_Foreach.scala 32:18:@29787.4]
  wire  x206_inr_Foreach_sm_io_done; // @[sm_x206_inr_Foreach.scala 32:18:@29787.4]
  wire  x206_inr_Foreach_sm_io_doneLatch; // @[sm_x206_inr_Foreach.scala 32:18:@29787.4]
  wire  x206_inr_Foreach_sm_io_ctrDone; // @[sm_x206_inr_Foreach.scala 32:18:@29787.4]
  wire  x206_inr_Foreach_sm_io_datapathEn; // @[sm_x206_inr_Foreach.scala 32:18:@29787.4]
  wire  x206_inr_Foreach_sm_io_ctrInc; // @[sm_x206_inr_Foreach.scala 32:18:@29787.4]
  wire  x206_inr_Foreach_sm_io_ctrRst; // @[sm_x206_inr_Foreach.scala 32:18:@29787.4]
  wire  x206_inr_Foreach_sm_io_parentAck; // @[sm_x206_inr_Foreach.scala 32:18:@29787.4]
  wire  x206_inr_Foreach_sm_io_backpressure; // @[sm_x206_inr_Foreach.scala 32:18:@29787.4]
  wire  x206_inr_Foreach_sm_io_break; // @[sm_x206_inr_Foreach.scala 32:18:@29787.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@29815.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@29815.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@29815.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@29815.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@29815.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@29861.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@29861.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@29861.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@29861.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@29861.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@29869.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@29869.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@29869.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@29869.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@29869.4]
  wire  x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_clock; // @[sm_x206_inr_Foreach.scala 96:24:@29904.4]
  wire  x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_reset; // @[sm_x206_inr_Foreach.scala 96:24:@29904.4]
  wire  x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_in_x188_fifoinpacked_0_wPort_0_en_0; // @[sm_x206_inr_Foreach.scala 96:24:@29904.4]
  wire  x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_in_x188_fifoinpacked_0_full; // @[sm_x206_inr_Foreach.scala 96:24:@29904.4]
  wire  x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_in_x188_fifoinpacked_0_active_0_in; // @[sm_x206_inr_Foreach.scala 96:24:@29904.4]
  wire  x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_in_x188_fifoinpacked_0_active_0_out; // @[sm_x206_inr_Foreach.scala 96:24:@29904.4]
  wire  x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x206_inr_Foreach.scala 96:24:@29904.4]
  wire  x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x206_inr_Foreach.scala 96:24:@29904.4]
  wire  x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x206_inr_Foreach.scala 96:24:@29904.4]
  wire [31:0] x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x206_inr_Foreach.scala 96:24:@29904.4]
  wire [31:0] x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x206_inr_Foreach.scala 96:24:@29904.4]
  wire  x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x206_inr_Foreach.scala 96:24:@29904.4]
  wire  x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x206_inr_Foreach.scala 96:24:@29904.4]
  wire  x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_rr; // @[sm_x206_inr_Foreach.scala 96:24:@29904.4]
  wire  x320_outr_UnitPipe_sm_clock; // @[sm_x320_outr_UnitPipe.scala 32:18:@30036.4]
  wire  x320_outr_UnitPipe_sm_reset; // @[sm_x320_outr_UnitPipe.scala 32:18:@30036.4]
  wire  x320_outr_UnitPipe_sm_io_enable; // @[sm_x320_outr_UnitPipe.scala 32:18:@30036.4]
  wire  x320_outr_UnitPipe_sm_io_done; // @[sm_x320_outr_UnitPipe.scala 32:18:@30036.4]
  wire  x320_outr_UnitPipe_sm_io_rst; // @[sm_x320_outr_UnitPipe.scala 32:18:@30036.4]
  wire  x320_outr_UnitPipe_sm_io_ctrDone; // @[sm_x320_outr_UnitPipe.scala 32:18:@30036.4]
  wire  x320_outr_UnitPipe_sm_io_ctrInc; // @[sm_x320_outr_UnitPipe.scala 32:18:@30036.4]
  wire  x320_outr_UnitPipe_sm_io_parentAck; // @[sm_x320_outr_UnitPipe.scala 32:18:@30036.4]
  wire  x320_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x320_outr_UnitPipe.scala 32:18:@30036.4]
  wire  x320_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x320_outr_UnitPipe.scala 32:18:@30036.4]
  wire  x320_outr_UnitPipe_sm_io_childAck_0; // @[sm_x320_outr_UnitPipe.scala 32:18:@30036.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@30093.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@30093.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@30093.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@30093.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@30093.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@30101.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@30101.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@30101.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@30101.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@30101.4]
  wire  x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_clock; // @[sm_x320_outr_UnitPipe.scala 76:24:@30131.4]
  wire  x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_reset; // @[sm_x320_outr_UnitPipe.scala 76:24:@30131.4]
  wire  x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x185_TVALID; // @[sm_x320_outr_UnitPipe.scala 76:24:@30131.4]
  wire  x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x185_TREADY; // @[sm_x320_outr_UnitPipe.scala 76:24:@30131.4]
  wire [255:0] x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x185_TDATA; // @[sm_x320_outr_UnitPipe.scala 76:24:@30131.4]
  wire  x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x184_TVALID; // @[sm_x320_outr_UnitPipe.scala 76:24:@30131.4]
  wire  x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x184_TREADY; // @[sm_x320_outr_UnitPipe.scala 76:24:@30131.4]
  wire [255:0] x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x184_TDATA; // @[sm_x320_outr_UnitPipe.scala 76:24:@30131.4]
  wire [7:0] x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x184_TID; // @[sm_x320_outr_UnitPipe.scala 76:24:@30131.4]
  wire [7:0] x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x184_TDEST; // @[sm_x320_outr_UnitPipe.scala 76:24:@30131.4]
  wire  x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x320_outr_UnitPipe.scala 76:24:@30131.4]
  wire  x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x320_outr_UnitPipe.scala 76:24:@30131.4]
  wire  x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x320_outr_UnitPipe.scala 76:24:@30131.4]
  wire  x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_rr; // @[sm_x320_outr_UnitPipe.scala 76:24:@30131.4]
  wire  _T_254; // @[package.scala 96:25:@29820.4 package.scala 96:25:@29821.4]
  wire  _T_260; // @[implicits.scala 47:10:@29824.4]
  wire  _T_261; // @[sm_x321_outr_UnitPipe.scala 70:41:@29825.4]
  wire  _T_262; // @[sm_x321_outr_UnitPipe.scala 70:78:@29826.4]
  wire  _T_263; // @[sm_x321_outr_UnitPipe.scala 70:76:@29827.4]
  wire  _T_275; // @[package.scala 96:25:@29866.4 package.scala 96:25:@29867.4]
  wire  _T_281; // @[package.scala 96:25:@29874.4 package.scala 96:25:@29875.4]
  wire  _T_284; // @[SpatialBlocks.scala 138:93:@29877.4]
  wire  _T_286; // @[SpatialBlocks.scala 157:36:@29886.4]
  wire  _T_287; // @[SpatialBlocks.scala 157:78:@29887.4]
  wire  _T_354; // @[package.scala 100:49:@30064.4]
  reg  _T_357; // @[package.scala 48:56:@30065.4]
  reg [31:0] _RAND_0;
  wire  _T_371; // @[package.scala 96:25:@30098.4 package.scala 96:25:@30099.4]
  wire  _T_377; // @[package.scala 96:25:@30106.4 package.scala 96:25:@30107.4]
  wire  _T_380; // @[SpatialBlocks.scala 138:93:@30109.4]
  x187_fifoinraw_0 x187_fifoinraw_0 ( // @[m_x187_fifoinraw_0.scala 27:17:@29655.4]
    .clock(x187_fifoinraw_0_clock),
    .reset(x187_fifoinraw_0_reset)
  );
  x188_fifoinpacked_0 x188_fifoinpacked_0 ( // @[m_x188_fifoinpacked_0.scala 27:17:@29679.4]
    .clock(x188_fifoinpacked_0_clock),
    .reset(x188_fifoinpacked_0_reset),
    .io_wPort_0_en_0(x188_fifoinpacked_0_io_wPort_0_en_0),
    .io_full(x188_fifoinpacked_0_io_full),
    .io_active_0_in(x188_fifoinpacked_0_io_active_0_in),
    .io_active_0_out(x188_fifoinpacked_0_io_active_0_out)
  );
  x187_fifoinraw_0 x189_fifooutraw_0 ( // @[m_x189_fifooutraw_0.scala 27:17:@29703.4]
    .clock(x189_fifooutraw_0_clock),
    .reset(x189_fifooutraw_0_reset)
  );
  x192_ctrchain x192_ctrchain ( // @[SpatialBlocks.scala 37:22:@29727.4]
    .clock(x192_ctrchain_clock),
    .reset(x192_ctrchain_reset),
    .io_input_reset(x192_ctrchain_io_input_reset),
    .io_input_enable(x192_ctrchain_io_input_enable),
    .io_output_counts_1(x192_ctrchain_io_output_counts_1),
    .io_output_counts_0(x192_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x192_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x192_ctrchain_io_output_oobs_1),
    .io_output_done(x192_ctrchain_io_output_done)
  );
  x206_inr_Foreach_sm x206_inr_Foreach_sm ( // @[sm_x206_inr_Foreach.scala 32:18:@29787.4]
    .clock(x206_inr_Foreach_sm_clock),
    .reset(x206_inr_Foreach_sm_reset),
    .io_enable(x206_inr_Foreach_sm_io_enable),
    .io_done(x206_inr_Foreach_sm_io_done),
    .io_doneLatch(x206_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x206_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x206_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x206_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x206_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x206_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x206_inr_Foreach_sm_io_backpressure),
    .io_break(x206_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@29815.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@29861.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@29869.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x206_inr_Foreach_kernelx206_inr_Foreach_concrete1 x206_inr_Foreach_kernelx206_inr_Foreach_concrete1 ( // @[sm_x206_inr_Foreach.scala 96:24:@29904.4]
    .clock(x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_clock),
    .reset(x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_reset),
    .io_in_x188_fifoinpacked_0_wPort_0_en_0(x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_in_x188_fifoinpacked_0_wPort_0_en_0),
    .io_in_x188_fifoinpacked_0_full(x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_in_x188_fifoinpacked_0_full),
    .io_in_x188_fifoinpacked_0_active_0_in(x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_in_x188_fifoinpacked_0_active_0_in),
    .io_in_x188_fifoinpacked_0_active_0_out(x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_in_x188_fifoinpacked_0_active_0_out),
    .io_sigsIn_backpressure(x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_rr)
  );
  RootController_sm x320_outr_UnitPipe_sm ( // @[sm_x320_outr_UnitPipe.scala 32:18:@30036.4]
    .clock(x320_outr_UnitPipe_sm_clock),
    .reset(x320_outr_UnitPipe_sm_reset),
    .io_enable(x320_outr_UnitPipe_sm_io_enable),
    .io_done(x320_outr_UnitPipe_sm_io_done),
    .io_rst(x320_outr_UnitPipe_sm_io_rst),
    .io_ctrDone(x320_outr_UnitPipe_sm_io_ctrDone),
    .io_ctrInc(x320_outr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x320_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x320_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x320_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x320_outr_UnitPipe_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@30093.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@30101.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1 x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1 ( // @[sm_x320_outr_UnitPipe.scala 76:24:@30131.4]
    .clock(x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_clock),
    .reset(x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_reset),
    .io_in_x185_TVALID(x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x185_TVALID),
    .io_in_x185_TREADY(x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x185_TREADY),
    .io_in_x185_TDATA(x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x185_TDATA),
    .io_in_x184_TVALID(x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x184_TVALID),
    .io_in_x184_TREADY(x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x184_TREADY),
    .io_in_x184_TDATA(x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x184_TDATA),
    .io_in_x184_TID(x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x184_TID),
    .io_in_x184_TDEST(x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x184_TDEST),
    .io_sigsIn_smEnableOuts_0(x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_254 = RetimeWrapper_io_out; // @[package.scala 96:25:@29820.4 package.scala 96:25:@29821.4]
  assign _T_260 = x188_fifoinpacked_0_io_full; // @[implicits.scala 47:10:@29824.4]
  assign _T_261 = ~ _T_260; // @[sm_x321_outr_UnitPipe.scala 70:41:@29825.4]
  assign _T_262 = ~ x188_fifoinpacked_0_io_active_0_out; // @[sm_x321_outr_UnitPipe.scala 70:78:@29826.4]
  assign _T_263 = _T_261 | _T_262; // @[sm_x321_outr_UnitPipe.scala 70:76:@29827.4]
  assign _T_275 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@29866.4 package.scala 96:25:@29867.4]
  assign _T_281 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@29874.4 package.scala 96:25:@29875.4]
  assign _T_284 = ~ _T_281; // @[SpatialBlocks.scala 138:93:@29877.4]
  assign _T_286 = x206_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@29886.4]
  assign _T_287 = ~ x206_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@29887.4]
  assign _T_354 = x320_outr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@30064.4]
  assign _T_371 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@30098.4 package.scala 96:25:@30099.4]
  assign _T_377 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@30106.4 package.scala 96:25:@30107.4]
  assign _T_380 = ~ _T_377; // @[SpatialBlocks.scala 138:93:@30109.4]
  assign io_in_x185_TVALID = x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x185_TVALID; // @[sm_x320_outr_UnitPipe.scala 48:23:@30188.4]
  assign io_in_x185_TDATA = x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x185_TDATA; // @[sm_x320_outr_UnitPipe.scala 48:23:@30186.4]
  assign io_in_x184_TREADY = x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x184_TREADY; // @[sm_x320_outr_UnitPipe.scala 49:23:@30196.4]
  assign io_sigsOut_smDoneIn_0 = x206_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@29884.4]
  assign io_sigsOut_smDoneIn_1 = x320_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@30116.4]
  assign io_sigsOut_smCtrCopyDone_0 = x206_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@29903.4]
  assign io_sigsOut_smCtrCopyDone_1 = x320_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@30130.4]
  assign x187_fifoinraw_0_clock = clock; // @[:@29656.4]
  assign x187_fifoinraw_0_reset = reset; // @[:@29657.4]
  assign x188_fifoinpacked_0_clock = clock; // @[:@29680.4]
  assign x188_fifoinpacked_0_reset = reset; // @[:@29681.4]
  assign x188_fifoinpacked_0_io_wPort_0_en_0 = x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_in_x188_fifoinpacked_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@29964.4]
  assign x188_fifoinpacked_0_io_active_0_in = x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_in_x188_fifoinpacked_0_active_0_in; // @[MemInterfaceType.scala 167:86:@29963.4]
  assign x189_fifooutraw_0_clock = clock; // @[:@29704.4]
  assign x189_fifooutraw_0_reset = reset; // @[:@29705.4]
  assign x192_ctrchain_clock = clock; // @[:@29728.4]
  assign x192_ctrchain_reset = reset; // @[:@29729.4]
  assign x192_ctrchain_io_input_reset = x206_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@29902.4]
  assign x192_ctrchain_io_input_enable = x206_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@29854.4 SpatialBlocks.scala 159:42:@29901.4]
  assign x206_inr_Foreach_sm_clock = clock; // @[:@29788.4]
  assign x206_inr_Foreach_sm_reset = reset; // @[:@29789.4]
  assign x206_inr_Foreach_sm_io_enable = _T_275 & _T_284; // @[SpatialBlocks.scala 140:18:@29881.4]
  assign x206_inr_Foreach_sm_io_ctrDone = io_rr ? _T_254 : 1'h0; // @[sm_x321_outr_UnitPipe.scala 69:38:@29823.4]
  assign x206_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@29883.4]
  assign x206_inr_Foreach_sm_io_backpressure = _T_263 | x206_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@29855.4]
  assign x206_inr_Foreach_sm_io_break = 1'h0; // @[sm_x321_outr_UnitPipe.scala 73:36:@29833.4]
  assign RetimeWrapper_clock = clock; // @[:@29816.4]
  assign RetimeWrapper_reset = reset; // @[:@29817.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@29819.4]
  assign RetimeWrapper_io_in = x192_ctrchain_io_output_done; // @[package.scala 94:16:@29818.4]
  assign RetimeWrapper_1_clock = clock; // @[:@29862.4]
  assign RetimeWrapper_1_reset = reset; // @[:@29863.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@29865.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@29864.4]
  assign RetimeWrapper_2_clock = clock; // @[:@29870.4]
  assign RetimeWrapper_2_reset = reset; // @[:@29871.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@29873.4]
  assign RetimeWrapper_2_io_in = x206_inr_Foreach_sm_io_done; // @[package.scala 94:16:@29872.4]
  assign x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_clock = clock; // @[:@29905.4]
  assign x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_reset = reset; // @[:@29906.4]
  assign x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_in_x188_fifoinpacked_0_full = x188_fifoinpacked_0_io_full; // @[MemInterfaceType.scala 159:15:@29958.4]
  assign x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_in_x188_fifoinpacked_0_active_0_out = x188_fifoinpacked_0_io_active_0_out; // @[MemInterfaceType.scala 158:75:@29957.4]
  assign x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_263 | x206_inr_Foreach_sm_io_doneLatch; // @[sm_x206_inr_Foreach.scala 101:22:@29987.4]
  assign x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_286 & _T_287; // @[sm_x206_inr_Foreach.scala 101:22:@29985.4]
  assign x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_break = x206_inr_Foreach_sm_io_break; // @[sm_x206_inr_Foreach.scala 101:22:@29983.4]
  assign x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x192_ctrchain_io_output_counts_1[12]}},x192_ctrchain_io_output_counts_1}; // @[sm_x206_inr_Foreach.scala 101:22:@29978.4]
  assign x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x192_ctrchain_io_output_counts_0[12]}},x192_ctrchain_io_output_counts_0}; // @[sm_x206_inr_Foreach.scala 101:22:@29977.4]
  assign x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x192_ctrchain_io_output_oobs_0; // @[sm_x206_inr_Foreach.scala 101:22:@29975.4]
  assign x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x192_ctrchain_io_output_oobs_1; // @[sm_x206_inr_Foreach.scala 101:22:@29976.4]
  assign x206_inr_Foreach_kernelx206_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x206_inr_Foreach.scala 100:18:@29971.4]
  assign x320_outr_UnitPipe_sm_clock = clock; // @[:@30037.4]
  assign x320_outr_UnitPipe_sm_reset = reset; // @[:@30038.4]
  assign x320_outr_UnitPipe_sm_io_enable = _T_371 & _T_380; // @[SpatialBlocks.scala 140:18:@30113.4]
  assign x320_outr_UnitPipe_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 134:15:@30088.4]
  assign x320_outr_UnitPipe_sm_io_ctrDone = x320_outr_UnitPipe_sm_io_ctrInc & _T_357; // @[sm_x321_outr_UnitPipe.scala 78:40:@30068.4]
  assign x320_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@30115.4]
  assign x320_outr_UnitPipe_sm_io_doneIn_0 = x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@30085.4]
  assign RetimeWrapper_3_clock = clock; // @[:@30094.4]
  assign RetimeWrapper_3_reset = reset; // @[:@30095.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@30097.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@30096.4]
  assign RetimeWrapper_4_clock = clock; // @[:@30102.4]
  assign RetimeWrapper_4_reset = reset; // @[:@30103.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@30105.4]
  assign RetimeWrapper_4_io_in = x320_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@30104.4]
  assign x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_clock = clock; // @[:@30132.4]
  assign x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_reset = reset; // @[:@30133.4]
  assign x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x185_TREADY = io_in_x185_TREADY; // @[sm_x320_outr_UnitPipe.scala 48:23:@30187.4]
  assign x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x184_TVALID = io_in_x184_TVALID; // @[sm_x320_outr_UnitPipe.scala 49:23:@30197.4]
  assign x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x184_TDATA = io_in_x184_TDATA; // @[sm_x320_outr_UnitPipe.scala 49:23:@30195.4]
  assign x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x184_TID = io_in_x184_TID; // @[sm_x320_outr_UnitPipe.scala 49:23:@30191.4]
  assign x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_in_x184_TDEST = io_in_x184_TDEST; // @[sm_x320_outr_UnitPipe.scala 49:23:@30190.4]
  assign x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x320_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x320_outr_UnitPipe.scala 81:22:@30206.4]
  assign x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x320_outr_UnitPipe_sm_io_childAck_0; // @[sm_x320_outr_UnitPipe.scala 81:22:@30204.4]
  assign x320_outr_UnitPipe_kernelx320_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x320_outr_UnitPipe.scala 80:18:@30198.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_357 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_357 <= 1'h0;
    end else begin
      _T_357 <= _T_354;
    end
  end
endmodule
module x343_outr_UnitPipe_sm( // @[:@30695.2]
  input   clock, // @[:@30696.4]
  input   reset, // @[:@30697.4]
  input   io_enable, // @[:@30698.4]
  output  io_done, // @[:@30698.4]
  input   io_parentAck, // @[:@30698.4]
  input   io_doneIn_0, // @[:@30698.4]
  input   io_doneIn_1, // @[:@30698.4]
  input   io_doneIn_2, // @[:@30698.4]
  output  io_enableOut_0, // @[:@30698.4]
  output  io_enableOut_1, // @[:@30698.4]
  output  io_enableOut_2, // @[:@30698.4]
  output  io_childAck_0, // @[:@30698.4]
  output  io_childAck_1, // @[:@30698.4]
  output  io_childAck_2, // @[:@30698.4]
  input   io_ctrCopyDone_0, // @[:@30698.4]
  input   io_ctrCopyDone_1, // @[:@30698.4]
  input   io_ctrCopyDone_2 // @[:@30698.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@30701.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@30701.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@30701.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@30701.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@30701.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@30701.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@30704.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@30704.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@30704.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@30704.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@30704.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@30704.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@30707.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@30707.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@30707.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@30707.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@30707.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@30707.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@30710.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@30710.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@30710.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@30710.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@30710.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@30710.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@30713.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@30713.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@30713.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@30713.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@30713.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@30713.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@30716.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@30716.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@30716.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@30716.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@30716.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@30716.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@30757.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@30757.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@30757.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@30757.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@30757.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@30757.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@30760.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@30760.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@30760.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@30760.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@30760.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@30760.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@30763.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@30763.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@30763.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@30763.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@30763.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@30763.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@30814.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@30814.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@30814.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@30814.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@30814.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@30828.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@30828.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@30828.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@30828.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@30828.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@30846.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@30846.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@30846.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@30846.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@30846.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@30883.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@30883.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@30883.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@30883.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@30883.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@30897.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@30897.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@30897.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@30897.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@30897.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@30915.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@30915.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@30915.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@30915.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@30915.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@30952.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@30952.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@30952.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@30952.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@30952.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@30966.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@30966.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@30966.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@30966.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@30966.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@30984.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@30984.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@30984.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@30984.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@30984.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@31041.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@31041.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@31041.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@31041.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@31041.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@31058.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@31058.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@31058.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@31058.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@31058.4]
  wire  _T_77; // @[Controllers.scala 80:47:@30719.4]
  wire  allDone; // @[Controllers.scala 80:47:@30720.4]
  wire  _T_151; // @[Controllers.scala 165:35:@30798.4]
  wire  _T_153; // @[Controllers.scala 165:60:@30799.4]
  wire  _T_154; // @[Controllers.scala 165:58:@30800.4]
  wire  _T_156; // @[Controllers.scala 165:76:@30801.4]
  wire  _T_157; // @[Controllers.scala 165:74:@30802.4]
  wire  _T_161; // @[Controllers.scala 165:109:@30805.4]
  wire  _T_164; // @[Controllers.scala 165:141:@30807.4]
  wire  _T_172; // @[package.scala 96:25:@30819.4 package.scala 96:25:@30820.4]
  wire  _T_176; // @[Controllers.scala 167:54:@30822.4]
  wire  _T_177; // @[Controllers.scala 167:52:@30823.4]
  wire  _T_184; // @[package.scala 96:25:@30833.4 package.scala 96:25:@30834.4]
  wire  _T_202; // @[package.scala 96:25:@30851.4 package.scala 96:25:@30852.4]
  wire  _T_206; // @[Controllers.scala 169:67:@30854.4]
  wire  _T_207; // @[Controllers.scala 169:86:@30855.4]
  wire  _T_219; // @[Controllers.scala 165:35:@30867.4]
  wire  _T_221; // @[Controllers.scala 165:60:@30868.4]
  wire  _T_222; // @[Controllers.scala 165:58:@30869.4]
  wire  _T_224; // @[Controllers.scala 165:76:@30870.4]
  wire  _T_225; // @[Controllers.scala 165:74:@30871.4]
  wire  _T_229; // @[Controllers.scala 165:109:@30874.4]
  wire  _T_232; // @[Controllers.scala 165:141:@30876.4]
  wire  _T_240; // @[package.scala 96:25:@30888.4 package.scala 96:25:@30889.4]
  wire  _T_244; // @[Controllers.scala 167:54:@30891.4]
  wire  _T_245; // @[Controllers.scala 167:52:@30892.4]
  wire  _T_252; // @[package.scala 96:25:@30902.4 package.scala 96:25:@30903.4]
  wire  _T_270; // @[package.scala 96:25:@30920.4 package.scala 96:25:@30921.4]
  wire  _T_274; // @[Controllers.scala 169:67:@30923.4]
  wire  _T_275; // @[Controllers.scala 169:86:@30924.4]
  wire  _T_287; // @[Controllers.scala 165:35:@30936.4]
  wire  _T_289; // @[Controllers.scala 165:60:@30937.4]
  wire  _T_290; // @[Controllers.scala 165:58:@30938.4]
  wire  _T_292; // @[Controllers.scala 165:76:@30939.4]
  wire  _T_293; // @[Controllers.scala 165:74:@30940.4]
  wire  _T_297; // @[Controllers.scala 165:109:@30943.4]
  wire  _T_300; // @[Controllers.scala 165:141:@30945.4]
  wire  _T_308; // @[package.scala 96:25:@30957.4 package.scala 96:25:@30958.4]
  wire  _T_312; // @[Controllers.scala 167:54:@30960.4]
  wire  _T_313; // @[Controllers.scala 167:52:@30961.4]
  wire  _T_320; // @[package.scala 96:25:@30971.4 package.scala 96:25:@30972.4]
  wire  _T_338; // @[package.scala 96:25:@30989.4 package.scala 96:25:@30990.4]
  wire  _T_342; // @[Controllers.scala 169:67:@30992.4]
  wire  _T_343; // @[Controllers.scala 169:86:@30993.4]
  wire  _T_358; // @[Controllers.scala 213:68:@31011.4]
  wire  _T_360; // @[Controllers.scala 213:90:@31013.4]
  wire  _T_362; // @[Controllers.scala 213:132:@31015.4]
  wire  _T_366; // @[Controllers.scala 213:68:@31020.4]
  wire  _T_368; // @[Controllers.scala 213:90:@31022.4]
  wire  _T_374; // @[Controllers.scala 213:68:@31028.4]
  wire  _T_376; // @[Controllers.scala 213:90:@31030.4]
  wire  _T_383; // @[package.scala 100:49:@31036.4]
  reg  _T_386; // @[package.scala 48:56:@31037.4]
  reg [31:0] _RAND_0;
  wire  _T_387; // @[package.scala 100:41:@31039.4]
  reg  _T_400; // @[package.scala 48:56:@31055.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@30701.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@30704.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@30707.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@30710.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@30713.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@30716.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@30757.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@30760.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@30763.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@30814.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@30828.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@30846.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@30883.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@30897.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@30915.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@30952.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@30966.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@30984.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@31041.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@31058.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@30719.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@30720.4]
  assign _T_151 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@30798.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@30799.4]
  assign _T_154 = _T_151 & _T_153; // @[Controllers.scala 165:58:@30800.4]
  assign _T_156 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@30801.4]
  assign _T_157 = _T_154 & _T_156; // @[Controllers.scala 165:74:@30802.4]
  assign _T_161 = _T_157 & io_enable; // @[Controllers.scala 165:109:@30805.4]
  assign _T_164 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@30807.4]
  assign _T_172 = RetimeWrapper_io_out; // @[package.scala 96:25:@30819.4 package.scala 96:25:@30820.4]
  assign _T_176 = _T_172 == 1'h0; // @[Controllers.scala 167:54:@30822.4]
  assign _T_177 = io_doneIn_0 | _T_176; // @[Controllers.scala 167:52:@30823.4]
  assign _T_184 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@30833.4 package.scala 96:25:@30834.4]
  assign _T_202 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@30851.4 package.scala 96:25:@30852.4]
  assign _T_206 = _T_202 == 1'h0; // @[Controllers.scala 169:67:@30854.4]
  assign _T_207 = _T_206 & io_enable; // @[Controllers.scala 169:86:@30855.4]
  assign _T_219 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@30867.4]
  assign _T_221 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@30868.4]
  assign _T_222 = _T_219 & _T_221; // @[Controllers.scala 165:58:@30869.4]
  assign _T_224 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@30870.4]
  assign _T_225 = _T_222 & _T_224; // @[Controllers.scala 165:74:@30871.4]
  assign _T_229 = _T_225 & io_enable; // @[Controllers.scala 165:109:@30874.4]
  assign _T_232 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@30876.4]
  assign _T_240 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@30888.4 package.scala 96:25:@30889.4]
  assign _T_244 = _T_240 == 1'h0; // @[Controllers.scala 167:54:@30891.4]
  assign _T_245 = io_doneIn_1 | _T_244; // @[Controllers.scala 167:52:@30892.4]
  assign _T_252 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@30902.4 package.scala 96:25:@30903.4]
  assign _T_270 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@30920.4 package.scala 96:25:@30921.4]
  assign _T_274 = _T_270 == 1'h0; // @[Controllers.scala 169:67:@30923.4]
  assign _T_275 = _T_274 & io_enable; // @[Controllers.scala 169:86:@30924.4]
  assign _T_287 = ~ iterDone_2_io_output; // @[Controllers.scala 165:35:@30936.4]
  assign _T_289 = io_doneIn_2 == 1'h0; // @[Controllers.scala 165:60:@30937.4]
  assign _T_290 = _T_287 & _T_289; // @[Controllers.scala 165:58:@30938.4]
  assign _T_292 = done_2_io_output == 1'h0; // @[Controllers.scala 165:76:@30939.4]
  assign _T_293 = _T_290 & _T_292; // @[Controllers.scala 165:74:@30940.4]
  assign _T_297 = _T_293 & io_enable; // @[Controllers.scala 165:109:@30943.4]
  assign _T_300 = io_ctrCopyDone_2 == 1'h0; // @[Controllers.scala 165:141:@30945.4]
  assign _T_308 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@30957.4 package.scala 96:25:@30958.4]
  assign _T_312 = _T_308 == 1'h0; // @[Controllers.scala 167:54:@30960.4]
  assign _T_313 = io_doneIn_2 | _T_312; // @[Controllers.scala 167:52:@30961.4]
  assign _T_320 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@30971.4 package.scala 96:25:@30972.4]
  assign _T_338 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@30989.4 package.scala 96:25:@30990.4]
  assign _T_342 = _T_338 == 1'h0; // @[Controllers.scala 169:67:@30992.4]
  assign _T_343 = _T_342 & io_enable; // @[Controllers.scala 169:86:@30993.4]
  assign _T_358 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@31011.4]
  assign _T_360 = _T_358 & _T_151; // @[Controllers.scala 213:90:@31013.4]
  assign _T_362 = ~ allDone; // @[Controllers.scala 213:132:@31015.4]
  assign _T_366 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@31020.4]
  assign _T_368 = _T_366 & _T_219; // @[Controllers.scala 213:90:@31022.4]
  assign _T_374 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@31028.4]
  assign _T_376 = _T_374 & _T_287; // @[Controllers.scala 213:90:@31030.4]
  assign _T_383 = allDone == 1'h0; // @[package.scala 100:49:@31036.4]
  assign _T_387 = allDone & _T_386; // @[package.scala 100:41:@31039.4]
  assign io_done = RetimeWrapper_10_io_out; // @[Controllers.scala 245:13:@31065.4]
  assign io_enableOut_0 = _T_360 & _T_362; // @[Controllers.scala 213:55:@31019.4]
  assign io_enableOut_1 = _T_368 & _T_362; // @[Controllers.scala 213:55:@31027.4]
  assign io_enableOut_2 = _T_376 & _T_362; // @[Controllers.scala 213:55:@31035.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@31006.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@31008.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@31010.4]
  assign active_0_clock = clock; // @[:@30702.4]
  assign active_0_reset = reset; // @[:@30703.4]
  assign active_0_io_input_set = _T_161 & _T_164; // @[Controllers.scala 165:32:@30809.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@30813.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@30723.4]
  assign active_1_clock = clock; // @[:@30705.4]
  assign active_1_reset = reset; // @[:@30706.4]
  assign active_1_io_input_set = _T_229 & _T_232; // @[Controllers.scala 165:32:@30878.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@30882.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@30724.4]
  assign active_2_clock = clock; // @[:@30708.4]
  assign active_2_reset = reset; // @[:@30709.4]
  assign active_2_io_input_set = _T_297 & _T_300; // @[Controllers.scala 165:32:@30947.4]
  assign active_2_io_input_reset = io_ctrCopyDone_2 | io_parentAck; // @[Controllers.scala 166:34:@30951.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@30725.4]
  assign done_0_clock = clock; // @[:@30711.4]
  assign done_0_reset = reset; // @[:@30712.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_207; // @[Controllers.scala 169:30:@30859.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@30737.4 Controllers.scala 170:32:@30866.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@30726.4]
  assign done_1_clock = clock; // @[:@30714.4]
  assign done_1_reset = reset; // @[:@30715.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_275; // @[Controllers.scala 169:30:@30928.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@30746.4 Controllers.scala 170:32:@30935.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@30727.4]
  assign done_2_clock = clock; // @[:@30717.4]
  assign done_2_reset = reset; // @[:@30718.4]
  assign done_2_io_input_set = io_ctrCopyDone_2 | _T_343; // @[Controllers.scala 169:30:@30997.4]
  assign done_2_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@30755.4 Controllers.scala 170:32:@31004.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@30728.4]
  assign iterDone_0_clock = clock; // @[:@30758.4]
  assign iterDone_0_reset = reset; // @[:@30759.4]
  assign iterDone_0_io_input_set = _T_177 & io_enable; // @[Controllers.scala 167:34:@30827.4]
  assign iterDone_0_io_input_reset = _T_184 | io_parentAck; // @[Controllers.scala 92:37:@30777.4 Controllers.scala 168:36:@30843.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@30766.4]
  assign iterDone_1_clock = clock; // @[:@30761.4]
  assign iterDone_1_reset = reset; // @[:@30762.4]
  assign iterDone_1_io_input_set = _T_245 & io_enable; // @[Controllers.scala 167:34:@30896.4]
  assign iterDone_1_io_input_reset = _T_252 | io_parentAck; // @[Controllers.scala 92:37:@30786.4 Controllers.scala 168:36:@30912.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@30767.4]
  assign iterDone_2_clock = clock; // @[:@30764.4]
  assign iterDone_2_reset = reset; // @[:@30765.4]
  assign iterDone_2_io_input_set = _T_313 & io_enable; // @[Controllers.scala 167:34:@30965.4]
  assign iterDone_2_io_input_reset = _T_320 | io_parentAck; // @[Controllers.scala 92:37:@30795.4 Controllers.scala 168:36:@30981.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@30768.4]
  assign RetimeWrapper_clock = clock; // @[:@30815.4]
  assign RetimeWrapper_reset = reset; // @[:@30816.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@30818.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@30817.4]
  assign RetimeWrapper_1_clock = clock; // @[:@30829.4]
  assign RetimeWrapper_1_reset = reset; // @[:@30830.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@30832.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@30831.4]
  assign RetimeWrapper_2_clock = clock; // @[:@30847.4]
  assign RetimeWrapper_2_reset = reset; // @[:@30848.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@30850.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@30849.4]
  assign RetimeWrapper_3_clock = clock; // @[:@30884.4]
  assign RetimeWrapper_3_reset = reset; // @[:@30885.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@30887.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@30886.4]
  assign RetimeWrapper_4_clock = clock; // @[:@30898.4]
  assign RetimeWrapper_4_reset = reset; // @[:@30899.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@30901.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@30900.4]
  assign RetimeWrapper_5_clock = clock; // @[:@30916.4]
  assign RetimeWrapper_5_reset = reset; // @[:@30917.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@30919.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@30918.4]
  assign RetimeWrapper_6_clock = clock; // @[:@30953.4]
  assign RetimeWrapper_6_reset = reset; // @[:@30954.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@30956.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@30955.4]
  assign RetimeWrapper_7_clock = clock; // @[:@30967.4]
  assign RetimeWrapper_7_reset = reset; // @[:@30968.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@30970.4]
  assign RetimeWrapper_7_io_in = io_doneIn_2; // @[package.scala 94:16:@30969.4]
  assign RetimeWrapper_8_clock = clock; // @[:@30985.4]
  assign RetimeWrapper_8_reset = reset; // @[:@30986.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@30988.4]
  assign RetimeWrapper_8_io_in = 1'h1; // @[package.scala 94:16:@30987.4]
  assign RetimeWrapper_9_clock = clock; // @[:@31042.4]
  assign RetimeWrapper_9_reset = reset; // @[:@31043.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@31045.4]
  assign RetimeWrapper_9_io_in = _T_387 | io_parentAck; // @[package.scala 94:16:@31044.4]
  assign RetimeWrapper_10_clock = clock; // @[:@31059.4]
  assign RetimeWrapper_10_reset = reset; // @[:@31060.4]
  assign RetimeWrapper_10_io_flow = io_enable; // @[package.scala 95:18:@31062.4]
  assign RetimeWrapper_10_io_in = allDone & _T_400; // @[package.scala 94:16:@31061.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_386 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_400 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_386 <= 1'h0;
    end else begin
      _T_386 <= _T_383;
    end
    if (reset) begin
      _T_400 <= 1'h0;
    end else begin
      _T_400 <= _T_383;
    end
  end
endmodule
module x329_inr_UnitPipe_sm( // @[:@31238.2]
  input   clock, // @[:@31239.4]
  input   reset, // @[:@31240.4]
  input   io_enable, // @[:@31241.4]
  output  io_done, // @[:@31241.4]
  output  io_doneLatch, // @[:@31241.4]
  input   io_ctrDone, // @[:@31241.4]
  output  io_datapathEn, // @[:@31241.4]
  output  io_ctrInc, // @[:@31241.4]
  input   io_parentAck, // @[:@31241.4]
  input   io_backpressure // @[:@31241.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@31243.4]
  wire  active_reset; // @[Controllers.scala 261:22:@31243.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@31243.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@31243.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@31243.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@31243.4]
  wire  done_clock; // @[Controllers.scala 262:20:@31246.4]
  wire  done_reset; // @[Controllers.scala 262:20:@31246.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@31246.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@31246.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@31246.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@31246.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@31300.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@31300.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@31300.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@31300.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@31300.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@31308.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@31308.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@31308.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@31308.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@31308.4]
  wire  _T_80; // @[Controllers.scala 264:48:@31251.4]
  wire  _T_81; // @[Controllers.scala 264:46:@31252.4]
  wire  _T_82; // @[Controllers.scala 264:62:@31253.4]
  wire  _T_83; // @[Controllers.scala 264:60:@31254.4]
  wire  _T_100; // @[package.scala 100:49:@31271.4]
  reg  _T_103; // @[package.scala 48:56:@31272.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 100:49:@31280.4]
  wire  _T_116; // @[Controllers.scala 283:41:@31288.4]
  wire  _T_117; // @[Controllers.scala 283:59:@31289.4]
  wire  _T_119; // @[Controllers.scala 284:37:@31292.4]
  reg  _T_125; // @[package.scala 48:56:@31296.4]
  reg [31:0] _RAND_1;
  reg  _T_142; // @[Controllers.scala 291:31:@31318.4]
  reg [31:0] _RAND_2;
  reg  _T_149; // @[package.scala 48:56:@31321.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:41:@31323.4]
  wire  _T_152; // @[Controllers.scala 292:61:@31324.4]
  wire  _T_153; // @[Controllers.scala 292:24:@31325.4]
  SRFF active ( // @[Controllers.scala 261:22:@31243.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@31246.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@31300.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@31308.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@31251.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@31252.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@31253.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@31254.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@31271.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 100:49:@31280.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@31288.4]
  assign _T_117 = _T_116 & io_enable; // @[Controllers.scala 283:59:@31289.4]
  assign _T_119 = active_io_output & io_enable; // @[Controllers.scala 284:37:@31292.4]
  assign _T_150 = done_io_output & _T_149; // @[package.scala 100:41:@31323.4]
  assign _T_152 = _T_150 ? 1'h1 : _T_142; // @[Controllers.scala 292:61:@31324.4]
  assign _T_153 = io_parentAck ? 1'h0 : _T_152; // @[Controllers.scala 292:24:@31325.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@31299.4]
  assign io_doneLatch = _T_142; // @[Controllers.scala 293:18:@31327.4]
  assign io_datapathEn = _T_117 & io_backpressure; // @[Controllers.scala 283:21:@31291.4]
  assign io_ctrInc = _T_119 & io_backpressure; // @[Controllers.scala 284:17:@31294.4]
  assign active_clock = clock; // @[:@31244.4]
  assign active_reset = reset; // @[:@31245.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@31256.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@31260.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@31261.4]
  assign done_clock = clock; // @[:@31247.4]
  assign done_reset = reset; // @[:@31248.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@31276.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@31269.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@31270.4]
  assign RetimeWrapper_clock = clock; // @[:@31301.4]
  assign RetimeWrapper_reset = reset; // @[:@31302.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@31304.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@31303.4]
  assign RetimeWrapper_1_clock = clock; // @[:@31309.4]
  assign RetimeWrapper_1_reset = reset; // @[:@31310.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@31312.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 94:16:@31311.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_125 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_142 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_149 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_142 <= 1'h0;
      end else begin
        if (_T_150) begin
          _T_142 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_108;
    end
  end
endmodule
module x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1( // @[:@31402.2]
  input  [63:0] io_in_x182_outdram_number, // @[:@31405.4]
  output        io_in_x322_valid, // @[:@31405.4]
  output [63:0] io_in_x322_bits_addr, // @[:@31405.4]
  output [31:0] io_in_x322_bits_size, // @[:@31405.4]
  input         io_sigsIn_backpressure, // @[:@31405.4]
  input         io_sigsIn_datapathEn, // @[:@31405.4]
  input         io_rr // @[:@31405.4]
);
  wire [96:0] x326_tuple; // @[Cat.scala 30:58:@31419.4]
  wire  _T_135; // @[implicits.scala 55:10:@31422.4]
  assign x326_tuple = {33'h7e9000,io_in_x182_outdram_number}; // @[Cat.scala 30:58:@31419.4]
  assign _T_135 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@31422.4]
  assign io_in_x322_valid = _T_135 & io_sigsIn_backpressure; // @[sm_x329_inr_UnitPipe.scala 65:18:@31425.4]
  assign io_in_x322_bits_addr = x326_tuple[63:0]; // @[sm_x329_inr_UnitPipe.scala 66:22:@31427.4]
  assign io_in_x322_bits_size = x326_tuple[95:64]; // @[sm_x329_inr_UnitPipe.scala 67:22:@31429.4]
endmodule
module FF_13( // @[:@31431.2]
  input         clock, // @[:@31432.4]
  input         reset, // @[:@31433.4]
  output [22:0] io_rPort_0_output_0, // @[:@31434.4]
  input  [22:0] io_wPort_0_data_0, // @[:@31434.4]
  input         io_wPort_0_reset, // @[:@31434.4]
  input         io_wPort_0_en_0 // @[:@31434.4]
);
  reg [22:0] ff; // @[MemPrimitives.scala 321:19:@31449.4]
  reg [31:0] _RAND_0;
  wire [22:0] _T_68; // @[MemPrimitives.scala 325:32:@31451.4]
  wire [22:0] _T_69; // @[MemPrimitives.scala 325:12:@31452.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@31451.4]
  assign _T_69 = io_wPort_0_reset ? 23'h0 : _T_68; // @[MemPrimitives.scala 325:12:@31452.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@31454.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[22:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 23'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 23'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_5( // @[:@31469.2]
  input         clock, // @[:@31470.4]
  input         reset, // @[:@31471.4]
  input         io_input_reset, // @[:@31472.4]
  input         io_input_enable, // @[:@31472.4]
  output [22:0] io_output_count_0, // @[:@31472.4]
  output        io_output_oobs_0, // @[:@31472.4]
  output        io_output_done // @[:@31472.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@31485.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@31485.4]
  wire [22:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@31485.4]
  wire [22:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@31485.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@31485.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@31485.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@31501.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@31501.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@31501.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@31501.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@31501.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@31501.4]
  wire  _T_36; // @[Counter.scala 264:45:@31504.4]
  wire [22:0] _T_48; // @[Counter.scala 287:52:@31529.4]
  wire [23:0] _T_50; // @[Counter.scala 291:33:@31530.4]
  wire [22:0] _T_51; // @[Counter.scala 291:33:@31531.4]
  wire [22:0] _T_52; // @[Counter.scala 291:33:@31532.4]
  wire  _T_57; // @[Counter.scala 293:18:@31534.4]
  wire [22:0] _T_68; // @[Counter.scala 299:115:@31542.4]
  wire [22:0] _T_71; // @[Counter.scala 299:152:@31545.4]
  wire [22:0] _T_72; // @[Counter.scala 299:74:@31546.4]
  wire  _T_75; // @[Counter.scala 322:102:@31550.4]
  wire  _T_77; // @[Counter.scala 322:130:@31551.4]
  FF_13 bases_0 ( // @[Counter.scala 261:53:@31485.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@31501.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@31504.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@31529.4]
  assign _T_50 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@31530.4]
  assign _T_51 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@31531.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@31532.4]
  assign _T_57 = $signed(_T_52) >= $signed(23'sh1fa400); // @[Counter.scala 293:18:@31534.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@31542.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@31545.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@31546.4]
  assign _T_75 = $signed(_T_48) < $signed(23'sh0); // @[Counter.scala 322:102:@31550.4]
  assign _T_77 = $signed(_T_48) >= $signed(23'sh1fa400); // @[Counter.scala 322:130:@31551.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@31549.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@31553.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@31555.4]
  assign bases_0_clock = clock; // @[:@31486.4]
  assign bases_0_reset = reset; // @[:@31487.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 23'h0 : _T_72; // @[Counter.scala 299:31:@31548.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@31527.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@31528.4]
  assign SRFF_clock = clock; // @[:@31502.4]
  assign SRFF_reset = reset; // @[:@31503.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@31506.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@31508.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@31509.4]
endmodule
module x331_ctrchain( // @[:@31560.2]
  input         clock, // @[:@31561.4]
  input         reset, // @[:@31562.4]
  input         io_input_reset, // @[:@31563.4]
  input         io_input_enable, // @[:@31563.4]
  output [22:0] io_output_counts_0, // @[:@31563.4]
  output        io_output_oobs_0, // @[:@31563.4]
  output        io_output_done // @[:@31563.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@31565.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@31565.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@31565.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@31565.4]
  wire [22:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@31565.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@31565.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@31565.4]
  reg  wasDone; // @[Counter.scala 542:24:@31574.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 546:69:@31580.4]
  wire  _T_47; // @[Counter.scala 546:80:@31581.4]
  reg  doneLatch; // @[Counter.scala 550:26:@31586.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 551:48:@31587.4]
  wire  _T_55; // @[Counter.scala 551:19:@31588.4]
  SingleCounter_5 ctrs_0 ( // @[Counter.scala 513:46:@31565.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 546:69:@31580.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 546:80:@31581.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@31587.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 551:19:@31588.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@31590.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@31592.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 546:18:@31583.4]
  assign ctrs_0_clock = clock; // @[:@31566.4]
  assign ctrs_0_reset = reset; // @[:@31567.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@31571.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@31572.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x338_inr_Foreach_sm( // @[:@31780.2]
  input   clock, // @[:@31781.4]
  input   reset, // @[:@31782.4]
  input   io_enable, // @[:@31783.4]
  output  io_done, // @[:@31783.4]
  output  io_doneLatch, // @[:@31783.4]
  input   io_ctrDone, // @[:@31783.4]
  output  io_datapathEn, // @[:@31783.4]
  output  io_ctrInc, // @[:@31783.4]
  output  io_ctrRst, // @[:@31783.4]
  input   io_parentAck, // @[:@31783.4]
  input   io_backpressure, // @[:@31783.4]
  input   io_break // @[:@31783.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@31785.4]
  wire  active_reset; // @[Controllers.scala 261:22:@31785.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@31785.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@31785.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@31785.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@31785.4]
  wire  done_clock; // @[Controllers.scala 262:20:@31788.4]
  wire  done_reset; // @[Controllers.scala 262:20:@31788.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@31788.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@31788.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@31788.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@31788.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@31822.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@31822.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@31822.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@31822.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@31822.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@31844.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@31844.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@31844.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@31844.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@31844.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@31856.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@31856.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@31856.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@31856.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@31856.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@31864.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@31864.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@31864.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@31864.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@31864.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@31880.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@31880.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@31880.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@31880.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@31880.4]
  wire  _T_80; // @[Controllers.scala 264:48:@31793.4]
  wire  _T_81; // @[Controllers.scala 264:46:@31794.4]
  wire  _T_82; // @[Controllers.scala 264:62:@31795.4]
  wire  _T_83; // @[Controllers.scala 264:60:@31796.4]
  wire  _T_100; // @[package.scala 100:49:@31813.4]
  reg  _T_103; // @[package.scala 48:56:@31814.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@31827.4 package.scala 96:25:@31828.4]
  wire  _T_110; // @[package.scala 100:49:@31829.4]
  reg  _T_113; // @[package.scala 48:56:@31830.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@31832.4]
  wire  _T_118; // @[Controllers.scala 283:41:@31837.4]
  wire  _T_119; // @[Controllers.scala 283:59:@31838.4]
  wire  _T_121; // @[Controllers.scala 284:37:@31841.4]
  wire  _T_124; // @[package.scala 96:25:@31849.4 package.scala 96:25:@31850.4]
  wire  _T_126; // @[package.scala 100:49:@31851.4]
  reg  _T_129; // @[package.scala 48:56:@31852.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@31874.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@31876.4]
  reg  _T_153; // @[package.scala 48:56:@31877.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@31885.4 package.scala 96:25:@31886.4]
  wire  _T_158; // @[Controllers.scala 292:61:@31887.4]
  wire  _T_159; // @[Controllers.scala 292:24:@31888.4]
  SRFF active ( // @[Controllers.scala 261:22:@31785.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@31788.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@31822.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@31844.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@31856.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@31864.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@31880.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@31793.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@31794.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@31795.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@31796.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@31813.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@31827.4 package.scala 96:25:@31828.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@31829.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@31832.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@31837.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@31838.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@31841.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@31849.4 package.scala 96:25:@31850.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@31851.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@31876.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@31885.4 package.scala 96:25:@31886.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@31887.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@31888.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@31855.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@31890.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@31840.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@31843.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@31835.4]
  assign active_clock = clock; // @[:@31786.4]
  assign active_reset = reset; // @[:@31787.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@31798.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@31802.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@31803.4]
  assign done_clock = clock; // @[:@31789.4]
  assign done_reset = reset; // @[:@31790.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@31818.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@31811.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@31812.4]
  assign RetimeWrapper_clock = clock; // @[:@31823.4]
  assign RetimeWrapper_reset = reset; // @[:@31824.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@31826.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@31825.4]
  assign RetimeWrapper_1_clock = clock; // @[:@31845.4]
  assign RetimeWrapper_1_reset = reset; // @[:@31846.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@31848.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@31847.4]
  assign RetimeWrapper_2_clock = clock; // @[:@31857.4]
  assign RetimeWrapper_2_reset = reset; // @[:@31858.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@31860.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@31859.4]
  assign RetimeWrapper_3_clock = clock; // @[:@31865.4]
  assign RetimeWrapper_3_reset = reset; // @[:@31866.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@31868.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@31867.4]
  assign RetimeWrapper_4_clock = clock; // @[:@31881.4]
  assign RetimeWrapper_4_reset = reset; // @[:@31882.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@31884.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@31883.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x338_inr_Foreach_kernelx338_inr_Foreach_concrete1( // @[:@32097.2]
  input         clock, // @[:@32098.4]
  input         reset, // @[:@32099.4]
  output        io_in_x323_valid, // @[:@32100.4]
  output [31:0] io_in_x323_bits_wdata_0, // @[:@32100.4]
  output        io_in_x323_bits_wstrb, // @[:@32100.4]
  output [20:0] io_in_x186_outbuf_0_rPort_0_ofs_0, // @[:@32100.4]
  output        io_in_x186_outbuf_0_rPort_0_en_0, // @[:@32100.4]
  output        io_in_x186_outbuf_0_rPort_0_backpressure, // @[:@32100.4]
  input  [31:0] io_in_x186_outbuf_0_rPort_0_output_0, // @[:@32100.4]
  input         io_sigsIn_backpressure, // @[:@32100.4]
  input         io_sigsIn_datapathEn, // @[:@32100.4]
  input         io_sigsIn_break, // @[:@32100.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@32100.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@32100.4]
  input         io_rr // @[:@32100.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@32127.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@32127.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@32156.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@32156.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@32156.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@32156.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@32156.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32165.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32165.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32165.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@32165.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@32165.4]
  wire  b333; // @[sm_x338_inr_Foreach.scala 62:18:@32135.4]
  wire  _T_274; // @[sm_x338_inr_Foreach.scala 67:129:@32139.4]
  wire  _T_278; // @[implicits.scala 55:10:@32142.4]
  wire  _T_279; // @[sm_x338_inr_Foreach.scala 67:146:@32143.4]
  wire [32:0] x336_tuple; // @[Cat.scala 30:58:@32153.4]
  wire  _T_290; // @[package.scala 96:25:@32170.4 package.scala 96:25:@32171.4]
  wire  _T_292; // @[implicits.scala 55:10:@32172.4]
  wire  x505_b333_D2; // @[package.scala 96:25:@32161.4 package.scala 96:25:@32162.4]
  wire  _T_293; // @[sm_x338_inr_Foreach.scala 74:112:@32173.4]
  wire [31:0] b332_number; // @[Math.scala 723:22:@32132.4 Math.scala 724:14:@32133.4]
  _ _ ( // @[Math.scala 720:24:@32127.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@32156.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@32165.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign b333 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x338_inr_Foreach.scala 62:18:@32135.4]
  assign _T_274 = ~ io_sigsIn_break; // @[sm_x338_inr_Foreach.scala 67:129:@32139.4]
  assign _T_278 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@32142.4]
  assign _T_279 = _T_274 & _T_278; // @[sm_x338_inr_Foreach.scala 67:146:@32143.4]
  assign x336_tuple = {1'h1,io_in_x186_outbuf_0_rPort_0_output_0}; // @[Cat.scala 30:58:@32153.4]
  assign _T_290 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@32170.4 package.scala 96:25:@32171.4]
  assign _T_292 = io_rr ? _T_290 : 1'h0; // @[implicits.scala 55:10:@32172.4]
  assign x505_b333_D2 = RetimeWrapper_io_out; // @[package.scala 96:25:@32161.4 package.scala 96:25:@32162.4]
  assign _T_293 = _T_292 & x505_b333_D2; // @[sm_x338_inr_Foreach.scala 74:112:@32173.4]
  assign b332_number = __io_result; // @[Math.scala 723:22:@32132.4 Math.scala 724:14:@32133.4]
  assign io_in_x323_valid = _T_293 & io_sigsIn_backpressure; // @[sm_x338_inr_Foreach.scala 74:18:@32175.4]
  assign io_in_x323_bits_wdata_0 = x336_tuple[31:0]; // @[sm_x338_inr_Foreach.scala 75:26:@32177.4]
  assign io_in_x323_bits_wstrb = x336_tuple[32]; // @[sm_x338_inr_Foreach.scala 76:23:@32179.4]
  assign io_in_x186_outbuf_0_rPort_0_ofs_0 = b332_number[20:0]; // @[MemInterfaceType.scala 107:54:@32146.4]
  assign io_in_x186_outbuf_0_rPort_0_en_0 = _T_279 & b333; // @[MemInterfaceType.scala 110:79:@32148.4]
  assign io_in_x186_outbuf_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32147.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@32130.4]
  assign RetimeWrapper_clock = clock; // @[:@32157.4]
  assign RetimeWrapper_reset = reset; // @[:@32158.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32160.4]
  assign RetimeWrapper_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@32159.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32166.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32167.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32169.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32168.4]
endmodule
module x342_inr_UnitPipe_sm( // @[:@32335.2]
  input   clock, // @[:@32336.4]
  input   reset, // @[:@32337.4]
  input   io_enable, // @[:@32338.4]
  output  io_done, // @[:@32338.4]
  output  io_doneLatch, // @[:@32338.4]
  input   io_ctrDone, // @[:@32338.4]
  output  io_datapathEn, // @[:@32338.4]
  output  io_ctrInc, // @[:@32338.4]
  input   io_parentAck // @[:@32338.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@32340.4]
  wire  active_reset; // @[Controllers.scala 261:22:@32340.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@32340.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@32340.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@32340.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@32340.4]
  wire  done_clock; // @[Controllers.scala 262:20:@32343.4]
  wire  done_reset; // @[Controllers.scala 262:20:@32343.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@32343.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@32343.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@32343.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@32343.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@32377.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@32377.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@32377.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@32377.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@32377.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32399.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32399.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32399.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@32399.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@32399.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@32411.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@32411.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@32411.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@32411.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@32411.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@32419.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@32419.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@32419.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@32419.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@32419.4]
  wire  _T_80; // @[Controllers.scala 264:48:@32348.4]
  wire  _T_81; // @[Controllers.scala 264:46:@32349.4]
  wire  _T_82; // @[Controllers.scala 264:62:@32350.4]
  wire  _T_100; // @[package.scala 100:49:@32368.4]
  reg  _T_103; // @[package.scala 48:56:@32369.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@32392.4]
  wire  _T_124; // @[package.scala 96:25:@32404.4 package.scala 96:25:@32405.4]
  wire  _T_126; // @[package.scala 100:49:@32406.4]
  reg  _T_129; // @[package.scala 48:56:@32407.4]
  reg [31:0] _RAND_1;
  reg  _T_146; // @[Controllers.scala 291:31:@32429.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@32431.4]
  reg  _T_153; // @[package.scala 48:56:@32432.4]
  reg [31:0] _RAND_3;
  wire  _T_154; // @[package.scala 100:41:@32434.4]
  wire  _T_156; // @[Controllers.scala 292:61:@32435.4]
  wire  _T_157; // @[Controllers.scala 292:24:@32436.4]
  SRFF active ( // @[Controllers.scala 261:22:@32340.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@32343.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@32377.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@32399.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@32411.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@32419.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@32348.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@32349.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@32350.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@32368.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@32392.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@32404.4 package.scala 96:25:@32405.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@32406.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@32431.4]
  assign _T_154 = done_io_output & _T_153; // @[package.scala 100:41:@32434.4]
  assign _T_156 = _T_154 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@32435.4]
  assign _T_157 = io_parentAck ? 1'h0 : _T_156; // @[Controllers.scala 292:24:@32436.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@32410.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@32438.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@32395.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@32398.4]
  assign active_clock = clock; // @[:@32341.4]
  assign active_reset = reset; // @[:@32342.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@32353.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@32357.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@32358.4]
  assign done_clock = clock; // @[:@32344.4]
  assign done_reset = reset; // @[:@32345.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@32373.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@32366.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@32367.4]
  assign RetimeWrapper_clock = clock; // @[:@32378.4]
  assign RetimeWrapper_reset = reset; // @[:@32379.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@32381.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@32380.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32400.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32401.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@32403.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@32402.4]
  assign RetimeWrapper_2_clock = clock; // @[:@32412.4]
  assign RetimeWrapper_2_reset = reset; // @[:@32413.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@32415.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@32414.4]
  assign RetimeWrapper_3_clock = clock; // @[:@32420.4]
  assign RetimeWrapper_3_reset = reset; // @[:@32421.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@32423.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@32422.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_154) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x342_inr_UnitPipe_kernelx342_inr_UnitPipe_concrete1( // @[:@32513.2]
  output  io_in_x324_ready, // @[:@32516.4]
  input   io_sigsIn_datapathEn // @[:@32516.4]
);
  assign io_in_x324_ready = io_sigsIn_datapathEn; // @[sm_x342_inr_UnitPipe.scala 57:18:@32528.4]
endmodule
module x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1( // @[:@32531.2]
  input         clock, // @[:@32532.4]
  input         reset, // @[:@32533.4]
  output        io_in_x324_ready, // @[:@32534.4]
  input         io_in_x324_valid, // @[:@32534.4]
  input         io_in_x323_ready, // @[:@32534.4]
  output        io_in_x323_valid, // @[:@32534.4]
  output [31:0] io_in_x323_bits_wdata_0, // @[:@32534.4]
  output        io_in_x323_bits_wstrb, // @[:@32534.4]
  input  [63:0] io_in_x182_outdram_number, // @[:@32534.4]
  output [20:0] io_in_x186_outbuf_0_rPort_0_ofs_0, // @[:@32534.4]
  output        io_in_x186_outbuf_0_rPort_0_en_0, // @[:@32534.4]
  output        io_in_x186_outbuf_0_rPort_0_backpressure, // @[:@32534.4]
  input  [31:0] io_in_x186_outbuf_0_rPort_0_output_0, // @[:@32534.4]
  input         io_in_x322_ready, // @[:@32534.4]
  output        io_in_x322_valid, // @[:@32534.4]
  output [63:0] io_in_x322_bits_addr, // @[:@32534.4]
  output [31:0] io_in_x322_bits_size, // @[:@32534.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@32534.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@32534.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@32534.4]
  input         io_sigsIn_smChildAcks_0, // @[:@32534.4]
  input         io_sigsIn_smChildAcks_1, // @[:@32534.4]
  input         io_sigsIn_smChildAcks_2, // @[:@32534.4]
  output        io_sigsOut_smDoneIn_0, // @[:@32534.4]
  output        io_sigsOut_smDoneIn_1, // @[:@32534.4]
  output        io_sigsOut_smDoneIn_2, // @[:@32534.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@32534.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@32534.4]
  output        io_sigsOut_smCtrCopyDone_2, // @[:@32534.4]
  input         io_rr // @[:@32534.4]
);
  wire  x329_inr_UnitPipe_sm_clock; // @[sm_x329_inr_UnitPipe.scala 33:18:@32601.4]
  wire  x329_inr_UnitPipe_sm_reset; // @[sm_x329_inr_UnitPipe.scala 33:18:@32601.4]
  wire  x329_inr_UnitPipe_sm_io_enable; // @[sm_x329_inr_UnitPipe.scala 33:18:@32601.4]
  wire  x329_inr_UnitPipe_sm_io_done; // @[sm_x329_inr_UnitPipe.scala 33:18:@32601.4]
  wire  x329_inr_UnitPipe_sm_io_doneLatch; // @[sm_x329_inr_UnitPipe.scala 33:18:@32601.4]
  wire  x329_inr_UnitPipe_sm_io_ctrDone; // @[sm_x329_inr_UnitPipe.scala 33:18:@32601.4]
  wire  x329_inr_UnitPipe_sm_io_datapathEn; // @[sm_x329_inr_UnitPipe.scala 33:18:@32601.4]
  wire  x329_inr_UnitPipe_sm_io_ctrInc; // @[sm_x329_inr_UnitPipe.scala 33:18:@32601.4]
  wire  x329_inr_UnitPipe_sm_io_parentAck; // @[sm_x329_inr_UnitPipe.scala 33:18:@32601.4]
  wire  x329_inr_UnitPipe_sm_io_backpressure; // @[sm_x329_inr_UnitPipe.scala 33:18:@32601.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@32658.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@32658.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@32658.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@32658.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@32658.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32666.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32666.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32666.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@32666.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@32666.4]
  wire [63:0] x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_in_x182_outdram_number; // @[sm_x329_inr_UnitPipe.scala 69:24:@32696.4]
  wire  x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_in_x322_valid; // @[sm_x329_inr_UnitPipe.scala 69:24:@32696.4]
  wire [63:0] x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_in_x322_bits_addr; // @[sm_x329_inr_UnitPipe.scala 69:24:@32696.4]
  wire [31:0] x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_in_x322_bits_size; // @[sm_x329_inr_UnitPipe.scala 69:24:@32696.4]
  wire  x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x329_inr_UnitPipe.scala 69:24:@32696.4]
  wire  x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x329_inr_UnitPipe.scala 69:24:@32696.4]
  wire  x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_rr; // @[sm_x329_inr_UnitPipe.scala 69:24:@32696.4]
  wire  x331_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@32764.4]
  wire  x331_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@32764.4]
  wire  x331_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@32764.4]
  wire  x331_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@32764.4]
  wire [22:0] x331_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@32764.4]
  wire  x331_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@32764.4]
  wire  x331_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@32764.4]
  wire  x338_inr_Foreach_sm_clock; // @[sm_x338_inr_Foreach.scala 33:18:@32817.4]
  wire  x338_inr_Foreach_sm_reset; // @[sm_x338_inr_Foreach.scala 33:18:@32817.4]
  wire  x338_inr_Foreach_sm_io_enable; // @[sm_x338_inr_Foreach.scala 33:18:@32817.4]
  wire  x338_inr_Foreach_sm_io_done; // @[sm_x338_inr_Foreach.scala 33:18:@32817.4]
  wire  x338_inr_Foreach_sm_io_doneLatch; // @[sm_x338_inr_Foreach.scala 33:18:@32817.4]
  wire  x338_inr_Foreach_sm_io_ctrDone; // @[sm_x338_inr_Foreach.scala 33:18:@32817.4]
  wire  x338_inr_Foreach_sm_io_datapathEn; // @[sm_x338_inr_Foreach.scala 33:18:@32817.4]
  wire  x338_inr_Foreach_sm_io_ctrInc; // @[sm_x338_inr_Foreach.scala 33:18:@32817.4]
  wire  x338_inr_Foreach_sm_io_ctrRst; // @[sm_x338_inr_Foreach.scala 33:18:@32817.4]
  wire  x338_inr_Foreach_sm_io_parentAck; // @[sm_x338_inr_Foreach.scala 33:18:@32817.4]
  wire  x338_inr_Foreach_sm_io_backpressure; // @[sm_x338_inr_Foreach.scala 33:18:@32817.4]
  wire  x338_inr_Foreach_sm_io_break; // @[sm_x338_inr_Foreach.scala 33:18:@32817.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@32845.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@32845.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@32845.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@32845.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@32845.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@32885.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@32885.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@32885.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@32885.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@32885.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@32893.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@32893.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@32893.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@32893.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@32893.4]
  wire  x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_clock; // @[sm_x338_inr_Foreach.scala 78:24:@32928.4]
  wire  x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_reset; // @[sm_x338_inr_Foreach.scala 78:24:@32928.4]
  wire  x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x323_valid; // @[sm_x338_inr_Foreach.scala 78:24:@32928.4]
  wire [31:0] x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x323_bits_wdata_0; // @[sm_x338_inr_Foreach.scala 78:24:@32928.4]
  wire  x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x323_bits_wstrb; // @[sm_x338_inr_Foreach.scala 78:24:@32928.4]
  wire [20:0] x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x186_outbuf_0_rPort_0_ofs_0; // @[sm_x338_inr_Foreach.scala 78:24:@32928.4]
  wire  x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x186_outbuf_0_rPort_0_en_0; // @[sm_x338_inr_Foreach.scala 78:24:@32928.4]
  wire  x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x186_outbuf_0_rPort_0_backpressure; // @[sm_x338_inr_Foreach.scala 78:24:@32928.4]
  wire [31:0] x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x186_outbuf_0_rPort_0_output_0; // @[sm_x338_inr_Foreach.scala 78:24:@32928.4]
  wire  x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x338_inr_Foreach.scala 78:24:@32928.4]
  wire  x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x338_inr_Foreach.scala 78:24:@32928.4]
  wire  x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x338_inr_Foreach.scala 78:24:@32928.4]
  wire [31:0] x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x338_inr_Foreach.scala 78:24:@32928.4]
  wire  x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x338_inr_Foreach.scala 78:24:@32928.4]
  wire  x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_rr; // @[sm_x338_inr_Foreach.scala 78:24:@32928.4]
  wire  x342_inr_UnitPipe_sm_clock; // @[sm_x342_inr_UnitPipe.scala 32:18:@33048.4]
  wire  x342_inr_UnitPipe_sm_reset; // @[sm_x342_inr_UnitPipe.scala 32:18:@33048.4]
  wire  x342_inr_UnitPipe_sm_io_enable; // @[sm_x342_inr_UnitPipe.scala 32:18:@33048.4]
  wire  x342_inr_UnitPipe_sm_io_done; // @[sm_x342_inr_UnitPipe.scala 32:18:@33048.4]
  wire  x342_inr_UnitPipe_sm_io_doneLatch; // @[sm_x342_inr_UnitPipe.scala 32:18:@33048.4]
  wire  x342_inr_UnitPipe_sm_io_ctrDone; // @[sm_x342_inr_UnitPipe.scala 32:18:@33048.4]
  wire  x342_inr_UnitPipe_sm_io_datapathEn; // @[sm_x342_inr_UnitPipe.scala 32:18:@33048.4]
  wire  x342_inr_UnitPipe_sm_io_ctrInc; // @[sm_x342_inr_UnitPipe.scala 32:18:@33048.4]
  wire  x342_inr_UnitPipe_sm_io_parentAck; // @[sm_x342_inr_UnitPipe.scala 32:18:@33048.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@33105.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@33105.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@33105.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@33105.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@33105.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@33113.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@33113.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@33113.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@33113.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@33113.4]
  wire  x342_inr_UnitPipe_kernelx342_inr_UnitPipe_concrete1_io_in_x324_ready; // @[sm_x342_inr_UnitPipe.scala 60:24:@33143.4]
  wire  x342_inr_UnitPipe_kernelx342_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x342_inr_UnitPipe.scala 60:24:@33143.4]
  wire  _T_359; // @[package.scala 100:49:@32629.4]
  reg  _T_362; // @[package.scala 48:56:@32630.4]
  reg [31:0] _RAND_0;
  wire  _T_375; // @[package.scala 96:25:@32663.4 package.scala 96:25:@32664.4]
  wire  _T_381; // @[package.scala 96:25:@32671.4 package.scala 96:25:@32672.4]
  wire  _T_384; // @[SpatialBlocks.scala 138:93:@32674.4]
  wire  _T_454; // @[package.scala 96:25:@32850.4 package.scala 96:25:@32851.4]
  wire  _T_468; // @[package.scala 96:25:@32890.4 package.scala 96:25:@32891.4]
  wire  _T_474; // @[package.scala 96:25:@32898.4 package.scala 96:25:@32899.4]
  wire  _T_477; // @[SpatialBlocks.scala 138:93:@32901.4]
  wire  _T_479; // @[SpatialBlocks.scala 157:36:@32910.4]
  wire  _T_480; // @[SpatialBlocks.scala 157:78:@32911.4]
  wire  _T_547; // @[package.scala 100:49:@33076.4]
  reg  _T_550; // @[package.scala 48:56:@33077.4]
  reg [31:0] _RAND_1;
  wire  x342_inr_UnitPipe_sigsIn_forwardpressure; // @[sm_x343_outr_UnitPipe.scala 101:55:@33083.4]
  wire  _T_563; // @[package.scala 96:25:@33110.4 package.scala 96:25:@33111.4]
  wire  _T_569; // @[package.scala 96:25:@33118.4 package.scala 96:25:@33119.4]
  wire  _T_572; // @[SpatialBlocks.scala 138:93:@33121.4]
  wire  x342_inr_UnitPipe_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@33122.4]
  x329_inr_UnitPipe_sm x329_inr_UnitPipe_sm ( // @[sm_x329_inr_UnitPipe.scala 33:18:@32601.4]
    .clock(x329_inr_UnitPipe_sm_clock),
    .reset(x329_inr_UnitPipe_sm_reset),
    .io_enable(x329_inr_UnitPipe_sm_io_enable),
    .io_done(x329_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x329_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x329_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x329_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x329_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x329_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x329_inr_UnitPipe_sm_io_backpressure)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@32658.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@32666.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1 x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1 ( // @[sm_x329_inr_UnitPipe.scala 69:24:@32696.4]
    .io_in_x182_outdram_number(x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_in_x182_outdram_number),
    .io_in_x322_valid(x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_in_x322_valid),
    .io_in_x322_bits_addr(x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_in_x322_bits_addr),
    .io_in_x322_bits_size(x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_in_x322_bits_size),
    .io_sigsIn_backpressure(x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_rr(x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_rr)
  );
  x331_ctrchain x331_ctrchain ( // @[SpatialBlocks.scala 37:22:@32764.4]
    .clock(x331_ctrchain_clock),
    .reset(x331_ctrchain_reset),
    .io_input_reset(x331_ctrchain_io_input_reset),
    .io_input_enable(x331_ctrchain_io_input_enable),
    .io_output_counts_0(x331_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x331_ctrchain_io_output_oobs_0),
    .io_output_done(x331_ctrchain_io_output_done)
  );
  x338_inr_Foreach_sm x338_inr_Foreach_sm ( // @[sm_x338_inr_Foreach.scala 33:18:@32817.4]
    .clock(x338_inr_Foreach_sm_clock),
    .reset(x338_inr_Foreach_sm_reset),
    .io_enable(x338_inr_Foreach_sm_io_enable),
    .io_done(x338_inr_Foreach_sm_io_done),
    .io_doneLatch(x338_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x338_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x338_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x338_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x338_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x338_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x338_inr_Foreach_sm_io_backpressure),
    .io_break(x338_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@32845.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@32885.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@32893.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x338_inr_Foreach_kernelx338_inr_Foreach_concrete1 x338_inr_Foreach_kernelx338_inr_Foreach_concrete1 ( // @[sm_x338_inr_Foreach.scala 78:24:@32928.4]
    .clock(x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_clock),
    .reset(x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_reset),
    .io_in_x323_valid(x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x323_valid),
    .io_in_x323_bits_wdata_0(x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x323_bits_wdata_0),
    .io_in_x323_bits_wstrb(x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x323_bits_wstrb),
    .io_in_x186_outbuf_0_rPort_0_ofs_0(x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x186_outbuf_0_rPort_0_ofs_0),
    .io_in_x186_outbuf_0_rPort_0_en_0(x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x186_outbuf_0_rPort_0_en_0),
    .io_in_x186_outbuf_0_rPort_0_backpressure(x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x186_outbuf_0_rPort_0_backpressure),
    .io_in_x186_outbuf_0_rPort_0_output_0(x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x186_outbuf_0_rPort_0_output_0),
    .io_sigsIn_backpressure(x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_rr)
  );
  x342_inr_UnitPipe_sm x342_inr_UnitPipe_sm ( // @[sm_x342_inr_UnitPipe.scala 32:18:@33048.4]
    .clock(x342_inr_UnitPipe_sm_clock),
    .reset(x342_inr_UnitPipe_sm_reset),
    .io_enable(x342_inr_UnitPipe_sm_io_enable),
    .io_done(x342_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x342_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x342_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x342_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x342_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x342_inr_UnitPipe_sm_io_parentAck)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@33105.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@33113.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x342_inr_UnitPipe_kernelx342_inr_UnitPipe_concrete1 x342_inr_UnitPipe_kernelx342_inr_UnitPipe_concrete1 ( // @[sm_x342_inr_UnitPipe.scala 60:24:@33143.4]
    .io_in_x324_ready(x342_inr_UnitPipe_kernelx342_inr_UnitPipe_concrete1_io_in_x324_ready),
    .io_sigsIn_datapathEn(x342_inr_UnitPipe_kernelx342_inr_UnitPipe_concrete1_io_sigsIn_datapathEn)
  );
  assign _T_359 = x329_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@32629.4]
  assign _T_375 = RetimeWrapper_io_out; // @[package.scala 96:25:@32663.4 package.scala 96:25:@32664.4]
  assign _T_381 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@32671.4 package.scala 96:25:@32672.4]
  assign _T_384 = ~ _T_381; // @[SpatialBlocks.scala 138:93:@32674.4]
  assign _T_454 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@32850.4 package.scala 96:25:@32851.4]
  assign _T_468 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@32890.4 package.scala 96:25:@32891.4]
  assign _T_474 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@32898.4 package.scala 96:25:@32899.4]
  assign _T_477 = ~ _T_474; // @[SpatialBlocks.scala 138:93:@32901.4]
  assign _T_479 = x338_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@32910.4]
  assign _T_480 = ~ x338_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@32911.4]
  assign _T_547 = x342_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@33076.4]
  assign x342_inr_UnitPipe_sigsIn_forwardpressure = io_in_x324_valid | x342_inr_UnitPipe_sm_io_doneLatch; // @[sm_x343_outr_UnitPipe.scala 101:55:@33083.4]
  assign _T_563 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@33110.4 package.scala 96:25:@33111.4]
  assign _T_569 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@33118.4 package.scala 96:25:@33119.4]
  assign _T_572 = ~ _T_569; // @[SpatialBlocks.scala 138:93:@33121.4]
  assign x342_inr_UnitPipe_sigsIn_baseEn = _T_563 & _T_572; // @[SpatialBlocks.scala 138:90:@33122.4]
  assign io_in_x324_ready = x342_inr_UnitPipe_kernelx342_inr_UnitPipe_concrete1_io_in_x324_ready; // @[sm_x342_inr_UnitPipe.scala 46:23:@33179.4]
  assign io_in_x323_valid = x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x323_valid; // @[sm_x338_inr_Foreach.scala 49:23:@32978.4]
  assign io_in_x323_bits_wdata_0 = x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x323_bits_wdata_0; // @[sm_x338_inr_Foreach.scala 49:23:@32977.4]
  assign io_in_x323_bits_wstrb = x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x323_bits_wstrb; // @[sm_x338_inr_Foreach.scala 49:23:@32976.4]
  assign io_in_x186_outbuf_0_rPort_0_ofs_0 = x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x186_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@32983.4]
  assign io_in_x186_outbuf_0_rPort_0_en_0 = x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x186_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@32982.4]
  assign io_in_x186_outbuf_0_rPort_0_backpressure = x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x186_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@32981.4]
  assign io_in_x322_valid = x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_in_x322_valid; // @[sm_x329_inr_UnitPipe.scala 50:23:@32735.4]
  assign io_in_x322_bits_addr = x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_in_x322_bits_addr; // @[sm_x329_inr_UnitPipe.scala 50:23:@32734.4]
  assign io_in_x322_bits_size = x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_in_x322_bits_size; // @[sm_x329_inr_UnitPipe.scala 50:23:@32733.4]
  assign io_sigsOut_smDoneIn_0 = x329_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@32681.4]
  assign io_sigsOut_smDoneIn_1 = x338_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@32908.4]
  assign io_sigsOut_smDoneIn_2 = x342_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@33128.4]
  assign io_sigsOut_smCtrCopyDone_0 = x329_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@32695.4]
  assign io_sigsOut_smCtrCopyDone_1 = x338_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@32927.4]
  assign io_sigsOut_smCtrCopyDone_2 = x342_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@33142.4]
  assign x329_inr_UnitPipe_sm_clock = clock; // @[:@32602.4]
  assign x329_inr_UnitPipe_sm_reset = reset; // @[:@32603.4]
  assign x329_inr_UnitPipe_sm_io_enable = _T_375 & _T_384; // @[SpatialBlocks.scala 140:18:@32678.4]
  assign x329_inr_UnitPipe_sm_io_ctrDone = x329_inr_UnitPipe_sm_io_ctrInc & _T_362; // @[sm_x343_outr_UnitPipe.scala 77:39:@32633.4]
  assign x329_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@32680.4]
  assign x329_inr_UnitPipe_sm_io_backpressure = io_in_x322_ready | x329_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@32652.4]
  assign RetimeWrapper_clock = clock; // @[:@32659.4]
  assign RetimeWrapper_reset = reset; // @[:@32660.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@32662.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@32661.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32667.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32668.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@32670.4]
  assign RetimeWrapper_1_io_in = x329_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@32669.4]
  assign x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_in_x182_outdram_number = io_in_x182_outdram_number; // @[sm_x329_inr_UnitPipe.scala 49:31:@32732.4]
  assign x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x322_ready | x329_inr_UnitPipe_sm_io_doneLatch; // @[sm_x329_inr_UnitPipe.scala 74:22:@32751.4]
  assign x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x329_inr_UnitPipe_sm_io_datapathEn; // @[sm_x329_inr_UnitPipe.scala 74:22:@32749.4]
  assign x329_inr_UnitPipe_kernelx329_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x329_inr_UnitPipe.scala 73:18:@32737.4]
  assign x331_ctrchain_clock = clock; // @[:@32765.4]
  assign x331_ctrchain_reset = reset; // @[:@32766.4]
  assign x331_ctrchain_io_input_reset = x338_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@32926.4]
  assign x331_ctrchain_io_input_enable = x338_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@32878.4 SpatialBlocks.scala 159:42:@32925.4]
  assign x338_inr_Foreach_sm_clock = clock; // @[:@32818.4]
  assign x338_inr_Foreach_sm_reset = reset; // @[:@32819.4]
  assign x338_inr_Foreach_sm_io_enable = _T_468 & _T_477; // @[SpatialBlocks.scala 140:18:@32905.4]
  assign x338_inr_Foreach_sm_io_ctrDone = io_rr ? _T_454 : 1'h0; // @[sm_x343_outr_UnitPipe.scala 90:38:@32853.4]
  assign x338_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@32907.4]
  assign x338_inr_Foreach_sm_io_backpressure = io_in_x323_ready | x338_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@32879.4]
  assign x338_inr_Foreach_sm_io_break = 1'h0; // @[sm_x343_outr_UnitPipe.scala 94:36:@32859.4]
  assign RetimeWrapper_2_clock = clock; // @[:@32846.4]
  assign RetimeWrapper_2_reset = reset; // @[:@32847.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@32849.4]
  assign RetimeWrapper_2_io_in = x331_ctrchain_io_output_done; // @[package.scala 94:16:@32848.4]
  assign RetimeWrapper_3_clock = clock; // @[:@32886.4]
  assign RetimeWrapper_3_reset = reset; // @[:@32887.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@32889.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@32888.4]
  assign RetimeWrapper_4_clock = clock; // @[:@32894.4]
  assign RetimeWrapper_4_reset = reset; // @[:@32895.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@32897.4]
  assign RetimeWrapper_4_io_in = x338_inr_Foreach_sm_io_done; // @[package.scala 94:16:@32896.4]
  assign x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_clock = clock; // @[:@32929.4]
  assign x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_reset = reset; // @[:@32930.4]
  assign x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_in_x186_outbuf_0_rPort_0_output_0 = io_in_x186_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@32980.4]
  assign x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x323_ready | x338_inr_Foreach_sm_io_doneLatch; // @[sm_x338_inr_Foreach.scala 83:22:@32999.4]
  assign x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_479 & _T_480; // @[sm_x338_inr_Foreach.scala 83:22:@32997.4]
  assign x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_sigsIn_break = x338_inr_Foreach_sm_io_break; // @[sm_x338_inr_Foreach.scala 83:22:@32995.4]
  assign x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{9{x331_ctrchain_io_output_counts_0[22]}},x331_ctrchain_io_output_counts_0}; // @[sm_x338_inr_Foreach.scala 83:22:@32990.4]
  assign x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x331_ctrchain_io_output_oobs_0; // @[sm_x338_inr_Foreach.scala 83:22:@32989.4]
  assign x338_inr_Foreach_kernelx338_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x338_inr_Foreach.scala 82:18:@32985.4]
  assign x342_inr_UnitPipe_sm_clock = clock; // @[:@33049.4]
  assign x342_inr_UnitPipe_sm_reset = reset; // @[:@33050.4]
  assign x342_inr_UnitPipe_sm_io_enable = x342_inr_UnitPipe_sigsIn_baseEn & x342_inr_UnitPipe_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@33125.4]
  assign x342_inr_UnitPipe_sm_io_ctrDone = x342_inr_UnitPipe_sm_io_ctrInc & _T_550; // @[sm_x343_outr_UnitPipe.scala 99:39:@33080.4]
  assign x342_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 142:21:@33127.4]
  assign RetimeWrapper_5_clock = clock; // @[:@33106.4]
  assign RetimeWrapper_5_reset = reset; // @[:@33107.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@33109.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@33108.4]
  assign RetimeWrapper_6_clock = clock; // @[:@33114.4]
  assign RetimeWrapper_6_reset = reset; // @[:@33115.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@33117.4]
  assign RetimeWrapper_6_io_in = x342_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@33116.4]
  assign x342_inr_UnitPipe_kernelx342_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x342_inr_UnitPipe_sm_io_datapathEn; // @[sm_x342_inr_UnitPipe.scala 65:22:@33192.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_362 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_550 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_362 <= 1'h0;
    end else begin
      _T_362 <= _T_359;
    end
    if (reset) begin
      _T_550 <= 1'h0;
    end else begin
      _T_550 <= _T_547;
    end
  end
endmodule
module x455_kernelx455_concrete1( // @[:@33208.2]
  input          clock, // @[:@33209.4]
  input          reset, // @[:@33210.4]
  output         io_in_x185_TVALID, // @[:@33211.4]
  input          io_in_x185_TREADY, // @[:@33211.4]
  output [255:0] io_in_x185_TDATA, // @[:@33211.4]
  input          io_in_x184_TVALID, // @[:@33211.4]
  output         io_in_x184_TREADY, // @[:@33211.4]
  input  [255:0] io_in_x184_TDATA, // @[:@33211.4]
  input  [7:0]   io_in_x184_TID, // @[:@33211.4]
  input  [7:0]   io_in_x184_TDEST, // @[:@33211.4]
  output         io_in_x324_ready, // @[:@33211.4]
  input          io_in_x324_valid, // @[:@33211.4]
  input          io_in_x323_ready, // @[:@33211.4]
  output         io_in_x323_valid, // @[:@33211.4]
  output [31:0]  io_in_x323_bits_wdata_0, // @[:@33211.4]
  output         io_in_x323_bits_wstrb, // @[:@33211.4]
  input  [63:0]  io_in_x182_outdram_number, // @[:@33211.4]
  output [20:0]  io_in_x186_outbuf_0_rPort_0_ofs_0, // @[:@33211.4]
  output         io_in_x186_outbuf_0_rPort_0_en_0, // @[:@33211.4]
  output         io_in_x186_outbuf_0_rPort_0_backpressure, // @[:@33211.4]
  input  [31:0]  io_in_x186_outbuf_0_rPort_0_output_0, // @[:@33211.4]
  input          io_in_x322_ready, // @[:@33211.4]
  output         io_in_x322_valid, // @[:@33211.4]
  output [63:0]  io_in_x322_bits_addr, // @[:@33211.4]
  output [31:0]  io_in_x322_bits_size, // @[:@33211.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@33211.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@33211.4]
  input          io_sigsIn_smChildAcks_0, // @[:@33211.4]
  input          io_sigsIn_smChildAcks_1, // @[:@33211.4]
  output         io_sigsOut_smDoneIn_0, // @[:@33211.4]
  output         io_sigsOut_smDoneIn_1, // @[:@33211.4]
  input          io_rr // @[:@33211.4]
);
  wire  x321_outr_UnitPipe_sm_clock; // @[sm_x321_outr_UnitPipe.scala 32:18:@33284.4]
  wire  x321_outr_UnitPipe_sm_reset; // @[sm_x321_outr_UnitPipe.scala 32:18:@33284.4]
  wire  x321_outr_UnitPipe_sm_io_enable; // @[sm_x321_outr_UnitPipe.scala 32:18:@33284.4]
  wire  x321_outr_UnitPipe_sm_io_done; // @[sm_x321_outr_UnitPipe.scala 32:18:@33284.4]
  wire  x321_outr_UnitPipe_sm_io_parentAck; // @[sm_x321_outr_UnitPipe.scala 32:18:@33284.4]
  wire  x321_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x321_outr_UnitPipe.scala 32:18:@33284.4]
  wire  x321_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x321_outr_UnitPipe.scala 32:18:@33284.4]
  wire  x321_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x321_outr_UnitPipe.scala 32:18:@33284.4]
  wire  x321_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x321_outr_UnitPipe.scala 32:18:@33284.4]
  wire  x321_outr_UnitPipe_sm_io_childAck_0; // @[sm_x321_outr_UnitPipe.scala 32:18:@33284.4]
  wire  x321_outr_UnitPipe_sm_io_childAck_1; // @[sm_x321_outr_UnitPipe.scala 32:18:@33284.4]
  wire  x321_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x321_outr_UnitPipe.scala 32:18:@33284.4]
  wire  x321_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x321_outr_UnitPipe.scala 32:18:@33284.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@33346.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@33346.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@33346.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@33346.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@33346.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@33354.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@33354.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@33354.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@33354.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@33354.4]
  wire  x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_clock; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire  x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_reset; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire  x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x185_TVALID; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire  x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x185_TREADY; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire [255:0] x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x185_TDATA; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire  x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x184_TVALID; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire  x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x184_TREADY; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire [255:0] x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x184_TDATA; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire [7:0] x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x184_TID; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire [7:0] x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x184_TDEST; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire  x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire  x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire  x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire  x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire  x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire  x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire  x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire  x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire  x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_rr; // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
  wire  x343_outr_UnitPipe_sm_clock; // @[sm_x343_outr_UnitPipe.scala 36:18:@33563.4]
  wire  x343_outr_UnitPipe_sm_reset; // @[sm_x343_outr_UnitPipe.scala 36:18:@33563.4]
  wire  x343_outr_UnitPipe_sm_io_enable; // @[sm_x343_outr_UnitPipe.scala 36:18:@33563.4]
  wire  x343_outr_UnitPipe_sm_io_done; // @[sm_x343_outr_UnitPipe.scala 36:18:@33563.4]
  wire  x343_outr_UnitPipe_sm_io_parentAck; // @[sm_x343_outr_UnitPipe.scala 36:18:@33563.4]
  wire  x343_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x343_outr_UnitPipe.scala 36:18:@33563.4]
  wire  x343_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x343_outr_UnitPipe.scala 36:18:@33563.4]
  wire  x343_outr_UnitPipe_sm_io_doneIn_2; // @[sm_x343_outr_UnitPipe.scala 36:18:@33563.4]
  wire  x343_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x343_outr_UnitPipe.scala 36:18:@33563.4]
  wire  x343_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x343_outr_UnitPipe.scala 36:18:@33563.4]
  wire  x343_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x343_outr_UnitPipe.scala 36:18:@33563.4]
  wire  x343_outr_UnitPipe_sm_io_childAck_0; // @[sm_x343_outr_UnitPipe.scala 36:18:@33563.4]
  wire  x343_outr_UnitPipe_sm_io_childAck_1; // @[sm_x343_outr_UnitPipe.scala 36:18:@33563.4]
  wire  x343_outr_UnitPipe_sm_io_childAck_2; // @[sm_x343_outr_UnitPipe.scala 36:18:@33563.4]
  wire  x343_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x343_outr_UnitPipe.scala 36:18:@33563.4]
  wire  x343_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x343_outr_UnitPipe.scala 36:18:@33563.4]
  wire  x343_outr_UnitPipe_sm_io_ctrCopyDone_2; // @[sm_x343_outr_UnitPipe.scala 36:18:@33563.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@33635.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@33635.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@33635.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@33635.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@33635.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@33643.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@33643.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@33643.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@33643.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@33643.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_clock; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_reset; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x324_ready; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x324_valid; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x323_ready; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x323_valid; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire [31:0] x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x323_bits_wdata_0; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x323_bits_wstrb; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire [63:0] x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x182_outdram_number; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire [20:0] x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x186_outbuf_0_rPort_0_ofs_0; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x186_outbuf_0_rPort_0_en_0; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x186_outbuf_0_rPort_0_backpressure; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire [31:0] x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x186_outbuf_0_rPort_0_output_0; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x322_ready; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x322_valid; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire [63:0] x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x322_bits_addr; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire [31:0] x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x322_bits_size; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_rr; // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
  wire  _T_408; // @[package.scala 96:25:@33351.4 package.scala 96:25:@33352.4]
  wire  _T_414; // @[package.scala 96:25:@33359.4 package.scala 96:25:@33360.4]
  wire  _T_417; // @[SpatialBlocks.scala 138:93:@33362.4]
  wire  _T_508; // @[package.scala 96:25:@33640.4 package.scala 96:25:@33641.4]
  wire  _T_514; // @[package.scala 96:25:@33648.4 package.scala 96:25:@33649.4]
  wire  _T_517; // @[SpatialBlocks.scala 138:93:@33651.4]
  x321_outr_UnitPipe_sm x321_outr_UnitPipe_sm ( // @[sm_x321_outr_UnitPipe.scala 32:18:@33284.4]
    .clock(x321_outr_UnitPipe_sm_clock),
    .reset(x321_outr_UnitPipe_sm_reset),
    .io_enable(x321_outr_UnitPipe_sm_io_enable),
    .io_done(x321_outr_UnitPipe_sm_io_done),
    .io_parentAck(x321_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x321_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x321_outr_UnitPipe_sm_io_doneIn_1),
    .io_enableOut_0(x321_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x321_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x321_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x321_outr_UnitPipe_sm_io_childAck_1),
    .io_ctrCopyDone_0(x321_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x321_outr_UnitPipe_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@33346.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@33354.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1 x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1 ( // @[sm_x321_outr_UnitPipe.scala 87:24:@33385.4]
    .clock(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_clock),
    .reset(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_reset),
    .io_in_x185_TVALID(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x185_TVALID),
    .io_in_x185_TREADY(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x185_TREADY),
    .io_in_x185_TDATA(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x185_TDATA),
    .io_in_x184_TVALID(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x184_TVALID),
    .io_in_x184_TREADY(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x184_TREADY),
    .io_in_x184_TDATA(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x184_TDATA),
    .io_in_x184_TID(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x184_TID),
    .io_in_x184_TDEST(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x184_TDEST),
    .io_sigsIn_smEnableOuts_0(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_rr)
  );
  x343_outr_UnitPipe_sm x343_outr_UnitPipe_sm ( // @[sm_x343_outr_UnitPipe.scala 36:18:@33563.4]
    .clock(x343_outr_UnitPipe_sm_clock),
    .reset(x343_outr_UnitPipe_sm_reset),
    .io_enable(x343_outr_UnitPipe_sm_io_enable),
    .io_done(x343_outr_UnitPipe_sm_io_done),
    .io_parentAck(x343_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x343_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x343_outr_UnitPipe_sm_io_doneIn_1),
    .io_doneIn_2(x343_outr_UnitPipe_sm_io_doneIn_2),
    .io_enableOut_0(x343_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x343_outr_UnitPipe_sm_io_enableOut_1),
    .io_enableOut_2(x343_outr_UnitPipe_sm_io_enableOut_2),
    .io_childAck_0(x343_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x343_outr_UnitPipe_sm_io_childAck_1),
    .io_childAck_2(x343_outr_UnitPipe_sm_io_childAck_2),
    .io_ctrCopyDone_0(x343_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x343_outr_UnitPipe_sm_io_ctrCopyDone_1),
    .io_ctrCopyDone_2(x343_outr_UnitPipe_sm_io_ctrCopyDone_2)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@33635.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@33643.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1 x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1 ( // @[sm_x343_outr_UnitPipe.scala 108:24:@33675.4]
    .clock(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_clock),
    .reset(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_reset),
    .io_in_x324_ready(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x324_ready),
    .io_in_x324_valid(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x324_valid),
    .io_in_x323_ready(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x323_ready),
    .io_in_x323_valid(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x323_valid),
    .io_in_x323_bits_wdata_0(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x323_bits_wdata_0),
    .io_in_x323_bits_wstrb(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x323_bits_wstrb),
    .io_in_x182_outdram_number(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x182_outdram_number),
    .io_in_x186_outbuf_0_rPort_0_ofs_0(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x186_outbuf_0_rPort_0_ofs_0),
    .io_in_x186_outbuf_0_rPort_0_en_0(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x186_outbuf_0_rPort_0_en_0),
    .io_in_x186_outbuf_0_rPort_0_backpressure(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x186_outbuf_0_rPort_0_backpressure),
    .io_in_x186_outbuf_0_rPort_0_output_0(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x186_outbuf_0_rPort_0_output_0),
    .io_in_x322_ready(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x322_ready),
    .io_in_x322_valid(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x322_valid),
    .io_in_x322_bits_addr(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x322_bits_addr),
    .io_in_x322_bits_size(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x322_bits_size),
    .io_sigsIn_smEnableOuts_0(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smCtrCopyDone_0(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_sigsOut_smCtrCopyDone_2(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2),
    .io_rr(x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_408 = RetimeWrapper_io_out; // @[package.scala 96:25:@33351.4 package.scala 96:25:@33352.4]
  assign _T_414 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@33359.4 package.scala 96:25:@33360.4]
  assign _T_417 = ~ _T_414; // @[SpatialBlocks.scala 138:93:@33362.4]
  assign _T_508 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@33640.4 package.scala 96:25:@33641.4]
  assign _T_514 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@33648.4 package.scala 96:25:@33649.4]
  assign _T_517 = ~ _T_514; // @[SpatialBlocks.scala 138:93:@33651.4]
  assign io_in_x185_TVALID = x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x185_TVALID; // @[sm_x321_outr_UnitPipe.scala 48:23:@33454.4]
  assign io_in_x185_TDATA = x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x185_TDATA; // @[sm_x321_outr_UnitPipe.scala 48:23:@33452.4]
  assign io_in_x184_TREADY = x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x184_TREADY; // @[sm_x321_outr_UnitPipe.scala 49:23:@33462.4]
  assign io_in_x324_ready = x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x324_ready; // @[sm_x343_outr_UnitPipe.scala 58:23:@33757.4]
  assign io_in_x323_valid = x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x323_valid; // @[sm_x343_outr_UnitPipe.scala 59:23:@33760.4]
  assign io_in_x323_bits_wdata_0 = x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x323_bits_wdata_0; // @[sm_x343_outr_UnitPipe.scala 59:23:@33759.4]
  assign io_in_x323_bits_wstrb = x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x323_bits_wstrb; // @[sm_x343_outr_UnitPipe.scala 59:23:@33758.4]
  assign io_in_x186_outbuf_0_rPort_0_ofs_0 = x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x186_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@33766.4]
  assign io_in_x186_outbuf_0_rPort_0_en_0 = x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x186_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@33765.4]
  assign io_in_x186_outbuf_0_rPort_0_backpressure = x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x186_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@33764.4]
  assign io_in_x322_valid = x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x322_valid; // @[sm_x343_outr_UnitPipe.scala 62:23:@33770.4]
  assign io_in_x322_bits_addr = x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x322_bits_addr; // @[sm_x343_outr_UnitPipe.scala 62:23:@33769.4]
  assign io_in_x322_bits_size = x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x322_bits_size; // @[sm_x343_outr_UnitPipe.scala 62:23:@33768.4]
  assign io_sigsOut_smDoneIn_0 = x321_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@33369.4]
  assign io_sigsOut_smDoneIn_1 = x343_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@33658.4]
  assign x321_outr_UnitPipe_sm_clock = clock; // @[:@33285.4]
  assign x321_outr_UnitPipe_sm_reset = reset; // @[:@33286.4]
  assign x321_outr_UnitPipe_sm_io_enable = _T_408 & _T_417; // @[SpatialBlocks.scala 140:18:@33366.4]
  assign x321_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@33368.4]
  assign x321_outr_UnitPipe_sm_io_doneIn_0 = x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@33336.4]
  assign x321_outr_UnitPipe_sm_io_doneIn_1 = x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@33337.4]
  assign x321_outr_UnitPipe_sm_io_ctrCopyDone_0 = x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@33383.4]
  assign x321_outr_UnitPipe_sm_io_ctrCopyDone_1 = x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@33384.4]
  assign RetimeWrapper_clock = clock; // @[:@33347.4]
  assign RetimeWrapper_reset = reset; // @[:@33348.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@33350.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@33349.4]
  assign RetimeWrapper_1_clock = clock; // @[:@33355.4]
  assign RetimeWrapper_1_reset = reset; // @[:@33356.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@33358.4]
  assign RetimeWrapper_1_io_in = x321_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@33357.4]
  assign x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_clock = clock; // @[:@33386.4]
  assign x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_reset = reset; // @[:@33387.4]
  assign x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x185_TREADY = io_in_x185_TREADY; // @[sm_x321_outr_UnitPipe.scala 48:23:@33453.4]
  assign x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x184_TVALID = io_in_x184_TVALID; // @[sm_x321_outr_UnitPipe.scala 49:23:@33463.4]
  assign x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x184_TDATA = io_in_x184_TDATA; // @[sm_x321_outr_UnitPipe.scala 49:23:@33461.4]
  assign x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x184_TID = io_in_x184_TID; // @[sm_x321_outr_UnitPipe.scala 49:23:@33457.4]
  assign x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_in_x184_TDEST = io_in_x184_TDEST; // @[sm_x321_outr_UnitPipe.scala 49:23:@33456.4]
  assign x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x321_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x321_outr_UnitPipe.scala 92:22:@33479.4]
  assign x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x321_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x321_outr_UnitPipe.scala 92:22:@33480.4]
  assign x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x321_outr_UnitPipe_sm_io_childAck_0; // @[sm_x321_outr_UnitPipe.scala 92:22:@33475.4]
  assign x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x321_outr_UnitPipe_sm_io_childAck_1; // @[sm_x321_outr_UnitPipe.scala 92:22:@33476.4]
  assign x321_outr_UnitPipe_kernelx321_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x321_outr_UnitPipe.scala 91:18:@33464.4]
  assign x343_outr_UnitPipe_sm_clock = clock; // @[:@33564.4]
  assign x343_outr_UnitPipe_sm_reset = reset; // @[:@33565.4]
  assign x343_outr_UnitPipe_sm_io_enable = _T_508 & _T_517; // @[SpatialBlocks.scala 140:18:@33655.4]
  assign x343_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@33657.4]
  assign x343_outr_UnitPipe_sm_io_doneIn_0 = x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@33623.4]
  assign x343_outr_UnitPipe_sm_io_doneIn_1 = x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@33624.4]
  assign x343_outr_UnitPipe_sm_io_doneIn_2 = x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:67:@33625.4]
  assign x343_outr_UnitPipe_sm_io_ctrCopyDone_0 = x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@33672.4]
  assign x343_outr_UnitPipe_sm_io_ctrCopyDone_1 = x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@33673.4]
  assign x343_outr_UnitPipe_sm_io_ctrCopyDone_2 = x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[SpatialBlocks.scala 161:90:@33674.4]
  assign RetimeWrapper_2_clock = clock; // @[:@33636.4]
  assign RetimeWrapper_2_reset = reset; // @[:@33637.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@33639.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@33638.4]
  assign RetimeWrapper_3_clock = clock; // @[:@33644.4]
  assign RetimeWrapper_3_reset = reset; // @[:@33645.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@33647.4]
  assign RetimeWrapper_3_io_in = x343_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@33646.4]
  assign x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_clock = clock; // @[:@33676.4]
  assign x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_reset = reset; // @[:@33677.4]
  assign x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x324_valid = io_in_x324_valid; // @[sm_x343_outr_UnitPipe.scala 58:23:@33756.4]
  assign x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x323_ready = io_in_x323_ready; // @[sm_x343_outr_UnitPipe.scala 59:23:@33761.4]
  assign x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x182_outdram_number = io_in_x182_outdram_number; // @[sm_x343_outr_UnitPipe.scala 60:31:@33762.4]
  assign x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x186_outbuf_0_rPort_0_output_0 = io_in_x186_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@33763.4]
  assign x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_in_x322_ready = io_in_x322_ready; // @[sm_x343_outr_UnitPipe.scala 62:23:@33771.4]
  assign x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x343_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x343_outr_UnitPipe.scala 113:22:@33794.4]
  assign x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x343_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x343_outr_UnitPipe.scala 113:22:@33795.4]
  assign x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2 = x343_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x343_outr_UnitPipe.scala 113:22:@33796.4]
  assign x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x343_outr_UnitPipe_sm_io_childAck_0; // @[sm_x343_outr_UnitPipe.scala 113:22:@33788.4]
  assign x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x343_outr_UnitPipe_sm_io_childAck_1; // @[sm_x343_outr_UnitPipe.scala 113:22:@33789.4]
  assign x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2 = x343_outr_UnitPipe_sm_io_childAck_2; // @[sm_x343_outr_UnitPipe.scala 113:22:@33790.4]
  assign x343_outr_UnitPipe_kernelx343_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x343_outr_UnitPipe.scala 112:18:@33772.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@33824.2]
  input          clock, // @[:@33825.4]
  input          reset, // @[:@33826.4]
  output         io_in_x185_TVALID, // @[:@33827.4]
  input          io_in_x185_TREADY, // @[:@33827.4]
  output [255:0] io_in_x185_TDATA, // @[:@33827.4]
  input          io_in_x184_TVALID, // @[:@33827.4]
  output         io_in_x184_TREADY, // @[:@33827.4]
  input  [255:0] io_in_x184_TDATA, // @[:@33827.4]
  input  [7:0]   io_in_x184_TID, // @[:@33827.4]
  input  [7:0]   io_in_x184_TDEST, // @[:@33827.4]
  output         io_in_x324_ready, // @[:@33827.4]
  input          io_in_x324_valid, // @[:@33827.4]
  input          io_in_x323_ready, // @[:@33827.4]
  output         io_in_x323_valid, // @[:@33827.4]
  output [31:0]  io_in_x323_bits_wdata_0, // @[:@33827.4]
  output         io_in_x323_bits_wstrb, // @[:@33827.4]
  input  [63:0]  io_in_x182_outdram_number, // @[:@33827.4]
  input          io_in_x322_ready, // @[:@33827.4]
  output         io_in_x322_valid, // @[:@33827.4]
  output [63:0]  io_in_x322_bits_addr, // @[:@33827.4]
  output [31:0]  io_in_x322_bits_size, // @[:@33827.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@33827.4]
  input          io_sigsIn_smChildAcks_0, // @[:@33827.4]
  output         io_sigsOut_smDoneIn_0, // @[:@33827.4]
  input          io_rr // @[:@33827.4]
);
  wire  x186_outbuf_0_clock; // @[m_x186_outbuf_0.scala 27:17:@33837.4]
  wire  x186_outbuf_0_reset; // @[m_x186_outbuf_0.scala 27:17:@33837.4]
  wire [20:0] x186_outbuf_0_io_rPort_0_ofs_0; // @[m_x186_outbuf_0.scala 27:17:@33837.4]
  wire  x186_outbuf_0_io_rPort_0_en_0; // @[m_x186_outbuf_0.scala 27:17:@33837.4]
  wire  x186_outbuf_0_io_rPort_0_backpressure; // @[m_x186_outbuf_0.scala 27:17:@33837.4]
  wire [31:0] x186_outbuf_0_io_rPort_0_output_0; // @[m_x186_outbuf_0.scala 27:17:@33837.4]
  wire  x455_sm_clock; // @[sm_x455.scala 37:18:@33895.4]
  wire  x455_sm_reset; // @[sm_x455.scala 37:18:@33895.4]
  wire  x455_sm_io_enable; // @[sm_x455.scala 37:18:@33895.4]
  wire  x455_sm_io_done; // @[sm_x455.scala 37:18:@33895.4]
  wire  x455_sm_io_ctrDone; // @[sm_x455.scala 37:18:@33895.4]
  wire  x455_sm_io_ctrInc; // @[sm_x455.scala 37:18:@33895.4]
  wire  x455_sm_io_parentAck; // @[sm_x455.scala 37:18:@33895.4]
  wire  x455_sm_io_doneIn_0; // @[sm_x455.scala 37:18:@33895.4]
  wire  x455_sm_io_doneIn_1; // @[sm_x455.scala 37:18:@33895.4]
  wire  x455_sm_io_enableOut_0; // @[sm_x455.scala 37:18:@33895.4]
  wire  x455_sm_io_enableOut_1; // @[sm_x455.scala 37:18:@33895.4]
  wire  x455_sm_io_childAck_0; // @[sm_x455.scala 37:18:@33895.4]
  wire  x455_sm_io_childAck_1; // @[sm_x455.scala 37:18:@33895.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@33962.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@33962.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@33962.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@33962.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@33962.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@33970.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@33970.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@33970.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@33970.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@33970.4]
  wire  x455_kernelx455_concrete1_clock; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_reset; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_in_x185_TVALID; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_in_x185_TREADY; // @[sm_x455.scala 102:24:@33999.4]
  wire [255:0] x455_kernelx455_concrete1_io_in_x185_TDATA; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_in_x184_TVALID; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_in_x184_TREADY; // @[sm_x455.scala 102:24:@33999.4]
  wire [255:0] x455_kernelx455_concrete1_io_in_x184_TDATA; // @[sm_x455.scala 102:24:@33999.4]
  wire [7:0] x455_kernelx455_concrete1_io_in_x184_TID; // @[sm_x455.scala 102:24:@33999.4]
  wire [7:0] x455_kernelx455_concrete1_io_in_x184_TDEST; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_in_x324_ready; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_in_x324_valid; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_in_x323_ready; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_in_x323_valid; // @[sm_x455.scala 102:24:@33999.4]
  wire [31:0] x455_kernelx455_concrete1_io_in_x323_bits_wdata_0; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_in_x323_bits_wstrb; // @[sm_x455.scala 102:24:@33999.4]
  wire [63:0] x455_kernelx455_concrete1_io_in_x182_outdram_number; // @[sm_x455.scala 102:24:@33999.4]
  wire [20:0] x455_kernelx455_concrete1_io_in_x186_outbuf_0_rPort_0_ofs_0; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_in_x186_outbuf_0_rPort_0_en_0; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_in_x186_outbuf_0_rPort_0_backpressure; // @[sm_x455.scala 102:24:@33999.4]
  wire [31:0] x455_kernelx455_concrete1_io_in_x186_outbuf_0_rPort_0_output_0; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_in_x322_ready; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_in_x322_valid; // @[sm_x455.scala 102:24:@33999.4]
  wire [63:0] x455_kernelx455_concrete1_io_in_x322_bits_addr; // @[sm_x455.scala 102:24:@33999.4]
  wire [31:0] x455_kernelx455_concrete1_io_in_x322_bits_size; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x455.scala 102:24:@33999.4]
  wire  x455_kernelx455_concrete1_io_rr; // @[sm_x455.scala 102:24:@33999.4]
  wire  _T_266; // @[package.scala 100:49:@33928.4]
  reg  _T_269; // @[package.scala 48:56:@33929.4]
  reg [31:0] _RAND_0;
  wire  _T_283; // @[package.scala 96:25:@33967.4 package.scala 96:25:@33968.4]
  wire  _T_289; // @[package.scala 96:25:@33975.4 package.scala 96:25:@33976.4]
  wire  _T_292; // @[SpatialBlocks.scala 138:93:@33978.4]
  x186_outbuf_0 x186_outbuf_0 ( // @[m_x186_outbuf_0.scala 27:17:@33837.4]
    .clock(x186_outbuf_0_clock),
    .reset(x186_outbuf_0_reset),
    .io_rPort_0_ofs_0(x186_outbuf_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x186_outbuf_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x186_outbuf_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x186_outbuf_0_io_rPort_0_output_0)
  );
  x455_sm x455_sm ( // @[sm_x455.scala 37:18:@33895.4]
    .clock(x455_sm_clock),
    .reset(x455_sm_reset),
    .io_enable(x455_sm_io_enable),
    .io_done(x455_sm_io_done),
    .io_ctrDone(x455_sm_io_ctrDone),
    .io_ctrInc(x455_sm_io_ctrInc),
    .io_parentAck(x455_sm_io_parentAck),
    .io_doneIn_0(x455_sm_io_doneIn_0),
    .io_doneIn_1(x455_sm_io_doneIn_1),
    .io_enableOut_0(x455_sm_io_enableOut_0),
    .io_enableOut_1(x455_sm_io_enableOut_1),
    .io_childAck_0(x455_sm_io_childAck_0),
    .io_childAck_1(x455_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@33962.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@33970.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x455_kernelx455_concrete1 x455_kernelx455_concrete1 ( // @[sm_x455.scala 102:24:@33999.4]
    .clock(x455_kernelx455_concrete1_clock),
    .reset(x455_kernelx455_concrete1_reset),
    .io_in_x185_TVALID(x455_kernelx455_concrete1_io_in_x185_TVALID),
    .io_in_x185_TREADY(x455_kernelx455_concrete1_io_in_x185_TREADY),
    .io_in_x185_TDATA(x455_kernelx455_concrete1_io_in_x185_TDATA),
    .io_in_x184_TVALID(x455_kernelx455_concrete1_io_in_x184_TVALID),
    .io_in_x184_TREADY(x455_kernelx455_concrete1_io_in_x184_TREADY),
    .io_in_x184_TDATA(x455_kernelx455_concrete1_io_in_x184_TDATA),
    .io_in_x184_TID(x455_kernelx455_concrete1_io_in_x184_TID),
    .io_in_x184_TDEST(x455_kernelx455_concrete1_io_in_x184_TDEST),
    .io_in_x324_ready(x455_kernelx455_concrete1_io_in_x324_ready),
    .io_in_x324_valid(x455_kernelx455_concrete1_io_in_x324_valid),
    .io_in_x323_ready(x455_kernelx455_concrete1_io_in_x323_ready),
    .io_in_x323_valid(x455_kernelx455_concrete1_io_in_x323_valid),
    .io_in_x323_bits_wdata_0(x455_kernelx455_concrete1_io_in_x323_bits_wdata_0),
    .io_in_x323_bits_wstrb(x455_kernelx455_concrete1_io_in_x323_bits_wstrb),
    .io_in_x182_outdram_number(x455_kernelx455_concrete1_io_in_x182_outdram_number),
    .io_in_x186_outbuf_0_rPort_0_ofs_0(x455_kernelx455_concrete1_io_in_x186_outbuf_0_rPort_0_ofs_0),
    .io_in_x186_outbuf_0_rPort_0_en_0(x455_kernelx455_concrete1_io_in_x186_outbuf_0_rPort_0_en_0),
    .io_in_x186_outbuf_0_rPort_0_backpressure(x455_kernelx455_concrete1_io_in_x186_outbuf_0_rPort_0_backpressure),
    .io_in_x186_outbuf_0_rPort_0_output_0(x455_kernelx455_concrete1_io_in_x186_outbuf_0_rPort_0_output_0),
    .io_in_x322_ready(x455_kernelx455_concrete1_io_in_x322_ready),
    .io_in_x322_valid(x455_kernelx455_concrete1_io_in_x322_valid),
    .io_in_x322_bits_addr(x455_kernelx455_concrete1_io_in_x322_bits_addr),
    .io_in_x322_bits_size(x455_kernelx455_concrete1_io_in_x322_bits_size),
    .io_sigsIn_smEnableOuts_0(x455_kernelx455_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x455_kernelx455_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x455_kernelx455_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x455_kernelx455_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x455_kernelx455_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x455_kernelx455_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(x455_kernelx455_concrete1_io_rr)
  );
  assign _T_266 = x455_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@33928.4]
  assign _T_283 = RetimeWrapper_io_out; // @[package.scala 96:25:@33967.4 package.scala 96:25:@33968.4]
  assign _T_289 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@33975.4 package.scala 96:25:@33976.4]
  assign _T_292 = ~ _T_289; // @[SpatialBlocks.scala 138:93:@33978.4]
  assign io_in_x185_TVALID = x455_kernelx455_concrete1_io_in_x185_TVALID; // @[sm_x455.scala 63:23:@34086.4]
  assign io_in_x185_TDATA = x455_kernelx455_concrete1_io_in_x185_TDATA; // @[sm_x455.scala 63:23:@34084.4]
  assign io_in_x184_TREADY = x455_kernelx455_concrete1_io_in_x184_TREADY; // @[sm_x455.scala 64:23:@34094.4]
  assign io_in_x324_ready = x455_kernelx455_concrete1_io_in_x324_ready; // @[sm_x455.scala 65:23:@34098.4]
  assign io_in_x323_valid = x455_kernelx455_concrete1_io_in_x323_valid; // @[sm_x455.scala 66:23:@34101.4]
  assign io_in_x323_bits_wdata_0 = x455_kernelx455_concrete1_io_in_x323_bits_wdata_0; // @[sm_x455.scala 66:23:@34100.4]
  assign io_in_x323_bits_wstrb = x455_kernelx455_concrete1_io_in_x323_bits_wstrb; // @[sm_x455.scala 66:23:@34099.4]
  assign io_in_x322_valid = x455_kernelx455_concrete1_io_in_x322_valid; // @[sm_x455.scala 69:23:@34111.4]
  assign io_in_x322_bits_addr = x455_kernelx455_concrete1_io_in_x322_bits_addr; // @[sm_x455.scala 69:23:@34110.4]
  assign io_in_x322_bits_size = x455_kernelx455_concrete1_io_in_x322_bits_size; // @[sm_x455.scala 69:23:@34109.4]
  assign io_sigsOut_smDoneIn_0 = x455_sm_io_done; // @[SpatialBlocks.scala 156:53:@33985.4]
  assign x186_outbuf_0_clock = clock; // @[:@33838.4]
  assign x186_outbuf_0_reset = reset; // @[:@33839.4]
  assign x186_outbuf_0_io_rPort_0_ofs_0 = x455_kernelx455_concrete1_io_in_x186_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@34107.4]
  assign x186_outbuf_0_io_rPort_0_en_0 = x455_kernelx455_concrete1_io_in_x186_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@34106.4]
  assign x186_outbuf_0_io_rPort_0_backpressure = x455_kernelx455_concrete1_io_in_x186_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@34105.4]
  assign x455_sm_clock = clock; // @[:@33896.4]
  assign x455_sm_reset = reset; // @[:@33897.4]
  assign x455_sm_io_enable = _T_283 & _T_292; // @[SpatialBlocks.scala 140:18:@33982.4]
  assign x455_sm_io_ctrDone = x455_sm_io_ctrInc & _T_269; // @[sm_RootController.scala 82:26:@33932.4]
  assign x455_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@33984.4]
  assign x455_sm_io_doneIn_0 = x455_kernelx455_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@33952.4]
  assign x455_sm_io_doneIn_1 = x455_kernelx455_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@33953.4]
  assign RetimeWrapper_clock = clock; // @[:@33963.4]
  assign RetimeWrapper_reset = reset; // @[:@33964.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@33966.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@33965.4]
  assign RetimeWrapper_1_clock = clock; // @[:@33971.4]
  assign RetimeWrapper_1_reset = reset; // @[:@33972.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@33974.4]
  assign RetimeWrapper_1_io_in = x455_sm_io_done; // @[package.scala 94:16:@33973.4]
  assign x455_kernelx455_concrete1_clock = clock; // @[:@34000.4]
  assign x455_kernelx455_concrete1_reset = reset; // @[:@34001.4]
  assign x455_kernelx455_concrete1_io_in_x185_TREADY = io_in_x185_TREADY; // @[sm_x455.scala 63:23:@34085.4]
  assign x455_kernelx455_concrete1_io_in_x184_TVALID = io_in_x184_TVALID; // @[sm_x455.scala 64:23:@34095.4]
  assign x455_kernelx455_concrete1_io_in_x184_TDATA = io_in_x184_TDATA; // @[sm_x455.scala 64:23:@34093.4]
  assign x455_kernelx455_concrete1_io_in_x184_TID = io_in_x184_TID; // @[sm_x455.scala 64:23:@34089.4]
  assign x455_kernelx455_concrete1_io_in_x184_TDEST = io_in_x184_TDEST; // @[sm_x455.scala 64:23:@34088.4]
  assign x455_kernelx455_concrete1_io_in_x324_valid = io_in_x324_valid; // @[sm_x455.scala 65:23:@34097.4]
  assign x455_kernelx455_concrete1_io_in_x323_ready = io_in_x323_ready; // @[sm_x455.scala 66:23:@34102.4]
  assign x455_kernelx455_concrete1_io_in_x182_outdram_number = io_in_x182_outdram_number; // @[sm_x455.scala 67:31:@34103.4]
  assign x455_kernelx455_concrete1_io_in_x186_outbuf_0_rPort_0_output_0 = x186_outbuf_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@34104.4]
  assign x455_kernelx455_concrete1_io_in_x322_ready = io_in_x322_ready; // @[sm_x455.scala 69:23:@34112.4]
  assign x455_kernelx455_concrete1_io_sigsIn_smEnableOuts_0 = x455_sm_io_enableOut_0; // @[sm_x455.scala 107:22:@34123.4]
  assign x455_kernelx455_concrete1_io_sigsIn_smEnableOuts_1 = x455_sm_io_enableOut_1; // @[sm_x455.scala 107:22:@34124.4]
  assign x455_kernelx455_concrete1_io_sigsIn_smChildAcks_0 = x455_sm_io_childAck_0; // @[sm_x455.scala 107:22:@34119.4]
  assign x455_kernelx455_concrete1_io_sigsIn_smChildAcks_1 = x455_sm_io_childAck_1; // @[sm_x455.scala 107:22:@34120.4]
  assign x455_kernelx455_concrete1_io_rr = io_rr; // @[sm_x455.scala 106:18:@34113.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_269 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_269 <= 1'h0;
    end else begin
      _T_269 <= _T_266;
    end
  end
endmodule
module AccelUnit( // @[:@34146.2]
  input          clock, // @[:@34147.4]
  input          reset, // @[:@34148.4]
  input          io_enable, // @[:@34149.4]
  output         io_done, // @[:@34149.4]
  input          io_reset, // @[:@34149.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@34149.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@34149.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@34149.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@34149.4]
  output         io_memStreams_loads_0_data_ready, // @[:@34149.4]
  input          io_memStreams_loads_0_data_valid, // @[:@34149.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@34149.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@34149.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@34149.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@34149.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@34149.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@34149.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@34149.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@34149.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@34149.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@34149.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@34149.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@34149.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@34149.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@34149.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@34149.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@34149.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@34149.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@34149.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@34149.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@34149.4]
  input          io_memStreams_stores_0_data_ready, // @[:@34149.4]
  output         io_memStreams_stores_0_data_valid, // @[:@34149.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@34149.4]
  output         io_memStreams_stores_0_data_bits_wstrb, // @[:@34149.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@34149.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@34149.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@34149.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@34149.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@34149.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@34149.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@34149.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@34149.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@34149.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@34149.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@34149.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@34149.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@34149.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@34149.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@34149.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@34149.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@34149.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@34149.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@34149.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@34149.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@34149.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@34149.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@34149.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@34149.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@34149.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@34149.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@34149.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@34149.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@34149.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@34149.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@34149.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@34149.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@34149.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@34149.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@34149.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@34149.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@34149.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@34149.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@34149.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@34149.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@34149.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@34149.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@34149.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@34149.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@34149.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@34149.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@34149.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@34149.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@34149.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@34149.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@34149.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@34149.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@34149.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@34149.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@34149.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@34149.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@34149.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@34149.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@34149.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@34149.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@34149.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@34149.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@34149.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@34149.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@34149.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@34149.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@34149.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@34149.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@34149.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@34149.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@34149.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@34149.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@34149.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@34149.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@34149.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@34149.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@34149.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@34149.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@34149.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@34149.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@34149.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@34149.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@34149.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@34149.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@34149.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@34149.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@34149.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@34149.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@34149.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@34149.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@34149.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@34149.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@34149.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@34149.4]
  output         io_heap_0_req_valid, // @[:@34149.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@34149.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@34149.4]
  input          io_heap_0_resp_valid, // @[:@34149.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@34149.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@34149.4]
  input  [63:0]  io_argIns_0, // @[:@34149.4]
  input  [63:0]  io_argIns_1, // @[:@34149.4]
  input          io_argOuts_0_port_ready, // @[:@34149.4]
  output         io_argOuts_0_port_valid, // @[:@34149.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@34149.4]
  input  [63:0]  io_argOuts_0_echo // @[:@34149.4]
);
  wire  SingleCounter_clock; // @[Main.scala 40:32:@34297.4]
  wire  SingleCounter_reset; // @[Main.scala 40:32:@34297.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 40:32:@34297.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 40:32:@34297.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@34315.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@34315.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@34315.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@34315.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@34315.4]
  wire  SRFF_clock; // @[Main.scala 44:28:@34324.4]
  wire  SRFF_reset; // @[Main.scala 44:28:@34324.4]
  wire  SRFF_io_input_set; // @[Main.scala 44:28:@34324.4]
  wire  SRFF_io_input_reset; // @[Main.scala 44:28:@34324.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 44:28:@34324.4]
  wire  SRFF_io_output; // @[Main.scala 44:28:@34324.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 36:18:@34363.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 36:18:@34363.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 36:18:@34363.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 36:18:@34363.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 36:18:@34363.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 36:18:@34363.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 36:18:@34363.4]
  wire  RootController_sm_io_parentAck; // @[sm_RootController.scala 36:18:@34363.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 36:18:@34363.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 36:18:@34363.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 36:18:@34363.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@34395.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@34395.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@34395.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@34395.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@34395.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 91:24:@34457.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 91:24:@34457.4]
  wire  RootController_kernelRootController_concrete1_io_in_x185_TVALID; // @[sm_RootController.scala 91:24:@34457.4]
  wire  RootController_kernelRootController_concrete1_io_in_x185_TREADY; // @[sm_RootController.scala 91:24:@34457.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x185_TDATA; // @[sm_RootController.scala 91:24:@34457.4]
  wire  RootController_kernelRootController_concrete1_io_in_x184_TVALID; // @[sm_RootController.scala 91:24:@34457.4]
  wire  RootController_kernelRootController_concrete1_io_in_x184_TREADY; // @[sm_RootController.scala 91:24:@34457.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x184_TDATA; // @[sm_RootController.scala 91:24:@34457.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x184_TID; // @[sm_RootController.scala 91:24:@34457.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x184_TDEST; // @[sm_RootController.scala 91:24:@34457.4]
  wire  RootController_kernelRootController_concrete1_io_in_x324_ready; // @[sm_RootController.scala 91:24:@34457.4]
  wire  RootController_kernelRootController_concrete1_io_in_x324_valid; // @[sm_RootController.scala 91:24:@34457.4]
  wire  RootController_kernelRootController_concrete1_io_in_x323_ready; // @[sm_RootController.scala 91:24:@34457.4]
  wire  RootController_kernelRootController_concrete1_io_in_x323_valid; // @[sm_RootController.scala 91:24:@34457.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x323_bits_wdata_0; // @[sm_RootController.scala 91:24:@34457.4]
  wire  RootController_kernelRootController_concrete1_io_in_x323_bits_wstrb; // @[sm_RootController.scala 91:24:@34457.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x182_outdram_number; // @[sm_RootController.scala 91:24:@34457.4]
  wire  RootController_kernelRootController_concrete1_io_in_x322_ready; // @[sm_RootController.scala 91:24:@34457.4]
  wire  RootController_kernelRootController_concrete1_io_in_x322_valid; // @[sm_RootController.scala 91:24:@34457.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x322_bits_addr; // @[sm_RootController.scala 91:24:@34457.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x322_bits_size; // @[sm_RootController.scala 91:24:@34457.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 91:24:@34457.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 91:24:@34457.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 91:24:@34457.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 91:24:@34457.4]
  wire  _T_599; // @[package.scala 96:25:@34320.4 package.scala 96:25:@34321.4]
  wire  _T_664; // @[Main.scala 46:50:@34391.4]
  wire  _T_665; // @[Main.scala 46:59:@34392.4]
  wire  _T_677; // @[package.scala 100:49:@34412.4]
  reg  _T_680; // @[package.scala 48:56:@34413.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 40:32:@34297.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@34315.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 44:28:@34324.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 36:18:@34363.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_parentAck(RootController_sm_io_parentAck),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@34395.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 91:24:@34457.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x185_TVALID(RootController_kernelRootController_concrete1_io_in_x185_TVALID),
    .io_in_x185_TREADY(RootController_kernelRootController_concrete1_io_in_x185_TREADY),
    .io_in_x185_TDATA(RootController_kernelRootController_concrete1_io_in_x185_TDATA),
    .io_in_x184_TVALID(RootController_kernelRootController_concrete1_io_in_x184_TVALID),
    .io_in_x184_TREADY(RootController_kernelRootController_concrete1_io_in_x184_TREADY),
    .io_in_x184_TDATA(RootController_kernelRootController_concrete1_io_in_x184_TDATA),
    .io_in_x184_TID(RootController_kernelRootController_concrete1_io_in_x184_TID),
    .io_in_x184_TDEST(RootController_kernelRootController_concrete1_io_in_x184_TDEST),
    .io_in_x324_ready(RootController_kernelRootController_concrete1_io_in_x324_ready),
    .io_in_x324_valid(RootController_kernelRootController_concrete1_io_in_x324_valid),
    .io_in_x323_ready(RootController_kernelRootController_concrete1_io_in_x323_ready),
    .io_in_x323_valid(RootController_kernelRootController_concrete1_io_in_x323_valid),
    .io_in_x323_bits_wdata_0(RootController_kernelRootController_concrete1_io_in_x323_bits_wdata_0),
    .io_in_x323_bits_wstrb(RootController_kernelRootController_concrete1_io_in_x323_bits_wstrb),
    .io_in_x182_outdram_number(RootController_kernelRootController_concrete1_io_in_x182_outdram_number),
    .io_in_x322_ready(RootController_kernelRootController_concrete1_io_in_x322_ready),
    .io_in_x322_valid(RootController_kernelRootController_concrete1_io_in_x322_valid),
    .io_in_x322_bits_addr(RootController_kernelRootController_concrete1_io_in_x322_bits_addr),
    .io_in_x322_bits_size(RootController_kernelRootController_concrete1_io_in_x322_bits_size),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@34320.4 package.scala 96:25:@34321.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 46:50:@34391.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 46:59:@34392.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@34412.4]
  assign io_done = SRFF_io_output; // @[Main.scala 53:23:@34411.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x322_valid; // @[sm_RootController.scala 65:23:@34546.4]
  assign io_memStreams_stores_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x322_bits_addr; // @[sm_RootController.scala 65:23:@34545.4]
  assign io_memStreams_stores_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x322_bits_size; // @[sm_RootController.scala 65:23:@34544.4]
  assign io_memStreams_stores_0_data_valid = RootController_kernelRootController_concrete1_io_in_x323_valid; // @[sm_RootController.scala 63:23:@34541.4]
  assign io_memStreams_stores_0_data_bits_wdata_0 = RootController_kernelRootController_concrete1_io_in_x323_bits_wdata_0; // @[sm_RootController.scala 63:23:@34540.4]
  assign io_memStreams_stores_0_data_bits_wstrb = RootController_kernelRootController_concrete1_io_in_x323_bits_wstrb; // @[sm_RootController.scala 63:23:@34539.4]
  assign io_memStreams_stores_0_wresp_ready = RootController_kernelRootController_concrete1_io_in_x324_ready; // @[sm_RootController.scala 62:23:@34538.4]
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x184_TREADY; // @[sm_RootController.scala 61:23:@34534.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x185_TVALID; // @[sm_RootController.scala 60:23:@34526.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x185_TDATA; // @[sm_RootController.scala 60:23:@34524.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 60:23:@34523.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 60:23:@34522.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 60:23:@34521.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 60:23:@34520.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 60:23:@34519.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 60:23:@34518.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@34298.4]
  assign SingleCounter_reset = reset; // @[:@34299.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 41:79:@34313.4]
  assign RetimeWrapper_clock = clock; // @[:@34316.4]
  assign RetimeWrapper_reset = reset; // @[:@34317.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@34319.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@34318.4]
  assign SRFF_clock = clock; // @[:@34325.4]
  assign SRFF_reset = reset; // @[:@34326.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 62:29:@34575.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 51:31:@34409.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 52:36:@34410.4]
  assign RootController_sm_clock = clock; // @[:@34364.4]
  assign RootController_sm_reset = reset; // @[:@34365.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 50:33:@34408.4 SpatialBlocks.scala 140:18:@34442.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@34436.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 54:34:@34416.4]
  assign RootController_sm_io_parentAck = 1'h0; // @[Main.scala 49:36:@34404.4 SpatialBlocks.scala 142:21:@34444.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@34433.4]
  assign RetimeWrapper_1_clock = clock; // @[:@34396.4]
  assign RetimeWrapper_1_reset = reset; // @[:@34397.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@34399.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@34398.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@34458.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@34459.4]
  assign RootController_kernelRootController_concrete1_io_in_x185_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 60:23:@34525.4]
  assign RootController_kernelRootController_concrete1_io_in_x184_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 61:23:@34535.4]
  assign RootController_kernelRootController_concrete1_io_in_x184_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 61:23:@34533.4]
  assign RootController_kernelRootController_concrete1_io_in_x184_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 61:23:@34529.4]
  assign RootController_kernelRootController_concrete1_io_in_x184_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 61:23:@34528.4]
  assign RootController_kernelRootController_concrete1_io_in_x324_valid = io_memStreams_stores_0_wresp_valid; // @[sm_RootController.scala 62:23:@34537.4]
  assign RootController_kernelRootController_concrete1_io_in_x323_ready = io_memStreams_stores_0_data_ready; // @[sm_RootController.scala 63:23:@34542.4]
  assign RootController_kernelRootController_concrete1_io_in_x182_outdram_number = io_argIns_1; // @[sm_RootController.scala 64:31:@34543.4]
  assign RootController_kernelRootController_concrete1_io_in_x322_ready = io_memStreams_stores_0_cmd_ready; // @[sm_RootController.scala 65:23:@34547.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 96:22:@34556.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 96:22:@34554.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 95:18:@34548.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module Counter( // @[:@34577.2]
  input        clock, // @[:@34578.4]
  input        reset, // @[:@34579.4]
  input        io_enable, // @[:@34580.4]
  output [5:0] io_out, // @[:@34580.4]
  output [5:0] io_next // @[:@34580.4]
);
  reg [5:0] count; // @[Counter.scala 15:22:@34582.4]
  reg [31:0] _RAND_0;
  wire [6:0] _T_17; // @[Counter.scala 17:24:@34583.4]
  wire [5:0] newCount; // @[Counter.scala 17:24:@34584.4]
  wire [5:0] _GEN_0; // @[Counter.scala 21:26:@34589.6]
  assign _T_17 = count + 6'h1; // @[Counter.scala 17:24:@34583.4]
  assign newCount = count + 6'h1; // @[Counter.scala 17:24:@34584.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@34589.6]
  assign io_out = count; // @[Counter.scala 25:10:@34592.4]
  assign io_next = count + 6'h1; // @[Counter.scala 26:11:@34593.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 6'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module SRAM_13( // @[:@34629.2]
  input         clock, // @[:@34630.4]
  input         reset, // @[:@34631.4]
  input  [5:0]  io_raddr, // @[:@34632.4]
  input         io_wen, // @[:@34632.4]
  input  [5:0]  io_waddr, // @[:@34632.4]
  input  [63:0] io_wdata_addr, // @[:@34632.4]
  input  [31:0] io_wdata_size, // @[:@34632.4]
  output [63:0] io_rdata_addr, // @[:@34632.4]
  output [31:0] io_rdata_size // @[:@34632.4]
);
  wire [95:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@34634.4]
  wire [95:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@34634.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@34634.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@34634.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@34634.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@34634.4]
  wire [5:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@34634.4]
  wire [5:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@34634.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@34634.4]
  wire [95:0] _T_17; // @[SRAM.scala 175:38:@34648.4]
  wire  _T_20; // @[SRAM.scala 182:49:@34653.4]
  wire  _T_21; // @[SRAM.scala 182:37:@34654.4]
  reg  _T_24; // @[SRAM.scala 182:29:@34655.4]
  reg [31:0] _RAND_0;
  reg [95:0] _T_28; // @[SRAM.scala 183:29:@34658.4]
  reg [95:0] _RAND_1;
  wire [95:0] _T_29; // @[SRAM.scala 184:22:@34660.4]
  SRAMVerilogAWS #(.DWIDTH(96), .WORDS(64), .AWIDTH(6)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@34634.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_17 = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:38:@34648.4]
  assign _T_20 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@34653.4]
  assign _T_21 = io_wen & _T_20; // @[SRAM.scala 182:37:@34654.4]
  assign _T_29 = _T_24 ? _T_28 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:22:@34660.4]
  assign io_rdata_addr = _T_29[95:32]; // @[SRAM.scala 184:16:@34669.4]
  assign io_rdata_size = _T_29[31:0]; // @[SRAM.scala 184:16:@34668.4]
  assign SRAMVerilogAWS_wdata = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:20:@34649.4]
  assign SRAMVerilogAWS_backpressure = 1'h1; // @[SRAM.scala 176:27:@34650.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@34646.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@34652.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@34651.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@34647.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@34645.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@34644.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_24 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  _T_28 = _RAND_1[95:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_24 <= 1'h0;
    end else begin
      _T_24 <= _T_21;
    end
    if (reset) begin
      _T_28 <= 96'h0;
    end else begin
      _T_28 <= _T_17;
    end
  end
endmodule
module FIFO( // @[:@34671.2]
  input         clock, // @[:@34672.4]
  input         reset, // @[:@34673.4]
  output        io_in_ready, // @[:@34674.4]
  input         io_in_valid, // @[:@34674.4]
  input  [63:0] io_in_bits_addr, // @[:@34674.4]
  input  [31:0] io_in_bits_size, // @[:@34674.4]
  input         io_out_ready, // @[:@34674.4]
  output        io_out_valid, // @[:@34674.4]
  output [63:0] io_out_bits_addr, // @[:@34674.4]
  output [31:0] io_out_bits_size // @[:@34674.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@35070.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@35070.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@35070.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@35070.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@35070.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@35080.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@35080.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@35080.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@35080.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@35080.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@35095.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@35095.4]
  wire [5:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@35095.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@35095.4]
  wire [5:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@35095.4]
  wire [63:0] SRAM_io_wdata_addr; // @[FIFO.scala 73:19:@35095.4]
  wire [31:0] SRAM_io_wdata_size; // @[FIFO.scala 73:19:@35095.4]
  wire [63:0] SRAM_io_rdata_addr; // @[FIFO.scala 73:19:@35095.4]
  wire [31:0] SRAM_io_rdata_size; // @[FIFO.scala 73:19:@35095.4]
  wire  writeEn; // @[FIFO.scala 30:29:@35068.4]
  wire  readEn; // @[FIFO.scala 31:29:@35069.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@35090.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@35091.4]
  wire  _T_824; // @[FIFO.scala 45:27:@35092.4]
  wire  empty; // @[FIFO.scala 45:24:@35093.4]
  wire  full; // @[FIFO.scala 46:23:@35094.4]
  wire  _T_827; // @[FIFO.scala 83:17:@35107.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@35108.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@35070.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@35080.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_13 SRAM ( // @[FIFO.scala 73:19:@35095.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata_addr(SRAM_io_wdata_addr),
    .io_wdata_size(SRAM_io_wdata_size),
    .io_rdata_addr(SRAM_io_rdata_addr),
    .io_rdata_size(SRAM_io_rdata_size)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@35068.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@35069.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@35091.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@35092.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@35093.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@35094.4]
  assign _T_827 = writeEn != readEn; // @[FIFO.scala 83:17:@35107.4]
  assign _GEN_0 = _T_827 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@35108.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@35114.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@35112.4]
  assign io_out_bits_addr = SRAM_io_rdata_addr; // @[FIFO.scala 79:17:@35105.4]
  assign io_out_bits_size = SRAM_io_rdata_size; // @[FIFO.scala 79:17:@35104.4]
  assign enqCounter_clock = clock; // @[:@35071.4]
  assign enqCounter_reset = reset; // @[:@35072.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@35078.4]
  assign deqCounter_clock = clock; // @[:@35081.4]
  assign deqCounter_reset = reset; // @[:@35082.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@35088.4]
  assign SRAM_clock = clock; // @[:@35096.4]
  assign SRAM_reset = reset; // @[:@35097.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@35099.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@35100.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@35101.4]
  assign SRAM_io_wdata_addr = io_in_bits_addr; // @[FIFO.scala 78:16:@35103.4]
  assign SRAM_io_wdata_size = io_in_bits_size; // @[FIFO.scala 78:16:@35102.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_827) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module Counter_2( // @[:@35116.2]
  input        clock, // @[:@35117.4]
  input        reset, // @[:@35118.4]
  input        io_enable, // @[:@35119.4]
  output [3:0] io_out // @[:@35119.4]
);
  reg [3:0] count; // @[Counter.scala 15:22:@35121.4]
  reg [31:0] _RAND_0;
  wire [4:0] _T_17; // @[Counter.scala 17:24:@35122.4]
  wire [3:0] newCount; // @[Counter.scala 17:24:@35123.4]
  wire [3:0] _GEN_0; // @[Counter.scala 21:26:@35128.6]
  assign _T_17 = count + 4'h1; // @[Counter.scala 17:24:@35122.4]
  assign newCount = count + 4'h1; // @[Counter.scala 17:24:@35123.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@35128.6]
  assign io_out = count; // @[Counter.scala 25:10:@35131.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 4'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module Counter_4( // @[:@35152.2]
  input        clock, // @[:@35153.4]
  input        reset, // @[:@35154.4]
  input        io_reset, // @[:@35155.4]
  input        io_enable, // @[:@35155.4]
  input  [1:0] io_stride, // @[:@35155.4]
  output [1:0] io_out, // @[:@35155.4]
  output [1:0] io_next // @[:@35155.4]
);
  reg [1:0] count; // @[Counter.scala 15:22:@35157.4]
  reg [31:0] _RAND_0;
  wire [2:0] _T_17; // @[Counter.scala 17:24:@35158.4]
  wire [1:0] newCount; // @[Counter.scala 17:24:@35159.4]
  wire [1:0] _GEN_0; // @[Counter.scala 21:26:@35164.6]
  wire [1:0] _GEN_1; // @[Counter.scala 19:18:@35160.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@35158.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@35159.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@35164.6]
  assign _GEN_1 = io_reset ? 2'h0 : _GEN_0; // @[Counter.scala 19:18:@35160.4]
  assign io_out = count; // @[Counter.scala 25:10:@35167.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@35168.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 2'h0;
    end else begin
      if (io_reset) begin
        count <= 2'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module SRAM_14( // @[:@35204.2]
  input         clock, // @[:@35205.4]
  input         reset, // @[:@35206.4]
  input  [1:0]  io_raddr, // @[:@35207.4]
  input         io_wen, // @[:@35207.4]
  input  [1:0]  io_waddr, // @[:@35207.4]
  input  [31:0] io_wdata, // @[:@35207.4]
  output [31:0] io_rdata, // @[:@35207.4]
  input         io_backpressure // @[:@35207.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@35209.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@35209.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@35209.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@35209.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@35209.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@35209.4]
  wire [1:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@35209.4]
  wire [1:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@35209.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@35209.4]
  wire  _T_19; // @[SRAM.scala 182:49:@35227.4]
  wire  _T_20; // @[SRAM.scala 182:37:@35228.4]
  reg  _T_23; // @[SRAM.scala 182:29:@35229.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@35231.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(4), .AWIDTH(2)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@35209.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@35227.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@35228.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@35236.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@35223.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@35224.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@35221.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@35226.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@35225.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@35222.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@35220.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@35219.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module FIFO_1( // @[:@35238.2]
  input         clock, // @[:@35239.4]
  input         reset, // @[:@35240.4]
  output        io_in_ready, // @[:@35241.4]
  input         io_in_valid, // @[:@35241.4]
  input  [31:0] io_in_bits, // @[:@35241.4]
  input         io_out_ready, // @[:@35241.4]
  output        io_out_valid, // @[:@35241.4]
  output [31:0] io_out_bits // @[:@35241.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@35267.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@35267.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@35267.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@35267.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@35267.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@35267.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@35267.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@35277.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@35277.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@35277.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@35277.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@35277.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@35277.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@35277.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@35292.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@35292.4]
  wire [1:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@35292.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@35292.4]
  wire [1:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@35292.4]
  wire [31:0] SRAM_io_wdata; // @[FIFO.scala 73:19:@35292.4]
  wire [31:0] SRAM_io_rdata; // @[FIFO.scala 73:19:@35292.4]
  wire  SRAM_io_backpressure; // @[FIFO.scala 73:19:@35292.4]
  wire  writeEn; // @[FIFO.scala 30:29:@35265.4]
  wire  readEn; // @[FIFO.scala 31:29:@35266.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@35287.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@35288.4]
  wire  _T_104; // @[FIFO.scala 45:27:@35289.4]
  wire  empty; // @[FIFO.scala 45:24:@35290.4]
  wire  full; // @[FIFO.scala 46:23:@35291.4]
  wire  _T_107; // @[FIFO.scala 83:17:@35302.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@35303.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@35267.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@35277.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_14 SRAM ( // @[FIFO.scala 73:19:@35292.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@35265.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@35266.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@35288.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@35289.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@35290.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@35291.4]
  assign _T_107 = writeEn != readEn; // @[FIFO.scala 83:17:@35302.4]
  assign _GEN_0 = _T_107 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@35303.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@35309.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@35307.4]
  assign io_out_bits = SRAM_io_rdata; // @[FIFO.scala 79:17:@35300.4]
  assign enqCounter_clock = clock; // @[:@35268.4]
  assign enqCounter_reset = reset; // @[:@35269.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@35275.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@35276.4]
  assign deqCounter_clock = clock; // @[:@35278.4]
  assign deqCounter_reset = reset; // @[:@35279.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@35285.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@35286.4]
  assign SRAM_clock = clock; // @[:@35293.4]
  assign SRAM_reset = reset; // @[:@35294.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@35296.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@35297.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@35298.4]
  assign SRAM_io_wdata = io_in_bits; // @[FIFO.scala 78:16:@35299.4]
  assign SRAM_io_backpressure = 1'h1; // @[FIFO.scala 80:23:@35301.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_107) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec( // @[:@37696.2]
  input         clock, // @[:@37697.4]
  input         reset, // @[:@37698.4]
  output        io_in_ready, // @[:@37699.4]
  input         io_in_valid, // @[:@37699.4]
  input  [31:0] io_in_bits_0, // @[:@37699.4]
  input         io_out_ready, // @[:@37699.4]
  output        io_out_valid, // @[:@37699.4]
  output [31:0] io_out_bits_0, // @[:@37699.4]
  output [31:0] io_out_bits_1, // @[:@37699.4]
  output [31:0] io_out_bits_2, // @[:@37699.4]
  output [31:0] io_out_bits_3, // @[:@37699.4]
  output [31:0] io_out_bits_4, // @[:@37699.4]
  output [31:0] io_out_bits_5, // @[:@37699.4]
  output [31:0] io_out_bits_6, // @[:@37699.4]
  output [31:0] io_out_bits_7, // @[:@37699.4]
  output [31:0] io_out_bits_8, // @[:@37699.4]
  output [31:0] io_out_bits_9, // @[:@37699.4]
  output [31:0] io_out_bits_10, // @[:@37699.4]
  output [31:0] io_out_bits_11, // @[:@37699.4]
  output [31:0] io_out_bits_12, // @[:@37699.4]
  output [31:0] io_out_bits_13, // @[:@37699.4]
  output [31:0] io_out_bits_14, // @[:@37699.4]
  output [31:0] io_out_bits_15 // @[:@37699.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@37703.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@37703.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@37703.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@37703.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@37714.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@37714.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@37714.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@37714.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@37727.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@37727.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@37727.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@37727.4]
  wire [31:0] fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@37727.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@37727.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@37727.4]
  wire [31:0] fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@37727.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@37762.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@37762.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@37762.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@37762.4]
  wire [31:0] fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@37762.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@37762.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@37762.4]
  wire [31:0] fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@37762.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@37797.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@37797.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@37797.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@37797.4]
  wire [31:0] fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@37797.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@37797.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@37797.4]
  wire [31:0] fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@37797.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@37832.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@37832.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@37832.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@37832.4]
  wire [31:0] fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@37832.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@37832.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@37832.4]
  wire [31:0] fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@37832.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@37867.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@37867.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@37867.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@37867.4]
  wire [31:0] fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@37867.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@37867.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@37867.4]
  wire [31:0] fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@37867.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@37902.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@37902.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@37902.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@37902.4]
  wire [31:0] fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@37902.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@37902.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@37902.4]
  wire [31:0] fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@37902.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@37937.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@37937.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@37937.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@37937.4]
  wire [31:0] fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@37937.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@37937.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@37937.4]
  wire [31:0] fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@37937.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@37972.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@37972.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@37972.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@37972.4]
  wire [31:0] fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@37972.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@37972.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@37972.4]
  wire [31:0] fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@37972.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@38007.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@38007.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@38007.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@38007.4]
  wire [31:0] fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@38007.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@38007.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@38007.4]
  wire [31:0] fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@38007.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@38042.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@38042.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@38042.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@38042.4]
  wire [31:0] fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@38042.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@38042.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@38042.4]
  wire [31:0] fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@38042.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@38077.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@38077.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@38077.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@38077.4]
  wire [31:0] fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@38077.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@38077.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@38077.4]
  wire [31:0] fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@38077.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@38112.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@38112.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@38112.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@38112.4]
  wire [31:0] fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@38112.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@38112.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@38112.4]
  wire [31:0] fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@38112.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@38147.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@38147.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@38147.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@38147.4]
  wire [31:0] fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@38147.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@38147.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@38147.4]
  wire [31:0] fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@38147.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@38182.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@38182.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@38182.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@38182.4]
  wire [31:0] fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@38182.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@38182.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@38182.4]
  wire [31:0] fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@38182.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@38217.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@38217.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@38217.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@38217.4]
  wire [31:0] fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@38217.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@38217.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@38217.4]
  wire [31:0] fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@38217.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@38252.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@38252.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@38252.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@38252.4]
  wire [31:0] fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@38252.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@38252.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@38252.4]
  wire [31:0] fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@38252.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@37702.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@37725.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@37752.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@37787.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@37822.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@37857.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@37892.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@37927.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@37962.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@37997.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@38032.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@38067.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@38102.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@38137.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@38172.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@38207.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@38242.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@38277.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38288.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38289.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@38319.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38290.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@38319.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38291.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@38319.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38292.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@38319.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38293.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@38319.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38294.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@38319.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38295.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@38319.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38296.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@38319.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38297.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@38319.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38298.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@38319.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38299.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@38319.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38300.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@38319.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38301.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@38319.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38302.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@38319.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38303.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@38338.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@38339.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@38340.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@38341.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@38342.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@38343.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@38344.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@38345.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@38346.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@38347.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@38348.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@38349.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@38350.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@38351.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@37703.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@37714.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_1 fifos_0 ( // @[FIFOVec.scala 40:19:@37727.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_1 fifos_1 ( // @[FIFOVec.scala 40:19:@37762.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_1 fifos_2 ( // @[FIFOVec.scala 40:19:@37797.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_1 fifos_3 ( // @[FIFOVec.scala 40:19:@37832.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_1 fifos_4 ( // @[FIFOVec.scala 40:19:@37867.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_1 fifos_5 ( // @[FIFOVec.scala 40:19:@37902.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_1 fifos_6 ( // @[FIFOVec.scala 40:19:@37937.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_1 fifos_7 ( // @[FIFOVec.scala 40:19:@37972.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_1 fifos_8 ( // @[FIFOVec.scala 40:19:@38007.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_1 fifos_9 ( // @[FIFOVec.scala 40:19:@38042.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_1 fifos_10 ( // @[FIFOVec.scala 40:19:@38077.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_1 fifos_11 ( // @[FIFOVec.scala 40:19:@38112.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_1 fifos_12 ( // @[FIFOVec.scala 40:19:@38147.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_1 fifos_13 ( // @[FIFOVec.scala 40:19:@38182.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_1 fifos_14 ( // @[FIFOVec.scala 40:19:@38217.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_1 fifos_15 ( // @[FIFOVec.scala 40:19:@38252.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@37702.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@37725.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@37752.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@37787.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@37822.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@37857.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@37892.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@37927.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@37962.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@37997.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@38032.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@38067.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@38102.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@38137.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@38172.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@38207.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@38242.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@38277.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38288.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38289.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@38319.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38290.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@38319.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38291.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@38319.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38292.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@38319.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38293.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@38319.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38294.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@38319.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38295.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@38319.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38296.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@38319.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38297.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@38319.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38298.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@38319.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38299.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@38319.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38300.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@38319.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38301.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@38319.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38302.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@38319.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@38287.4 FIFOVec.scala 49:42:@38303.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@38338.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@38339.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@38340.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@38341.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@38342.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@38343.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@38344.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@38345.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@38346.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@38347.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@38348.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@38349.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@38350.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@38351.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@38320.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@38354.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@38662.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@38663.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@38664.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@38665.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@38666.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@38667.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@38668.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@38669.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@38670.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@38671.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@38672.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@38673.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@38674.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@38675.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@38676.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@38677.4]
  assign enqCounter_clock = clock; // @[:@37704.4]
  assign enqCounter_reset = reset; // @[:@37705.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@37712.4]
  assign deqCounter_clock = clock; // @[:@37715.4]
  assign deqCounter_reset = reset; // @[:@37716.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@37723.4]
  assign fifos_0_clock = clock; // @[:@37728.4]
  assign fifos_0_reset = reset; // @[:@37729.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@37755.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37757.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37761.4]
  assign fifos_1_clock = clock; // @[:@37763.4]
  assign fifos_1_reset = reset; // @[:@37764.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@37790.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37792.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37796.4]
  assign fifos_2_clock = clock; // @[:@37798.4]
  assign fifos_2_reset = reset; // @[:@37799.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@37825.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37827.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37831.4]
  assign fifos_3_clock = clock; // @[:@37833.4]
  assign fifos_3_reset = reset; // @[:@37834.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@37860.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37862.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37866.4]
  assign fifos_4_clock = clock; // @[:@37868.4]
  assign fifos_4_reset = reset; // @[:@37869.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@37895.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37897.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37901.4]
  assign fifos_5_clock = clock; // @[:@37903.4]
  assign fifos_5_reset = reset; // @[:@37904.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@37930.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37932.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37936.4]
  assign fifos_6_clock = clock; // @[:@37938.4]
  assign fifos_6_reset = reset; // @[:@37939.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@37965.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@37967.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@37971.4]
  assign fifos_7_clock = clock; // @[:@37973.4]
  assign fifos_7_reset = reset; // @[:@37974.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@38000.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38002.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38006.4]
  assign fifos_8_clock = clock; // @[:@38008.4]
  assign fifos_8_reset = reset; // @[:@38009.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@38035.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38037.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38041.4]
  assign fifos_9_clock = clock; // @[:@38043.4]
  assign fifos_9_reset = reset; // @[:@38044.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@38070.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38072.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38076.4]
  assign fifos_10_clock = clock; // @[:@38078.4]
  assign fifos_10_reset = reset; // @[:@38079.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@38105.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38107.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38111.4]
  assign fifos_11_clock = clock; // @[:@38113.4]
  assign fifos_11_reset = reset; // @[:@38114.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@38140.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38142.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38146.4]
  assign fifos_12_clock = clock; // @[:@38148.4]
  assign fifos_12_reset = reset; // @[:@38149.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@38175.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38177.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38181.4]
  assign fifos_13_clock = clock; // @[:@38183.4]
  assign fifos_13_reset = reset; // @[:@38184.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@38210.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38212.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38216.4]
  assign fifos_14_clock = clock; // @[:@38218.4]
  assign fifos_14_reset = reset; // @[:@38219.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@38245.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38247.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38251.4]
  assign fifos_15_clock = clock; // @[:@38253.4]
  assign fifos_15_reset = reset; // @[:@38254.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@38280.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@38282.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@38286.4]
endmodule
module FFRAM( // @[:@38751.2]
  input        clock, // @[:@38752.4]
  input        reset, // @[:@38753.4]
  input  [1:0] io_raddr, // @[:@38754.4]
  input        io_wen, // @[:@38754.4]
  input  [1:0] io_waddr, // @[:@38754.4]
  input        io_wdata, // @[:@38754.4]
  output       io_rdata, // @[:@38754.4]
  input        io_banks_0_wdata_valid, // @[:@38754.4]
  input        io_banks_0_wdata_bits, // @[:@38754.4]
  input        io_banks_1_wdata_valid, // @[:@38754.4]
  input        io_banks_1_wdata_bits, // @[:@38754.4]
  input        io_banks_2_wdata_valid, // @[:@38754.4]
  input        io_banks_2_wdata_bits, // @[:@38754.4]
  input        io_banks_3_wdata_valid, // @[:@38754.4]
  input        io_banks_3_wdata_bits // @[:@38754.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@38758.4]
  reg [31:0] _RAND_0;
  wire  _T_88; // @[SRAM.scala 148:37:@38759.4]
  wire  _T_89; // @[SRAM.scala 148:25:@38760.4]
  wire  _T_90; // @[SRAM.scala 148:15:@38761.4]
  wire  _T_91; // @[SRAM.scala 149:15:@38763.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@38762.4]
  reg  regs_1; // @[SRAM.scala 145:20:@38769.4]
  reg [31:0] _RAND_1;
  wire  _T_97; // @[SRAM.scala 148:37:@38770.4]
  wire  _T_98; // @[SRAM.scala 148:25:@38771.4]
  wire  _T_99; // @[SRAM.scala 148:15:@38772.4]
  wire  _T_100; // @[SRAM.scala 149:15:@38774.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@38773.4]
  reg  regs_2; // @[SRAM.scala 145:20:@38780.4]
  reg [31:0] _RAND_2;
  wire  _T_106; // @[SRAM.scala 148:37:@38781.4]
  wire  _T_107; // @[SRAM.scala 148:25:@38782.4]
  wire  _T_108; // @[SRAM.scala 148:15:@38783.4]
  wire  _T_109; // @[SRAM.scala 149:15:@38785.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@38784.4]
  reg  regs_3; // @[SRAM.scala 145:20:@38791.4]
  reg [31:0] _RAND_3;
  wire  _T_115; // @[SRAM.scala 148:37:@38792.4]
  wire  _T_116; // @[SRAM.scala 148:25:@38793.4]
  wire  _T_117; // @[SRAM.scala 148:15:@38794.4]
  wire  _T_118; // @[SRAM.scala 149:15:@38796.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@38795.4]
  wire  _GEN_5; // @[SRAM.scala 155:12:@38805.4]
  wire  _GEN_6; // @[SRAM.scala 155:12:@38805.4]
  assign _T_88 = io_waddr == 2'h0; // @[SRAM.scala 148:37:@38759.4]
  assign _T_89 = io_wen & _T_88; // @[SRAM.scala 148:25:@38760.4]
  assign _T_90 = io_banks_0_wdata_valid | _T_89; // @[SRAM.scala 148:15:@38761.4]
  assign _T_91 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@38763.6]
  assign _GEN_0 = _T_90 ? _T_91 : regs_0; // @[SRAM.scala 148:48:@38762.4]
  assign _T_97 = io_waddr == 2'h1; // @[SRAM.scala 148:37:@38770.4]
  assign _T_98 = io_wen & _T_97; // @[SRAM.scala 148:25:@38771.4]
  assign _T_99 = io_banks_1_wdata_valid | _T_98; // @[SRAM.scala 148:15:@38772.4]
  assign _T_100 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@38774.6]
  assign _GEN_1 = _T_99 ? _T_100 : regs_1; // @[SRAM.scala 148:48:@38773.4]
  assign _T_106 = io_waddr == 2'h2; // @[SRAM.scala 148:37:@38781.4]
  assign _T_107 = io_wen & _T_106; // @[SRAM.scala 148:25:@38782.4]
  assign _T_108 = io_banks_2_wdata_valid | _T_107; // @[SRAM.scala 148:15:@38783.4]
  assign _T_109 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@38785.6]
  assign _GEN_2 = _T_108 ? _T_109 : regs_2; // @[SRAM.scala 148:48:@38784.4]
  assign _T_115 = io_waddr == 2'h3; // @[SRAM.scala 148:37:@38792.4]
  assign _T_116 = io_wen & _T_115; // @[SRAM.scala 148:25:@38793.4]
  assign _T_117 = io_banks_3_wdata_valid | _T_116; // @[SRAM.scala 148:15:@38794.4]
  assign _T_118 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@38796.6]
  assign _GEN_3 = _T_117 ? _T_118 : regs_3; // @[SRAM.scala 148:48:@38795.4]
  assign _GEN_5 = 2'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@38805.4]
  assign _GEN_6 = 2'h2 == io_raddr ? regs_2 : _GEN_5; // @[SRAM.scala 155:12:@38805.4]
  assign io_rdata = 2'h3 == io_raddr ? regs_3 : _GEN_6; // @[SRAM.scala 155:12:@38805.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_90) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_99) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_108) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_117) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_17( // @[:@38807.2]
  input   clock, // @[:@38808.4]
  input   reset, // @[:@38809.4]
  output  io_in_ready, // @[:@38810.4]
  input   io_in_valid, // @[:@38810.4]
  input   io_in_bits, // @[:@38810.4]
  input   io_out_ready, // @[:@38810.4]
  output  io_out_valid, // @[:@38810.4]
  output  io_out_bits // @[:@38810.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@38836.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@38836.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@38836.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@38836.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@38836.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@38836.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@38836.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@38846.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@38846.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@38846.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@38846.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@38846.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@38846.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@38846.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@38861.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@38861.4]
  wire [1:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@38861.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@38861.4]
  wire [1:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@38861.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@38861.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@38861.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@38861.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@38861.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@38861.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@38861.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@38861.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@38861.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@38861.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@38861.4]
  wire  writeEn; // @[FIFO.scala 30:29:@38834.4]
  wire  readEn; // @[FIFO.scala 31:29:@38835.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@38856.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@38857.4]
  wire  _T_104; // @[FIFO.scala 45:27:@38858.4]
  wire  empty; // @[FIFO.scala 45:24:@38859.4]
  wire  full; // @[FIFO.scala 46:23:@38860.4]
  wire  _T_157; // @[FIFO.scala 83:17:@38947.4]
  wire  _GEN_4; // @[FIFO.scala 83:29:@38948.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@38836.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@38846.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM FFRAM ( // @[FIFO.scala 49:19:@38861.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@38834.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@38835.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@38857.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@38858.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@38859.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@38860.4]
  assign _T_157 = writeEn != readEn; // @[FIFO.scala 83:17:@38947.4]
  assign _GEN_4 = _T_157 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@38948.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@38954.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@38952.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@38886.4]
  assign enqCounter_clock = clock; // @[:@38837.4]
  assign enqCounter_reset = reset; // @[:@38838.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@38844.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@38845.4]
  assign deqCounter_clock = clock; // @[:@38847.4]
  assign deqCounter_reset = reset; // @[:@38848.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@38854.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@38855.4]
  assign FFRAM_clock = clock; // @[:@38862.4]
  assign FFRAM_reset = reset; // @[:@38863.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@38882.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@38883.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@38884.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@38885.4]
  assign FFRAM_io_banks_0_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@38888.4]
  assign FFRAM_io_banks_0_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@38887.4]
  assign FFRAM_io_banks_1_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@38891.4]
  assign FFRAM_io_banks_1_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@38890.4]
  assign FFRAM_io_banks_2_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@38894.4]
  assign FFRAM_io_banks_2_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@38893.4]
  assign FFRAM_io_banks_3_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@38897.4]
  assign FFRAM_io_banks_3_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@38896.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_157) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec_1( // @[:@42571.2]
  input   clock, // @[:@42572.4]
  input   reset, // @[:@42573.4]
  output  io_in_ready, // @[:@42574.4]
  input   io_in_valid, // @[:@42574.4]
  input   io_in_bits_0, // @[:@42574.4]
  input   io_out_ready, // @[:@42574.4]
  output  io_out_valid, // @[:@42574.4]
  output  io_out_bits_0, // @[:@42574.4]
  output  io_out_bits_1, // @[:@42574.4]
  output  io_out_bits_2, // @[:@42574.4]
  output  io_out_bits_3, // @[:@42574.4]
  output  io_out_bits_4, // @[:@42574.4]
  output  io_out_bits_5, // @[:@42574.4]
  output  io_out_bits_6, // @[:@42574.4]
  output  io_out_bits_7, // @[:@42574.4]
  output  io_out_bits_8, // @[:@42574.4]
  output  io_out_bits_9, // @[:@42574.4]
  output  io_out_bits_10, // @[:@42574.4]
  output  io_out_bits_11, // @[:@42574.4]
  output  io_out_bits_12, // @[:@42574.4]
  output  io_out_bits_13, // @[:@42574.4]
  output  io_out_bits_14, // @[:@42574.4]
  output  io_out_bits_15 // @[:@42574.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@42578.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@42578.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@42578.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@42578.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@42589.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@42589.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@42589.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@42589.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@42602.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@42602.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@42602.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@42602.4]
  wire  fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@42602.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@42602.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@42602.4]
  wire  fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@42602.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@42637.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@42637.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@42637.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@42637.4]
  wire  fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@42637.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@42637.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@42637.4]
  wire  fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@42637.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@42672.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@42672.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@42672.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@42672.4]
  wire  fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@42672.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@42672.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@42672.4]
  wire  fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@42672.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@42707.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@42707.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@42707.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@42707.4]
  wire  fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@42707.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@42707.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@42707.4]
  wire  fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@42707.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@42742.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@42742.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@42742.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@42742.4]
  wire  fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@42742.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@42742.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@42742.4]
  wire  fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@42742.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@42777.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@42777.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@42777.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@42777.4]
  wire  fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@42777.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@42777.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@42777.4]
  wire  fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@42777.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@42812.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@42812.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@42812.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@42812.4]
  wire  fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@42812.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@42812.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@42812.4]
  wire  fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@42812.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@42847.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@42847.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@42847.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@42847.4]
  wire  fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@42847.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@42847.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@42847.4]
  wire  fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@42847.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@42882.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@42882.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@42882.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@42882.4]
  wire  fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@42882.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@42882.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@42882.4]
  wire  fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@42882.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@42917.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@42917.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@42917.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@42917.4]
  wire  fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@42917.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@42917.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@42917.4]
  wire  fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@42917.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@42952.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@42952.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@42952.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@42952.4]
  wire  fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@42952.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@42952.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@42952.4]
  wire  fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@42952.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@42987.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@42987.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@42987.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@42987.4]
  wire  fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@42987.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@42987.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@42987.4]
  wire  fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@42987.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@43022.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@43022.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@43022.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@43022.4]
  wire  fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@43022.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@43022.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@43022.4]
  wire  fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@43022.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@43057.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@43057.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@43057.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@43057.4]
  wire  fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@43057.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@43057.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@43057.4]
  wire  fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@43057.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@43092.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@43092.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@43092.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@43092.4]
  wire  fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@43092.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@43092.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@43092.4]
  wire  fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@43092.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@43127.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@43127.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@43127.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@43127.4]
  wire  fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@43127.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@43127.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@43127.4]
  wire  fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@43127.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@42577.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@42600.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@42627.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@42662.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@42697.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@42732.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@42767.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@42802.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@42837.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@42872.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@42907.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@42942.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@42977.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@43012.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@43047.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@43082.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@43117.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@43152.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43163.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43164.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@43194.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43165.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@43194.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43166.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@43194.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43167.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@43194.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43168.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@43194.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43169.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@43194.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43170.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@43194.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43171.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@43194.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43172.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@43194.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43173.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@43194.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43174.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@43194.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43175.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@43194.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43176.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@43194.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43177.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@43194.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43178.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@43213.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@43214.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@43215.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@43216.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@43217.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@43218.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@43219.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@43220.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@43221.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@43222.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@43223.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@43224.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@43225.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@43226.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@42578.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@42589.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_17 fifos_0 ( // @[FIFOVec.scala 40:19:@42602.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_17 fifos_1 ( // @[FIFOVec.scala 40:19:@42637.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_17 fifos_2 ( // @[FIFOVec.scala 40:19:@42672.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_17 fifos_3 ( // @[FIFOVec.scala 40:19:@42707.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_17 fifos_4 ( // @[FIFOVec.scala 40:19:@42742.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_17 fifos_5 ( // @[FIFOVec.scala 40:19:@42777.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_17 fifos_6 ( // @[FIFOVec.scala 40:19:@42812.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_17 fifos_7 ( // @[FIFOVec.scala 40:19:@42847.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_17 fifos_8 ( // @[FIFOVec.scala 40:19:@42882.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_17 fifos_9 ( // @[FIFOVec.scala 40:19:@42917.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_17 fifos_10 ( // @[FIFOVec.scala 40:19:@42952.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_17 fifos_11 ( // @[FIFOVec.scala 40:19:@42987.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_17 fifos_12 ( // @[FIFOVec.scala 40:19:@43022.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_17 fifos_13 ( // @[FIFOVec.scala 40:19:@43057.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_17 fifos_14 ( // @[FIFOVec.scala 40:19:@43092.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_17 fifos_15 ( // @[FIFOVec.scala 40:19:@43127.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@42577.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@42600.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@42627.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@42662.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@42697.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@42732.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@42767.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@42802.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@42837.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@42872.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@42907.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@42942.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@42977.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@43012.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@43047.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@43082.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@43117.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@43152.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43163.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43164.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@43194.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43165.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@43194.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43166.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@43194.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43167.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@43194.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43168.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@43194.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43169.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@43194.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43170.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@43194.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43171.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@43194.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43172.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@43194.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43173.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@43194.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43174.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@43194.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43175.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@43194.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43176.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@43194.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43177.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@43194.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@43162.4 FIFOVec.scala 49:42:@43178.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@43213.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@43214.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@43215.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@43216.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@43217.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@43218.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@43219.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@43220.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@43221.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@43222.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@43223.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@43224.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@43225.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@43226.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@43195.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@43229.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@43537.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@43538.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@43539.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@43540.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@43541.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@43542.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@43543.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@43544.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@43545.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@43546.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@43547.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@43548.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@43549.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@43550.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@43551.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@43552.4]
  assign enqCounter_clock = clock; // @[:@42579.4]
  assign enqCounter_reset = reset; // @[:@42580.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@42587.4]
  assign deqCounter_clock = clock; // @[:@42590.4]
  assign deqCounter_reset = reset; // @[:@42591.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@42598.4]
  assign fifos_0_clock = clock; // @[:@42603.4]
  assign fifos_0_reset = reset; // @[:@42604.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@42630.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42632.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42636.4]
  assign fifos_1_clock = clock; // @[:@42638.4]
  assign fifos_1_reset = reset; // @[:@42639.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@42665.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42667.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42671.4]
  assign fifos_2_clock = clock; // @[:@42673.4]
  assign fifos_2_reset = reset; // @[:@42674.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@42700.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42702.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42706.4]
  assign fifos_3_clock = clock; // @[:@42708.4]
  assign fifos_3_reset = reset; // @[:@42709.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@42735.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42737.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42741.4]
  assign fifos_4_clock = clock; // @[:@42743.4]
  assign fifos_4_reset = reset; // @[:@42744.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@42770.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42772.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42776.4]
  assign fifos_5_clock = clock; // @[:@42778.4]
  assign fifos_5_reset = reset; // @[:@42779.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@42805.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42807.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42811.4]
  assign fifos_6_clock = clock; // @[:@42813.4]
  assign fifos_6_reset = reset; // @[:@42814.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@42840.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42842.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42846.4]
  assign fifos_7_clock = clock; // @[:@42848.4]
  assign fifos_7_reset = reset; // @[:@42849.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@42875.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42877.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42881.4]
  assign fifos_8_clock = clock; // @[:@42883.4]
  assign fifos_8_reset = reset; // @[:@42884.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@42910.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42912.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42916.4]
  assign fifos_9_clock = clock; // @[:@42918.4]
  assign fifos_9_reset = reset; // @[:@42919.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@42945.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42947.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42951.4]
  assign fifos_10_clock = clock; // @[:@42953.4]
  assign fifos_10_reset = reset; // @[:@42954.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@42980.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@42982.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@42986.4]
  assign fifos_11_clock = clock; // @[:@42988.4]
  assign fifos_11_reset = reset; // @[:@42989.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@43015.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43017.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43021.4]
  assign fifos_12_clock = clock; // @[:@43023.4]
  assign fifos_12_reset = reset; // @[:@43024.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@43050.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43052.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43056.4]
  assign fifos_13_clock = clock; // @[:@43058.4]
  assign fifos_13_reset = reset; // @[:@43059.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@43085.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43087.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43091.4]
  assign fifos_14_clock = clock; // @[:@43093.4]
  assign fifos_14_reset = reset; // @[:@43094.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@43120.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43122.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43126.4]
  assign fifos_15_clock = clock; // @[:@43128.4]
  assign fifos_15_reset = reset; // @[:@43129.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@43155.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@43157.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@43161.4]
endmodule
module FIFOWidthConvert( // @[:@43554.2]
  input         clock, // @[:@43555.4]
  input         reset, // @[:@43556.4]
  output        io_in_ready, // @[:@43557.4]
  input         io_in_valid, // @[:@43557.4]
  input  [31:0] io_in_bits_data_0, // @[:@43557.4]
  input         io_in_bits_strobe, // @[:@43557.4]
  input         io_out_ready, // @[:@43557.4]
  output        io_out_valid, // @[:@43557.4]
  output [31:0] io_out_bits_data_0, // @[:@43557.4]
  output [31:0] io_out_bits_data_1, // @[:@43557.4]
  output [31:0] io_out_bits_data_2, // @[:@43557.4]
  output [31:0] io_out_bits_data_3, // @[:@43557.4]
  output [31:0] io_out_bits_data_4, // @[:@43557.4]
  output [31:0] io_out_bits_data_5, // @[:@43557.4]
  output [31:0] io_out_bits_data_6, // @[:@43557.4]
  output [31:0] io_out_bits_data_7, // @[:@43557.4]
  output [31:0] io_out_bits_data_8, // @[:@43557.4]
  output [31:0] io_out_bits_data_9, // @[:@43557.4]
  output [31:0] io_out_bits_data_10, // @[:@43557.4]
  output [31:0] io_out_bits_data_11, // @[:@43557.4]
  output [31:0] io_out_bits_data_12, // @[:@43557.4]
  output [31:0] io_out_bits_data_13, // @[:@43557.4]
  output [31:0] io_out_bits_data_14, // @[:@43557.4]
  output [31:0] io_out_bits_data_15, // @[:@43557.4]
  output [63:0] io_out_bits_strobe // @[:@43557.4]
);
  wire  FIFOVec_clock; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire  FIFOVec_reset; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire  FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire  FIFOVec_io_in_valid; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire [31:0] FIFOVec_io_in_bits_0; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire  FIFOVec_io_out_ready; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire  FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire [31:0] FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire [31:0] FIFOVec_io_out_bits_1; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire [31:0] FIFOVec_io_out_bits_2; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire [31:0] FIFOVec_io_out_bits_3; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire [31:0] FIFOVec_io_out_bits_4; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire [31:0] FIFOVec_io_out_bits_5; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire [31:0] FIFOVec_io_out_bits_6; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire [31:0] FIFOVec_io_out_bits_7; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire [31:0] FIFOVec_io_out_bits_8; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire [31:0] FIFOVec_io_out_bits_9; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire [31:0] FIFOVec_io_out_bits_10; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire [31:0] FIFOVec_io_out_bits_11; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire [31:0] FIFOVec_io_out_bits_12; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire [31:0] FIFOVec_io_out_bits_13; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire [31:0] FIFOVec_io_out_bits_14; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire [31:0] FIFOVec_io_out_bits_15; // @[FIFOWidthConvert.scala 61:22:@43559.4]
  wire  FIFOVec_1_clock; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_reset; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_in_ready; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_in_valid; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_in_bits_0; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_out_ready; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_out_valid; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_out_bits_0; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_out_bits_1; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_out_bits_2; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_out_bits_3; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_out_bits_4; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_out_bits_5; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_out_bits_6; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_out_bits_7; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_out_bits_8; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_out_bits_9; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_out_bits_10; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_out_bits_11; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_out_bits_12; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_out_bits_13; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_out_bits_14; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire  FIFOVec_1_io_out_bits_15; // @[FIFOWidthConvert.scala 62:26:@43600.4]
  wire [319:0] _T_55; // @[Cat.scala 30:58:@43659.4]
  wire [511:0] _T_61; // @[Cat.scala 30:58:@43665.4]
  wire [9:0] _T_108; // @[Cat.scala 30:58:@43723.4]
  wire [15:0] _T_114; // @[Cat.scala 30:58:@43729.4]
  wire  _T_115; // @[FIFOWidthConvert.scala 36:14:@43730.4]
  wire  _T_119; // @[FIFOWidthConvert.scala 36:14:@43734.4]
  wire  _T_123; // @[FIFOWidthConvert.scala 36:14:@43738.4]
  wire  _T_127; // @[FIFOWidthConvert.scala 36:14:@43742.4]
  wire  _T_131; // @[FIFOWidthConvert.scala 36:14:@43746.4]
  wire  _T_135; // @[FIFOWidthConvert.scala 36:14:@43750.4]
  wire  _T_139; // @[FIFOWidthConvert.scala 36:14:@43754.4]
  wire  _T_143; // @[FIFOWidthConvert.scala 36:14:@43758.4]
  wire  _T_147; // @[FIFOWidthConvert.scala 36:14:@43762.4]
  wire  _T_151; // @[FIFOWidthConvert.scala 36:14:@43766.4]
  wire  _T_155; // @[FIFOWidthConvert.scala 36:14:@43770.4]
  wire  _T_159; // @[FIFOWidthConvert.scala 36:14:@43774.4]
  wire  _T_163; // @[FIFOWidthConvert.scala 36:14:@43778.4]
  wire  _T_167; // @[FIFOWidthConvert.scala 36:14:@43782.4]
  wire  _T_171; // @[FIFOWidthConvert.scala 36:14:@43786.4]
  wire  _T_175; // @[FIFOWidthConvert.scala 36:14:@43790.4]
  wire [9:0] _T_257; // @[Cat.scala 30:58:@43867.4]
  wire [18:0] _T_266; // @[Cat.scala 30:58:@43876.4]
  wire [27:0] _T_275; // @[Cat.scala 30:58:@43885.4]
  wire [36:0] _T_284; // @[Cat.scala 30:58:@43894.4]
  wire [45:0] _T_293; // @[Cat.scala 30:58:@43903.4]
  wire [54:0] _T_302; // @[Cat.scala 30:58:@43912.4]
  wire [62:0] _T_310; // @[Cat.scala 30:58:@43920.4]
  FIFOVec FIFOVec ( // @[FIFOWidthConvert.scala 61:22:@43559.4]
    .clock(FIFOVec_clock),
    .reset(FIFOVec_reset),
    .io_in_ready(FIFOVec_io_in_ready),
    .io_in_valid(FIFOVec_io_in_valid),
    .io_in_bits_0(FIFOVec_io_in_bits_0),
    .io_out_ready(FIFOVec_io_out_ready),
    .io_out_valid(FIFOVec_io_out_valid),
    .io_out_bits_0(FIFOVec_io_out_bits_0),
    .io_out_bits_1(FIFOVec_io_out_bits_1),
    .io_out_bits_2(FIFOVec_io_out_bits_2),
    .io_out_bits_3(FIFOVec_io_out_bits_3),
    .io_out_bits_4(FIFOVec_io_out_bits_4),
    .io_out_bits_5(FIFOVec_io_out_bits_5),
    .io_out_bits_6(FIFOVec_io_out_bits_6),
    .io_out_bits_7(FIFOVec_io_out_bits_7),
    .io_out_bits_8(FIFOVec_io_out_bits_8),
    .io_out_bits_9(FIFOVec_io_out_bits_9),
    .io_out_bits_10(FIFOVec_io_out_bits_10),
    .io_out_bits_11(FIFOVec_io_out_bits_11),
    .io_out_bits_12(FIFOVec_io_out_bits_12),
    .io_out_bits_13(FIFOVec_io_out_bits_13),
    .io_out_bits_14(FIFOVec_io_out_bits_14),
    .io_out_bits_15(FIFOVec_io_out_bits_15)
  );
  FIFOVec_1 FIFOVec_1 ( // @[FIFOWidthConvert.scala 62:26:@43600.4]
    .clock(FIFOVec_1_clock),
    .reset(FIFOVec_1_reset),
    .io_in_ready(FIFOVec_1_io_in_ready),
    .io_in_valid(FIFOVec_1_io_in_valid),
    .io_in_bits_0(FIFOVec_1_io_in_bits_0),
    .io_out_ready(FIFOVec_1_io_out_ready),
    .io_out_valid(FIFOVec_1_io_out_valid),
    .io_out_bits_0(FIFOVec_1_io_out_bits_0),
    .io_out_bits_1(FIFOVec_1_io_out_bits_1),
    .io_out_bits_2(FIFOVec_1_io_out_bits_2),
    .io_out_bits_3(FIFOVec_1_io_out_bits_3),
    .io_out_bits_4(FIFOVec_1_io_out_bits_4),
    .io_out_bits_5(FIFOVec_1_io_out_bits_5),
    .io_out_bits_6(FIFOVec_1_io_out_bits_6),
    .io_out_bits_7(FIFOVec_1_io_out_bits_7),
    .io_out_bits_8(FIFOVec_1_io_out_bits_8),
    .io_out_bits_9(FIFOVec_1_io_out_bits_9),
    .io_out_bits_10(FIFOVec_1_io_out_bits_10),
    .io_out_bits_11(FIFOVec_1_io_out_bits_11),
    .io_out_bits_12(FIFOVec_1_io_out_bits_12),
    .io_out_bits_13(FIFOVec_1_io_out_bits_13),
    .io_out_bits_14(FIFOVec_1_io_out_bits_14),
    .io_out_bits_15(FIFOVec_1_io_out_bits_15)
  );
  assign _T_55 = {FIFOVec_io_out_bits_15,FIFOVec_io_out_bits_14,FIFOVec_io_out_bits_13,FIFOVec_io_out_bits_12,FIFOVec_io_out_bits_11,FIFOVec_io_out_bits_10,FIFOVec_io_out_bits_9,FIFOVec_io_out_bits_8,FIFOVec_io_out_bits_7,FIFOVec_io_out_bits_6}; // @[Cat.scala 30:58:@43659.4]
  assign _T_61 = {_T_55,FIFOVec_io_out_bits_5,FIFOVec_io_out_bits_4,FIFOVec_io_out_bits_3,FIFOVec_io_out_bits_2,FIFOVec_io_out_bits_1,FIFOVec_io_out_bits_0}; // @[Cat.scala 30:58:@43665.4]
  assign _T_108 = {FIFOVec_1_io_out_bits_0,FIFOVec_1_io_out_bits_1,FIFOVec_1_io_out_bits_2,FIFOVec_1_io_out_bits_3,FIFOVec_1_io_out_bits_4,FIFOVec_1_io_out_bits_5,FIFOVec_1_io_out_bits_6,FIFOVec_1_io_out_bits_7,FIFOVec_1_io_out_bits_8,FIFOVec_1_io_out_bits_9}; // @[Cat.scala 30:58:@43723.4]
  assign _T_114 = {_T_108,FIFOVec_1_io_out_bits_10,FIFOVec_1_io_out_bits_11,FIFOVec_1_io_out_bits_12,FIFOVec_1_io_out_bits_13,FIFOVec_1_io_out_bits_14,FIFOVec_1_io_out_bits_15}; // @[Cat.scala 30:58:@43729.4]
  assign _T_115 = _T_114[0]; // @[FIFOWidthConvert.scala 36:14:@43730.4]
  assign _T_119 = _T_114[1]; // @[FIFOWidthConvert.scala 36:14:@43734.4]
  assign _T_123 = _T_114[2]; // @[FIFOWidthConvert.scala 36:14:@43738.4]
  assign _T_127 = _T_114[3]; // @[FIFOWidthConvert.scala 36:14:@43742.4]
  assign _T_131 = _T_114[4]; // @[FIFOWidthConvert.scala 36:14:@43746.4]
  assign _T_135 = _T_114[5]; // @[FIFOWidthConvert.scala 36:14:@43750.4]
  assign _T_139 = _T_114[6]; // @[FIFOWidthConvert.scala 36:14:@43754.4]
  assign _T_143 = _T_114[7]; // @[FIFOWidthConvert.scala 36:14:@43758.4]
  assign _T_147 = _T_114[8]; // @[FIFOWidthConvert.scala 36:14:@43762.4]
  assign _T_151 = _T_114[9]; // @[FIFOWidthConvert.scala 36:14:@43766.4]
  assign _T_155 = _T_114[10]; // @[FIFOWidthConvert.scala 36:14:@43770.4]
  assign _T_159 = _T_114[11]; // @[FIFOWidthConvert.scala 36:14:@43774.4]
  assign _T_163 = _T_114[12]; // @[FIFOWidthConvert.scala 36:14:@43778.4]
  assign _T_167 = _T_114[13]; // @[FIFOWidthConvert.scala 36:14:@43782.4]
  assign _T_171 = _T_114[14]; // @[FIFOWidthConvert.scala 36:14:@43786.4]
  assign _T_175 = _T_114[15]; // @[FIFOWidthConvert.scala 36:14:@43790.4]
  assign _T_257 = {_T_175,_T_175,_T_175,_T_175,_T_171,_T_171,_T_171,_T_171,_T_167,_T_167}; // @[Cat.scala 30:58:@43867.4]
  assign _T_266 = {_T_257,_T_167,_T_167,_T_163,_T_163,_T_163,_T_163,_T_159,_T_159,_T_159}; // @[Cat.scala 30:58:@43876.4]
  assign _T_275 = {_T_266,_T_159,_T_155,_T_155,_T_155,_T_155,_T_151,_T_151,_T_151,_T_151}; // @[Cat.scala 30:58:@43885.4]
  assign _T_284 = {_T_275,_T_147,_T_147,_T_147,_T_147,_T_143,_T_143,_T_143,_T_143,_T_139}; // @[Cat.scala 30:58:@43894.4]
  assign _T_293 = {_T_284,_T_139,_T_139,_T_139,_T_135,_T_135,_T_135,_T_135,_T_131,_T_131}; // @[Cat.scala 30:58:@43903.4]
  assign _T_302 = {_T_293,_T_131,_T_131,_T_127,_T_127,_T_127,_T_127,_T_123,_T_123,_T_123}; // @[Cat.scala 30:58:@43912.4]
  assign _T_310 = {_T_302,_T_123,_T_119,_T_119,_T_119,_T_119,_T_115,_T_115,_T_115}; // @[Cat.scala 30:58:@43920.4]
  assign io_in_ready = FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 71:17:@43649.4]
  assign io_out_valid = FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 72:18:@43650.4]
  assign io_out_bits_data_0 = _T_61[31:0]; // @[FIFOWidthConvert.scala 73:22:@43699.4]
  assign io_out_bits_data_1 = _T_61[63:32]; // @[FIFOWidthConvert.scala 73:22:@43700.4]
  assign io_out_bits_data_2 = _T_61[95:64]; // @[FIFOWidthConvert.scala 73:22:@43701.4]
  assign io_out_bits_data_3 = _T_61[127:96]; // @[FIFOWidthConvert.scala 73:22:@43702.4]
  assign io_out_bits_data_4 = _T_61[159:128]; // @[FIFOWidthConvert.scala 73:22:@43703.4]
  assign io_out_bits_data_5 = _T_61[191:160]; // @[FIFOWidthConvert.scala 73:22:@43704.4]
  assign io_out_bits_data_6 = _T_61[223:192]; // @[FIFOWidthConvert.scala 73:22:@43705.4]
  assign io_out_bits_data_7 = _T_61[255:224]; // @[FIFOWidthConvert.scala 73:22:@43706.4]
  assign io_out_bits_data_8 = _T_61[287:256]; // @[FIFOWidthConvert.scala 73:22:@43707.4]
  assign io_out_bits_data_9 = _T_61[319:288]; // @[FIFOWidthConvert.scala 73:22:@43708.4]
  assign io_out_bits_data_10 = _T_61[351:320]; // @[FIFOWidthConvert.scala 73:22:@43709.4]
  assign io_out_bits_data_11 = _T_61[383:352]; // @[FIFOWidthConvert.scala 73:22:@43710.4]
  assign io_out_bits_data_12 = _T_61[415:384]; // @[FIFOWidthConvert.scala 73:22:@43711.4]
  assign io_out_bits_data_13 = _T_61[447:416]; // @[FIFOWidthConvert.scala 73:22:@43712.4]
  assign io_out_bits_data_14 = _T_61[479:448]; // @[FIFOWidthConvert.scala 73:22:@43713.4]
  assign io_out_bits_data_15 = _T_61[511:480]; // @[FIFOWidthConvert.scala 73:22:@43714.4]
  assign io_out_bits_strobe = {_T_310,_T_115}; // @[FIFOWidthConvert.scala 74:24:@43922.4]
  assign FIFOVec_clock = clock; // @[:@43560.4]
  assign FIFOVec_reset = reset; // @[:@43561.4]
  assign FIFOVec_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 68:22:@43646.4]
  assign FIFOVec_io_in_bits_0 = io_in_bits_data_0; // @[FIFOWidthConvert.scala 67:24:@43645.4]
  assign FIFOVec_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 75:23:@43923.4]
  assign FIFOVec_1_clock = clock; // @[:@43601.4]
  assign FIFOVec_1_reset = reset; // @[:@43602.4]
  assign FIFOVec_1_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 70:26:@43648.4]
  assign FIFOVec_1_io_in_bits_0 = io_in_bits_strobe; // @[FIFOWidthConvert.scala 69:28:@43647.4]
  assign FIFOVec_1_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 76:27:@43924.4]
endmodule
module FFRAM_16( // @[:@43962.2]
  input        clock, // @[:@43963.4]
  input        reset, // @[:@43964.4]
  input  [5:0] io_raddr, // @[:@43965.4]
  input        io_wen, // @[:@43965.4]
  input  [5:0] io_waddr, // @[:@43965.4]
  input        io_wdata, // @[:@43965.4]
  output       io_rdata, // @[:@43965.4]
  input        io_banks_0_wdata_valid, // @[:@43965.4]
  input        io_banks_0_wdata_bits, // @[:@43965.4]
  input        io_banks_1_wdata_valid, // @[:@43965.4]
  input        io_banks_1_wdata_bits, // @[:@43965.4]
  input        io_banks_2_wdata_valid, // @[:@43965.4]
  input        io_banks_2_wdata_bits, // @[:@43965.4]
  input        io_banks_3_wdata_valid, // @[:@43965.4]
  input        io_banks_3_wdata_bits, // @[:@43965.4]
  input        io_banks_4_wdata_valid, // @[:@43965.4]
  input        io_banks_4_wdata_bits, // @[:@43965.4]
  input        io_banks_5_wdata_valid, // @[:@43965.4]
  input        io_banks_5_wdata_bits, // @[:@43965.4]
  input        io_banks_6_wdata_valid, // @[:@43965.4]
  input        io_banks_6_wdata_bits, // @[:@43965.4]
  input        io_banks_7_wdata_valid, // @[:@43965.4]
  input        io_banks_7_wdata_bits, // @[:@43965.4]
  input        io_banks_8_wdata_valid, // @[:@43965.4]
  input        io_banks_8_wdata_bits, // @[:@43965.4]
  input        io_banks_9_wdata_valid, // @[:@43965.4]
  input        io_banks_9_wdata_bits, // @[:@43965.4]
  input        io_banks_10_wdata_valid, // @[:@43965.4]
  input        io_banks_10_wdata_bits, // @[:@43965.4]
  input        io_banks_11_wdata_valid, // @[:@43965.4]
  input        io_banks_11_wdata_bits, // @[:@43965.4]
  input        io_banks_12_wdata_valid, // @[:@43965.4]
  input        io_banks_12_wdata_bits, // @[:@43965.4]
  input        io_banks_13_wdata_valid, // @[:@43965.4]
  input        io_banks_13_wdata_bits, // @[:@43965.4]
  input        io_banks_14_wdata_valid, // @[:@43965.4]
  input        io_banks_14_wdata_bits, // @[:@43965.4]
  input        io_banks_15_wdata_valid, // @[:@43965.4]
  input        io_banks_15_wdata_bits, // @[:@43965.4]
  input        io_banks_16_wdata_valid, // @[:@43965.4]
  input        io_banks_16_wdata_bits, // @[:@43965.4]
  input        io_banks_17_wdata_valid, // @[:@43965.4]
  input        io_banks_17_wdata_bits, // @[:@43965.4]
  input        io_banks_18_wdata_valid, // @[:@43965.4]
  input        io_banks_18_wdata_bits, // @[:@43965.4]
  input        io_banks_19_wdata_valid, // @[:@43965.4]
  input        io_banks_19_wdata_bits, // @[:@43965.4]
  input        io_banks_20_wdata_valid, // @[:@43965.4]
  input        io_banks_20_wdata_bits, // @[:@43965.4]
  input        io_banks_21_wdata_valid, // @[:@43965.4]
  input        io_banks_21_wdata_bits, // @[:@43965.4]
  input        io_banks_22_wdata_valid, // @[:@43965.4]
  input        io_banks_22_wdata_bits, // @[:@43965.4]
  input        io_banks_23_wdata_valid, // @[:@43965.4]
  input        io_banks_23_wdata_bits, // @[:@43965.4]
  input        io_banks_24_wdata_valid, // @[:@43965.4]
  input        io_banks_24_wdata_bits, // @[:@43965.4]
  input        io_banks_25_wdata_valid, // @[:@43965.4]
  input        io_banks_25_wdata_bits, // @[:@43965.4]
  input        io_banks_26_wdata_valid, // @[:@43965.4]
  input        io_banks_26_wdata_bits, // @[:@43965.4]
  input        io_banks_27_wdata_valid, // @[:@43965.4]
  input        io_banks_27_wdata_bits, // @[:@43965.4]
  input        io_banks_28_wdata_valid, // @[:@43965.4]
  input        io_banks_28_wdata_bits, // @[:@43965.4]
  input        io_banks_29_wdata_valid, // @[:@43965.4]
  input        io_banks_29_wdata_bits, // @[:@43965.4]
  input        io_banks_30_wdata_valid, // @[:@43965.4]
  input        io_banks_30_wdata_bits, // @[:@43965.4]
  input        io_banks_31_wdata_valid, // @[:@43965.4]
  input        io_banks_31_wdata_bits, // @[:@43965.4]
  input        io_banks_32_wdata_valid, // @[:@43965.4]
  input        io_banks_32_wdata_bits, // @[:@43965.4]
  input        io_banks_33_wdata_valid, // @[:@43965.4]
  input        io_banks_33_wdata_bits, // @[:@43965.4]
  input        io_banks_34_wdata_valid, // @[:@43965.4]
  input        io_banks_34_wdata_bits, // @[:@43965.4]
  input        io_banks_35_wdata_valid, // @[:@43965.4]
  input        io_banks_35_wdata_bits, // @[:@43965.4]
  input        io_banks_36_wdata_valid, // @[:@43965.4]
  input        io_banks_36_wdata_bits, // @[:@43965.4]
  input        io_banks_37_wdata_valid, // @[:@43965.4]
  input        io_banks_37_wdata_bits, // @[:@43965.4]
  input        io_banks_38_wdata_valid, // @[:@43965.4]
  input        io_banks_38_wdata_bits, // @[:@43965.4]
  input        io_banks_39_wdata_valid, // @[:@43965.4]
  input        io_banks_39_wdata_bits, // @[:@43965.4]
  input        io_banks_40_wdata_valid, // @[:@43965.4]
  input        io_banks_40_wdata_bits, // @[:@43965.4]
  input        io_banks_41_wdata_valid, // @[:@43965.4]
  input        io_banks_41_wdata_bits, // @[:@43965.4]
  input        io_banks_42_wdata_valid, // @[:@43965.4]
  input        io_banks_42_wdata_bits, // @[:@43965.4]
  input        io_banks_43_wdata_valid, // @[:@43965.4]
  input        io_banks_43_wdata_bits, // @[:@43965.4]
  input        io_banks_44_wdata_valid, // @[:@43965.4]
  input        io_banks_44_wdata_bits, // @[:@43965.4]
  input        io_banks_45_wdata_valid, // @[:@43965.4]
  input        io_banks_45_wdata_bits, // @[:@43965.4]
  input        io_banks_46_wdata_valid, // @[:@43965.4]
  input        io_banks_46_wdata_bits, // @[:@43965.4]
  input        io_banks_47_wdata_valid, // @[:@43965.4]
  input        io_banks_47_wdata_bits, // @[:@43965.4]
  input        io_banks_48_wdata_valid, // @[:@43965.4]
  input        io_banks_48_wdata_bits, // @[:@43965.4]
  input        io_banks_49_wdata_valid, // @[:@43965.4]
  input        io_banks_49_wdata_bits, // @[:@43965.4]
  input        io_banks_50_wdata_valid, // @[:@43965.4]
  input        io_banks_50_wdata_bits, // @[:@43965.4]
  input        io_banks_51_wdata_valid, // @[:@43965.4]
  input        io_banks_51_wdata_bits, // @[:@43965.4]
  input        io_banks_52_wdata_valid, // @[:@43965.4]
  input        io_banks_52_wdata_bits, // @[:@43965.4]
  input        io_banks_53_wdata_valid, // @[:@43965.4]
  input        io_banks_53_wdata_bits, // @[:@43965.4]
  input        io_banks_54_wdata_valid, // @[:@43965.4]
  input        io_banks_54_wdata_bits, // @[:@43965.4]
  input        io_banks_55_wdata_valid, // @[:@43965.4]
  input        io_banks_55_wdata_bits, // @[:@43965.4]
  input        io_banks_56_wdata_valid, // @[:@43965.4]
  input        io_banks_56_wdata_bits, // @[:@43965.4]
  input        io_banks_57_wdata_valid, // @[:@43965.4]
  input        io_banks_57_wdata_bits, // @[:@43965.4]
  input        io_banks_58_wdata_valid, // @[:@43965.4]
  input        io_banks_58_wdata_bits, // @[:@43965.4]
  input        io_banks_59_wdata_valid, // @[:@43965.4]
  input        io_banks_59_wdata_bits, // @[:@43965.4]
  input        io_banks_60_wdata_valid, // @[:@43965.4]
  input        io_banks_60_wdata_bits, // @[:@43965.4]
  input        io_banks_61_wdata_valid, // @[:@43965.4]
  input        io_banks_61_wdata_bits, // @[:@43965.4]
  input        io_banks_62_wdata_valid, // @[:@43965.4]
  input        io_banks_62_wdata_bits, // @[:@43965.4]
  input        io_banks_63_wdata_valid, // @[:@43965.4]
  input        io_banks_63_wdata_bits // @[:@43965.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@43969.4]
  reg [31:0] _RAND_0;
  wire  _T_688; // @[SRAM.scala 148:37:@43970.4]
  wire  _T_689; // @[SRAM.scala 148:25:@43971.4]
  wire  _T_690; // @[SRAM.scala 148:15:@43972.4]
  wire  _T_691; // @[SRAM.scala 149:15:@43974.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@43973.4]
  reg  regs_1; // @[SRAM.scala 145:20:@43980.4]
  reg [31:0] _RAND_1;
  wire  _T_697; // @[SRAM.scala 148:37:@43981.4]
  wire  _T_698; // @[SRAM.scala 148:25:@43982.4]
  wire  _T_699; // @[SRAM.scala 148:15:@43983.4]
  wire  _T_700; // @[SRAM.scala 149:15:@43985.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@43984.4]
  reg  regs_2; // @[SRAM.scala 145:20:@43991.4]
  reg [31:0] _RAND_2;
  wire  _T_706; // @[SRAM.scala 148:37:@43992.4]
  wire  _T_707; // @[SRAM.scala 148:25:@43993.4]
  wire  _T_708; // @[SRAM.scala 148:15:@43994.4]
  wire  _T_709; // @[SRAM.scala 149:15:@43996.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@43995.4]
  reg  regs_3; // @[SRAM.scala 145:20:@44002.4]
  reg [31:0] _RAND_3;
  wire  _T_715; // @[SRAM.scala 148:37:@44003.4]
  wire  _T_716; // @[SRAM.scala 148:25:@44004.4]
  wire  _T_717; // @[SRAM.scala 148:15:@44005.4]
  wire  _T_718; // @[SRAM.scala 149:15:@44007.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@44006.4]
  reg  regs_4; // @[SRAM.scala 145:20:@44013.4]
  reg [31:0] _RAND_4;
  wire  _T_724; // @[SRAM.scala 148:37:@44014.4]
  wire  _T_725; // @[SRAM.scala 148:25:@44015.4]
  wire  _T_726; // @[SRAM.scala 148:15:@44016.4]
  wire  _T_727; // @[SRAM.scala 149:15:@44018.6]
  wire  _GEN_4; // @[SRAM.scala 148:48:@44017.4]
  reg  regs_5; // @[SRAM.scala 145:20:@44024.4]
  reg [31:0] _RAND_5;
  wire  _T_733; // @[SRAM.scala 148:37:@44025.4]
  wire  _T_734; // @[SRAM.scala 148:25:@44026.4]
  wire  _T_735; // @[SRAM.scala 148:15:@44027.4]
  wire  _T_736; // @[SRAM.scala 149:15:@44029.6]
  wire  _GEN_5; // @[SRAM.scala 148:48:@44028.4]
  reg  regs_6; // @[SRAM.scala 145:20:@44035.4]
  reg [31:0] _RAND_6;
  wire  _T_742; // @[SRAM.scala 148:37:@44036.4]
  wire  _T_743; // @[SRAM.scala 148:25:@44037.4]
  wire  _T_744; // @[SRAM.scala 148:15:@44038.4]
  wire  _T_745; // @[SRAM.scala 149:15:@44040.6]
  wire  _GEN_6; // @[SRAM.scala 148:48:@44039.4]
  reg  regs_7; // @[SRAM.scala 145:20:@44046.4]
  reg [31:0] _RAND_7;
  wire  _T_751; // @[SRAM.scala 148:37:@44047.4]
  wire  _T_752; // @[SRAM.scala 148:25:@44048.4]
  wire  _T_753; // @[SRAM.scala 148:15:@44049.4]
  wire  _T_754; // @[SRAM.scala 149:15:@44051.6]
  wire  _GEN_7; // @[SRAM.scala 148:48:@44050.4]
  reg  regs_8; // @[SRAM.scala 145:20:@44057.4]
  reg [31:0] _RAND_8;
  wire  _T_760; // @[SRAM.scala 148:37:@44058.4]
  wire  _T_761; // @[SRAM.scala 148:25:@44059.4]
  wire  _T_762; // @[SRAM.scala 148:15:@44060.4]
  wire  _T_763; // @[SRAM.scala 149:15:@44062.6]
  wire  _GEN_8; // @[SRAM.scala 148:48:@44061.4]
  reg  regs_9; // @[SRAM.scala 145:20:@44068.4]
  reg [31:0] _RAND_9;
  wire  _T_769; // @[SRAM.scala 148:37:@44069.4]
  wire  _T_770; // @[SRAM.scala 148:25:@44070.4]
  wire  _T_771; // @[SRAM.scala 148:15:@44071.4]
  wire  _T_772; // @[SRAM.scala 149:15:@44073.6]
  wire  _GEN_9; // @[SRAM.scala 148:48:@44072.4]
  reg  regs_10; // @[SRAM.scala 145:20:@44079.4]
  reg [31:0] _RAND_10;
  wire  _T_778; // @[SRAM.scala 148:37:@44080.4]
  wire  _T_779; // @[SRAM.scala 148:25:@44081.4]
  wire  _T_780; // @[SRAM.scala 148:15:@44082.4]
  wire  _T_781; // @[SRAM.scala 149:15:@44084.6]
  wire  _GEN_10; // @[SRAM.scala 148:48:@44083.4]
  reg  regs_11; // @[SRAM.scala 145:20:@44090.4]
  reg [31:0] _RAND_11;
  wire  _T_787; // @[SRAM.scala 148:37:@44091.4]
  wire  _T_788; // @[SRAM.scala 148:25:@44092.4]
  wire  _T_789; // @[SRAM.scala 148:15:@44093.4]
  wire  _T_790; // @[SRAM.scala 149:15:@44095.6]
  wire  _GEN_11; // @[SRAM.scala 148:48:@44094.4]
  reg  regs_12; // @[SRAM.scala 145:20:@44101.4]
  reg [31:0] _RAND_12;
  wire  _T_796; // @[SRAM.scala 148:37:@44102.4]
  wire  _T_797; // @[SRAM.scala 148:25:@44103.4]
  wire  _T_798; // @[SRAM.scala 148:15:@44104.4]
  wire  _T_799; // @[SRAM.scala 149:15:@44106.6]
  wire  _GEN_12; // @[SRAM.scala 148:48:@44105.4]
  reg  regs_13; // @[SRAM.scala 145:20:@44112.4]
  reg [31:0] _RAND_13;
  wire  _T_805; // @[SRAM.scala 148:37:@44113.4]
  wire  _T_806; // @[SRAM.scala 148:25:@44114.4]
  wire  _T_807; // @[SRAM.scala 148:15:@44115.4]
  wire  _T_808; // @[SRAM.scala 149:15:@44117.6]
  wire  _GEN_13; // @[SRAM.scala 148:48:@44116.4]
  reg  regs_14; // @[SRAM.scala 145:20:@44123.4]
  reg [31:0] _RAND_14;
  wire  _T_814; // @[SRAM.scala 148:37:@44124.4]
  wire  _T_815; // @[SRAM.scala 148:25:@44125.4]
  wire  _T_816; // @[SRAM.scala 148:15:@44126.4]
  wire  _T_817; // @[SRAM.scala 149:15:@44128.6]
  wire  _GEN_14; // @[SRAM.scala 148:48:@44127.4]
  reg  regs_15; // @[SRAM.scala 145:20:@44134.4]
  reg [31:0] _RAND_15;
  wire  _T_823; // @[SRAM.scala 148:37:@44135.4]
  wire  _T_824; // @[SRAM.scala 148:25:@44136.4]
  wire  _T_825; // @[SRAM.scala 148:15:@44137.4]
  wire  _T_826; // @[SRAM.scala 149:15:@44139.6]
  wire  _GEN_15; // @[SRAM.scala 148:48:@44138.4]
  reg  regs_16; // @[SRAM.scala 145:20:@44145.4]
  reg [31:0] _RAND_16;
  wire  _T_832; // @[SRAM.scala 148:37:@44146.4]
  wire  _T_833; // @[SRAM.scala 148:25:@44147.4]
  wire  _T_834; // @[SRAM.scala 148:15:@44148.4]
  wire  _T_835; // @[SRAM.scala 149:15:@44150.6]
  wire  _GEN_16; // @[SRAM.scala 148:48:@44149.4]
  reg  regs_17; // @[SRAM.scala 145:20:@44156.4]
  reg [31:0] _RAND_17;
  wire  _T_841; // @[SRAM.scala 148:37:@44157.4]
  wire  _T_842; // @[SRAM.scala 148:25:@44158.4]
  wire  _T_843; // @[SRAM.scala 148:15:@44159.4]
  wire  _T_844; // @[SRAM.scala 149:15:@44161.6]
  wire  _GEN_17; // @[SRAM.scala 148:48:@44160.4]
  reg  regs_18; // @[SRAM.scala 145:20:@44167.4]
  reg [31:0] _RAND_18;
  wire  _T_850; // @[SRAM.scala 148:37:@44168.4]
  wire  _T_851; // @[SRAM.scala 148:25:@44169.4]
  wire  _T_852; // @[SRAM.scala 148:15:@44170.4]
  wire  _T_853; // @[SRAM.scala 149:15:@44172.6]
  wire  _GEN_18; // @[SRAM.scala 148:48:@44171.4]
  reg  regs_19; // @[SRAM.scala 145:20:@44178.4]
  reg [31:0] _RAND_19;
  wire  _T_859; // @[SRAM.scala 148:37:@44179.4]
  wire  _T_860; // @[SRAM.scala 148:25:@44180.4]
  wire  _T_861; // @[SRAM.scala 148:15:@44181.4]
  wire  _T_862; // @[SRAM.scala 149:15:@44183.6]
  wire  _GEN_19; // @[SRAM.scala 148:48:@44182.4]
  reg  regs_20; // @[SRAM.scala 145:20:@44189.4]
  reg [31:0] _RAND_20;
  wire  _T_868; // @[SRAM.scala 148:37:@44190.4]
  wire  _T_869; // @[SRAM.scala 148:25:@44191.4]
  wire  _T_870; // @[SRAM.scala 148:15:@44192.4]
  wire  _T_871; // @[SRAM.scala 149:15:@44194.6]
  wire  _GEN_20; // @[SRAM.scala 148:48:@44193.4]
  reg  regs_21; // @[SRAM.scala 145:20:@44200.4]
  reg [31:0] _RAND_21;
  wire  _T_877; // @[SRAM.scala 148:37:@44201.4]
  wire  _T_878; // @[SRAM.scala 148:25:@44202.4]
  wire  _T_879; // @[SRAM.scala 148:15:@44203.4]
  wire  _T_880; // @[SRAM.scala 149:15:@44205.6]
  wire  _GEN_21; // @[SRAM.scala 148:48:@44204.4]
  reg  regs_22; // @[SRAM.scala 145:20:@44211.4]
  reg [31:0] _RAND_22;
  wire  _T_886; // @[SRAM.scala 148:37:@44212.4]
  wire  _T_887; // @[SRAM.scala 148:25:@44213.4]
  wire  _T_888; // @[SRAM.scala 148:15:@44214.4]
  wire  _T_889; // @[SRAM.scala 149:15:@44216.6]
  wire  _GEN_22; // @[SRAM.scala 148:48:@44215.4]
  reg  regs_23; // @[SRAM.scala 145:20:@44222.4]
  reg [31:0] _RAND_23;
  wire  _T_895; // @[SRAM.scala 148:37:@44223.4]
  wire  _T_896; // @[SRAM.scala 148:25:@44224.4]
  wire  _T_897; // @[SRAM.scala 148:15:@44225.4]
  wire  _T_898; // @[SRAM.scala 149:15:@44227.6]
  wire  _GEN_23; // @[SRAM.scala 148:48:@44226.4]
  reg  regs_24; // @[SRAM.scala 145:20:@44233.4]
  reg [31:0] _RAND_24;
  wire  _T_904; // @[SRAM.scala 148:37:@44234.4]
  wire  _T_905; // @[SRAM.scala 148:25:@44235.4]
  wire  _T_906; // @[SRAM.scala 148:15:@44236.4]
  wire  _T_907; // @[SRAM.scala 149:15:@44238.6]
  wire  _GEN_24; // @[SRAM.scala 148:48:@44237.4]
  reg  regs_25; // @[SRAM.scala 145:20:@44244.4]
  reg [31:0] _RAND_25;
  wire  _T_913; // @[SRAM.scala 148:37:@44245.4]
  wire  _T_914; // @[SRAM.scala 148:25:@44246.4]
  wire  _T_915; // @[SRAM.scala 148:15:@44247.4]
  wire  _T_916; // @[SRAM.scala 149:15:@44249.6]
  wire  _GEN_25; // @[SRAM.scala 148:48:@44248.4]
  reg  regs_26; // @[SRAM.scala 145:20:@44255.4]
  reg [31:0] _RAND_26;
  wire  _T_922; // @[SRAM.scala 148:37:@44256.4]
  wire  _T_923; // @[SRAM.scala 148:25:@44257.4]
  wire  _T_924; // @[SRAM.scala 148:15:@44258.4]
  wire  _T_925; // @[SRAM.scala 149:15:@44260.6]
  wire  _GEN_26; // @[SRAM.scala 148:48:@44259.4]
  reg  regs_27; // @[SRAM.scala 145:20:@44266.4]
  reg [31:0] _RAND_27;
  wire  _T_931; // @[SRAM.scala 148:37:@44267.4]
  wire  _T_932; // @[SRAM.scala 148:25:@44268.4]
  wire  _T_933; // @[SRAM.scala 148:15:@44269.4]
  wire  _T_934; // @[SRAM.scala 149:15:@44271.6]
  wire  _GEN_27; // @[SRAM.scala 148:48:@44270.4]
  reg  regs_28; // @[SRAM.scala 145:20:@44277.4]
  reg [31:0] _RAND_28;
  wire  _T_940; // @[SRAM.scala 148:37:@44278.4]
  wire  _T_941; // @[SRAM.scala 148:25:@44279.4]
  wire  _T_942; // @[SRAM.scala 148:15:@44280.4]
  wire  _T_943; // @[SRAM.scala 149:15:@44282.6]
  wire  _GEN_28; // @[SRAM.scala 148:48:@44281.4]
  reg  regs_29; // @[SRAM.scala 145:20:@44288.4]
  reg [31:0] _RAND_29;
  wire  _T_949; // @[SRAM.scala 148:37:@44289.4]
  wire  _T_950; // @[SRAM.scala 148:25:@44290.4]
  wire  _T_951; // @[SRAM.scala 148:15:@44291.4]
  wire  _T_952; // @[SRAM.scala 149:15:@44293.6]
  wire  _GEN_29; // @[SRAM.scala 148:48:@44292.4]
  reg  regs_30; // @[SRAM.scala 145:20:@44299.4]
  reg [31:0] _RAND_30;
  wire  _T_958; // @[SRAM.scala 148:37:@44300.4]
  wire  _T_959; // @[SRAM.scala 148:25:@44301.4]
  wire  _T_960; // @[SRAM.scala 148:15:@44302.4]
  wire  _T_961; // @[SRAM.scala 149:15:@44304.6]
  wire  _GEN_30; // @[SRAM.scala 148:48:@44303.4]
  reg  regs_31; // @[SRAM.scala 145:20:@44310.4]
  reg [31:0] _RAND_31;
  wire  _T_967; // @[SRAM.scala 148:37:@44311.4]
  wire  _T_968; // @[SRAM.scala 148:25:@44312.4]
  wire  _T_969; // @[SRAM.scala 148:15:@44313.4]
  wire  _T_970; // @[SRAM.scala 149:15:@44315.6]
  wire  _GEN_31; // @[SRAM.scala 148:48:@44314.4]
  reg  regs_32; // @[SRAM.scala 145:20:@44321.4]
  reg [31:0] _RAND_32;
  wire  _T_976; // @[SRAM.scala 148:37:@44322.4]
  wire  _T_977; // @[SRAM.scala 148:25:@44323.4]
  wire  _T_978; // @[SRAM.scala 148:15:@44324.4]
  wire  _T_979; // @[SRAM.scala 149:15:@44326.6]
  wire  _GEN_32; // @[SRAM.scala 148:48:@44325.4]
  reg  regs_33; // @[SRAM.scala 145:20:@44332.4]
  reg [31:0] _RAND_33;
  wire  _T_985; // @[SRAM.scala 148:37:@44333.4]
  wire  _T_986; // @[SRAM.scala 148:25:@44334.4]
  wire  _T_987; // @[SRAM.scala 148:15:@44335.4]
  wire  _T_988; // @[SRAM.scala 149:15:@44337.6]
  wire  _GEN_33; // @[SRAM.scala 148:48:@44336.4]
  reg  regs_34; // @[SRAM.scala 145:20:@44343.4]
  reg [31:0] _RAND_34;
  wire  _T_994; // @[SRAM.scala 148:37:@44344.4]
  wire  _T_995; // @[SRAM.scala 148:25:@44345.4]
  wire  _T_996; // @[SRAM.scala 148:15:@44346.4]
  wire  _T_997; // @[SRAM.scala 149:15:@44348.6]
  wire  _GEN_34; // @[SRAM.scala 148:48:@44347.4]
  reg  regs_35; // @[SRAM.scala 145:20:@44354.4]
  reg [31:0] _RAND_35;
  wire  _T_1003; // @[SRAM.scala 148:37:@44355.4]
  wire  _T_1004; // @[SRAM.scala 148:25:@44356.4]
  wire  _T_1005; // @[SRAM.scala 148:15:@44357.4]
  wire  _T_1006; // @[SRAM.scala 149:15:@44359.6]
  wire  _GEN_35; // @[SRAM.scala 148:48:@44358.4]
  reg  regs_36; // @[SRAM.scala 145:20:@44365.4]
  reg [31:0] _RAND_36;
  wire  _T_1012; // @[SRAM.scala 148:37:@44366.4]
  wire  _T_1013; // @[SRAM.scala 148:25:@44367.4]
  wire  _T_1014; // @[SRAM.scala 148:15:@44368.4]
  wire  _T_1015; // @[SRAM.scala 149:15:@44370.6]
  wire  _GEN_36; // @[SRAM.scala 148:48:@44369.4]
  reg  regs_37; // @[SRAM.scala 145:20:@44376.4]
  reg [31:0] _RAND_37;
  wire  _T_1021; // @[SRAM.scala 148:37:@44377.4]
  wire  _T_1022; // @[SRAM.scala 148:25:@44378.4]
  wire  _T_1023; // @[SRAM.scala 148:15:@44379.4]
  wire  _T_1024; // @[SRAM.scala 149:15:@44381.6]
  wire  _GEN_37; // @[SRAM.scala 148:48:@44380.4]
  reg  regs_38; // @[SRAM.scala 145:20:@44387.4]
  reg [31:0] _RAND_38;
  wire  _T_1030; // @[SRAM.scala 148:37:@44388.4]
  wire  _T_1031; // @[SRAM.scala 148:25:@44389.4]
  wire  _T_1032; // @[SRAM.scala 148:15:@44390.4]
  wire  _T_1033; // @[SRAM.scala 149:15:@44392.6]
  wire  _GEN_38; // @[SRAM.scala 148:48:@44391.4]
  reg  regs_39; // @[SRAM.scala 145:20:@44398.4]
  reg [31:0] _RAND_39;
  wire  _T_1039; // @[SRAM.scala 148:37:@44399.4]
  wire  _T_1040; // @[SRAM.scala 148:25:@44400.4]
  wire  _T_1041; // @[SRAM.scala 148:15:@44401.4]
  wire  _T_1042; // @[SRAM.scala 149:15:@44403.6]
  wire  _GEN_39; // @[SRAM.scala 148:48:@44402.4]
  reg  regs_40; // @[SRAM.scala 145:20:@44409.4]
  reg [31:0] _RAND_40;
  wire  _T_1048; // @[SRAM.scala 148:37:@44410.4]
  wire  _T_1049; // @[SRAM.scala 148:25:@44411.4]
  wire  _T_1050; // @[SRAM.scala 148:15:@44412.4]
  wire  _T_1051; // @[SRAM.scala 149:15:@44414.6]
  wire  _GEN_40; // @[SRAM.scala 148:48:@44413.4]
  reg  regs_41; // @[SRAM.scala 145:20:@44420.4]
  reg [31:0] _RAND_41;
  wire  _T_1057; // @[SRAM.scala 148:37:@44421.4]
  wire  _T_1058; // @[SRAM.scala 148:25:@44422.4]
  wire  _T_1059; // @[SRAM.scala 148:15:@44423.4]
  wire  _T_1060; // @[SRAM.scala 149:15:@44425.6]
  wire  _GEN_41; // @[SRAM.scala 148:48:@44424.4]
  reg  regs_42; // @[SRAM.scala 145:20:@44431.4]
  reg [31:0] _RAND_42;
  wire  _T_1066; // @[SRAM.scala 148:37:@44432.4]
  wire  _T_1067; // @[SRAM.scala 148:25:@44433.4]
  wire  _T_1068; // @[SRAM.scala 148:15:@44434.4]
  wire  _T_1069; // @[SRAM.scala 149:15:@44436.6]
  wire  _GEN_42; // @[SRAM.scala 148:48:@44435.4]
  reg  regs_43; // @[SRAM.scala 145:20:@44442.4]
  reg [31:0] _RAND_43;
  wire  _T_1075; // @[SRAM.scala 148:37:@44443.4]
  wire  _T_1076; // @[SRAM.scala 148:25:@44444.4]
  wire  _T_1077; // @[SRAM.scala 148:15:@44445.4]
  wire  _T_1078; // @[SRAM.scala 149:15:@44447.6]
  wire  _GEN_43; // @[SRAM.scala 148:48:@44446.4]
  reg  regs_44; // @[SRAM.scala 145:20:@44453.4]
  reg [31:0] _RAND_44;
  wire  _T_1084; // @[SRAM.scala 148:37:@44454.4]
  wire  _T_1085; // @[SRAM.scala 148:25:@44455.4]
  wire  _T_1086; // @[SRAM.scala 148:15:@44456.4]
  wire  _T_1087; // @[SRAM.scala 149:15:@44458.6]
  wire  _GEN_44; // @[SRAM.scala 148:48:@44457.4]
  reg  regs_45; // @[SRAM.scala 145:20:@44464.4]
  reg [31:0] _RAND_45;
  wire  _T_1093; // @[SRAM.scala 148:37:@44465.4]
  wire  _T_1094; // @[SRAM.scala 148:25:@44466.4]
  wire  _T_1095; // @[SRAM.scala 148:15:@44467.4]
  wire  _T_1096; // @[SRAM.scala 149:15:@44469.6]
  wire  _GEN_45; // @[SRAM.scala 148:48:@44468.4]
  reg  regs_46; // @[SRAM.scala 145:20:@44475.4]
  reg [31:0] _RAND_46;
  wire  _T_1102; // @[SRAM.scala 148:37:@44476.4]
  wire  _T_1103; // @[SRAM.scala 148:25:@44477.4]
  wire  _T_1104; // @[SRAM.scala 148:15:@44478.4]
  wire  _T_1105; // @[SRAM.scala 149:15:@44480.6]
  wire  _GEN_46; // @[SRAM.scala 148:48:@44479.4]
  reg  regs_47; // @[SRAM.scala 145:20:@44486.4]
  reg [31:0] _RAND_47;
  wire  _T_1111; // @[SRAM.scala 148:37:@44487.4]
  wire  _T_1112; // @[SRAM.scala 148:25:@44488.4]
  wire  _T_1113; // @[SRAM.scala 148:15:@44489.4]
  wire  _T_1114; // @[SRAM.scala 149:15:@44491.6]
  wire  _GEN_47; // @[SRAM.scala 148:48:@44490.4]
  reg  regs_48; // @[SRAM.scala 145:20:@44497.4]
  reg [31:0] _RAND_48;
  wire  _T_1120; // @[SRAM.scala 148:37:@44498.4]
  wire  _T_1121; // @[SRAM.scala 148:25:@44499.4]
  wire  _T_1122; // @[SRAM.scala 148:15:@44500.4]
  wire  _T_1123; // @[SRAM.scala 149:15:@44502.6]
  wire  _GEN_48; // @[SRAM.scala 148:48:@44501.4]
  reg  regs_49; // @[SRAM.scala 145:20:@44508.4]
  reg [31:0] _RAND_49;
  wire  _T_1129; // @[SRAM.scala 148:37:@44509.4]
  wire  _T_1130; // @[SRAM.scala 148:25:@44510.4]
  wire  _T_1131; // @[SRAM.scala 148:15:@44511.4]
  wire  _T_1132; // @[SRAM.scala 149:15:@44513.6]
  wire  _GEN_49; // @[SRAM.scala 148:48:@44512.4]
  reg  regs_50; // @[SRAM.scala 145:20:@44519.4]
  reg [31:0] _RAND_50;
  wire  _T_1138; // @[SRAM.scala 148:37:@44520.4]
  wire  _T_1139; // @[SRAM.scala 148:25:@44521.4]
  wire  _T_1140; // @[SRAM.scala 148:15:@44522.4]
  wire  _T_1141; // @[SRAM.scala 149:15:@44524.6]
  wire  _GEN_50; // @[SRAM.scala 148:48:@44523.4]
  reg  regs_51; // @[SRAM.scala 145:20:@44530.4]
  reg [31:0] _RAND_51;
  wire  _T_1147; // @[SRAM.scala 148:37:@44531.4]
  wire  _T_1148; // @[SRAM.scala 148:25:@44532.4]
  wire  _T_1149; // @[SRAM.scala 148:15:@44533.4]
  wire  _T_1150; // @[SRAM.scala 149:15:@44535.6]
  wire  _GEN_51; // @[SRAM.scala 148:48:@44534.4]
  reg  regs_52; // @[SRAM.scala 145:20:@44541.4]
  reg [31:0] _RAND_52;
  wire  _T_1156; // @[SRAM.scala 148:37:@44542.4]
  wire  _T_1157; // @[SRAM.scala 148:25:@44543.4]
  wire  _T_1158; // @[SRAM.scala 148:15:@44544.4]
  wire  _T_1159; // @[SRAM.scala 149:15:@44546.6]
  wire  _GEN_52; // @[SRAM.scala 148:48:@44545.4]
  reg  regs_53; // @[SRAM.scala 145:20:@44552.4]
  reg [31:0] _RAND_53;
  wire  _T_1165; // @[SRAM.scala 148:37:@44553.4]
  wire  _T_1166; // @[SRAM.scala 148:25:@44554.4]
  wire  _T_1167; // @[SRAM.scala 148:15:@44555.4]
  wire  _T_1168; // @[SRAM.scala 149:15:@44557.6]
  wire  _GEN_53; // @[SRAM.scala 148:48:@44556.4]
  reg  regs_54; // @[SRAM.scala 145:20:@44563.4]
  reg [31:0] _RAND_54;
  wire  _T_1174; // @[SRAM.scala 148:37:@44564.4]
  wire  _T_1175; // @[SRAM.scala 148:25:@44565.4]
  wire  _T_1176; // @[SRAM.scala 148:15:@44566.4]
  wire  _T_1177; // @[SRAM.scala 149:15:@44568.6]
  wire  _GEN_54; // @[SRAM.scala 148:48:@44567.4]
  reg  regs_55; // @[SRAM.scala 145:20:@44574.4]
  reg [31:0] _RAND_55;
  wire  _T_1183; // @[SRAM.scala 148:37:@44575.4]
  wire  _T_1184; // @[SRAM.scala 148:25:@44576.4]
  wire  _T_1185; // @[SRAM.scala 148:15:@44577.4]
  wire  _T_1186; // @[SRAM.scala 149:15:@44579.6]
  wire  _GEN_55; // @[SRAM.scala 148:48:@44578.4]
  reg  regs_56; // @[SRAM.scala 145:20:@44585.4]
  reg [31:0] _RAND_56;
  wire  _T_1192; // @[SRAM.scala 148:37:@44586.4]
  wire  _T_1193; // @[SRAM.scala 148:25:@44587.4]
  wire  _T_1194; // @[SRAM.scala 148:15:@44588.4]
  wire  _T_1195; // @[SRAM.scala 149:15:@44590.6]
  wire  _GEN_56; // @[SRAM.scala 148:48:@44589.4]
  reg  regs_57; // @[SRAM.scala 145:20:@44596.4]
  reg [31:0] _RAND_57;
  wire  _T_1201; // @[SRAM.scala 148:37:@44597.4]
  wire  _T_1202; // @[SRAM.scala 148:25:@44598.4]
  wire  _T_1203; // @[SRAM.scala 148:15:@44599.4]
  wire  _T_1204; // @[SRAM.scala 149:15:@44601.6]
  wire  _GEN_57; // @[SRAM.scala 148:48:@44600.4]
  reg  regs_58; // @[SRAM.scala 145:20:@44607.4]
  reg [31:0] _RAND_58;
  wire  _T_1210; // @[SRAM.scala 148:37:@44608.4]
  wire  _T_1211; // @[SRAM.scala 148:25:@44609.4]
  wire  _T_1212; // @[SRAM.scala 148:15:@44610.4]
  wire  _T_1213; // @[SRAM.scala 149:15:@44612.6]
  wire  _GEN_58; // @[SRAM.scala 148:48:@44611.4]
  reg  regs_59; // @[SRAM.scala 145:20:@44618.4]
  reg [31:0] _RAND_59;
  wire  _T_1219; // @[SRAM.scala 148:37:@44619.4]
  wire  _T_1220; // @[SRAM.scala 148:25:@44620.4]
  wire  _T_1221; // @[SRAM.scala 148:15:@44621.4]
  wire  _T_1222; // @[SRAM.scala 149:15:@44623.6]
  wire  _GEN_59; // @[SRAM.scala 148:48:@44622.4]
  reg  regs_60; // @[SRAM.scala 145:20:@44629.4]
  reg [31:0] _RAND_60;
  wire  _T_1228; // @[SRAM.scala 148:37:@44630.4]
  wire  _T_1229; // @[SRAM.scala 148:25:@44631.4]
  wire  _T_1230; // @[SRAM.scala 148:15:@44632.4]
  wire  _T_1231; // @[SRAM.scala 149:15:@44634.6]
  wire  _GEN_60; // @[SRAM.scala 148:48:@44633.4]
  reg  regs_61; // @[SRAM.scala 145:20:@44640.4]
  reg [31:0] _RAND_61;
  wire  _T_1237; // @[SRAM.scala 148:37:@44641.4]
  wire  _T_1238; // @[SRAM.scala 148:25:@44642.4]
  wire  _T_1239; // @[SRAM.scala 148:15:@44643.4]
  wire  _T_1240; // @[SRAM.scala 149:15:@44645.6]
  wire  _GEN_61; // @[SRAM.scala 148:48:@44644.4]
  reg  regs_62; // @[SRAM.scala 145:20:@44651.4]
  reg [31:0] _RAND_62;
  wire  _T_1246; // @[SRAM.scala 148:37:@44652.4]
  wire  _T_1247; // @[SRAM.scala 148:25:@44653.4]
  wire  _T_1248; // @[SRAM.scala 148:15:@44654.4]
  wire  _T_1249; // @[SRAM.scala 149:15:@44656.6]
  wire  _GEN_62; // @[SRAM.scala 148:48:@44655.4]
  reg  regs_63; // @[SRAM.scala 145:20:@44662.4]
  reg [31:0] _RAND_63;
  wire  _T_1255; // @[SRAM.scala 148:37:@44663.4]
  wire  _T_1256; // @[SRAM.scala 148:25:@44664.4]
  wire  _T_1257; // @[SRAM.scala 148:15:@44665.4]
  wire  _T_1258; // @[SRAM.scala 149:15:@44667.6]
  wire  _GEN_63; // @[SRAM.scala 148:48:@44666.4]
  wire  _GEN_65; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_66; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_67; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_68; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_69; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_70; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_71; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_72; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_73; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_74; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_75; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_76; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_77; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_78; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_79; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_80; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_81; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_82; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_83; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_84; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_85; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_86; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_87; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_88; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_89; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_90; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_91; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_92; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_93; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_94; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_95; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_96; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_97; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_98; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_99; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_100; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_101; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_102; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_103; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_104; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_105; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_106; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_107; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_108; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_109; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_110; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_111; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_112; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_113; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_114; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_115; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_116; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_117; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_118; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_119; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_120; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_121; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_122; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_123; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_124; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_125; // @[SRAM.scala 155:12:@44736.4]
  wire  _GEN_126; // @[SRAM.scala 155:12:@44736.4]
  assign _T_688 = io_waddr == 6'h0; // @[SRAM.scala 148:37:@43970.4]
  assign _T_689 = io_wen & _T_688; // @[SRAM.scala 148:25:@43971.4]
  assign _T_690 = io_banks_0_wdata_valid | _T_689; // @[SRAM.scala 148:15:@43972.4]
  assign _T_691 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43974.6]
  assign _GEN_0 = _T_690 ? _T_691 : regs_0; // @[SRAM.scala 148:48:@43973.4]
  assign _T_697 = io_waddr == 6'h1; // @[SRAM.scala 148:37:@43981.4]
  assign _T_698 = io_wen & _T_697; // @[SRAM.scala 148:25:@43982.4]
  assign _T_699 = io_banks_1_wdata_valid | _T_698; // @[SRAM.scala 148:15:@43983.4]
  assign _T_700 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43985.6]
  assign _GEN_1 = _T_699 ? _T_700 : regs_1; // @[SRAM.scala 148:48:@43984.4]
  assign _T_706 = io_waddr == 6'h2; // @[SRAM.scala 148:37:@43992.4]
  assign _T_707 = io_wen & _T_706; // @[SRAM.scala 148:25:@43993.4]
  assign _T_708 = io_banks_2_wdata_valid | _T_707; // @[SRAM.scala 148:15:@43994.4]
  assign _T_709 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@43996.6]
  assign _GEN_2 = _T_708 ? _T_709 : regs_2; // @[SRAM.scala 148:48:@43995.4]
  assign _T_715 = io_waddr == 6'h3; // @[SRAM.scala 148:37:@44003.4]
  assign _T_716 = io_wen & _T_715; // @[SRAM.scala 148:25:@44004.4]
  assign _T_717 = io_banks_3_wdata_valid | _T_716; // @[SRAM.scala 148:15:@44005.4]
  assign _T_718 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44007.6]
  assign _GEN_3 = _T_717 ? _T_718 : regs_3; // @[SRAM.scala 148:48:@44006.4]
  assign _T_724 = io_waddr == 6'h4; // @[SRAM.scala 148:37:@44014.4]
  assign _T_725 = io_wen & _T_724; // @[SRAM.scala 148:25:@44015.4]
  assign _T_726 = io_banks_4_wdata_valid | _T_725; // @[SRAM.scala 148:15:@44016.4]
  assign _T_727 = io_banks_4_wdata_valid ? io_banks_4_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44018.6]
  assign _GEN_4 = _T_726 ? _T_727 : regs_4; // @[SRAM.scala 148:48:@44017.4]
  assign _T_733 = io_waddr == 6'h5; // @[SRAM.scala 148:37:@44025.4]
  assign _T_734 = io_wen & _T_733; // @[SRAM.scala 148:25:@44026.4]
  assign _T_735 = io_banks_5_wdata_valid | _T_734; // @[SRAM.scala 148:15:@44027.4]
  assign _T_736 = io_banks_5_wdata_valid ? io_banks_5_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44029.6]
  assign _GEN_5 = _T_735 ? _T_736 : regs_5; // @[SRAM.scala 148:48:@44028.4]
  assign _T_742 = io_waddr == 6'h6; // @[SRAM.scala 148:37:@44036.4]
  assign _T_743 = io_wen & _T_742; // @[SRAM.scala 148:25:@44037.4]
  assign _T_744 = io_banks_6_wdata_valid | _T_743; // @[SRAM.scala 148:15:@44038.4]
  assign _T_745 = io_banks_6_wdata_valid ? io_banks_6_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44040.6]
  assign _GEN_6 = _T_744 ? _T_745 : regs_6; // @[SRAM.scala 148:48:@44039.4]
  assign _T_751 = io_waddr == 6'h7; // @[SRAM.scala 148:37:@44047.4]
  assign _T_752 = io_wen & _T_751; // @[SRAM.scala 148:25:@44048.4]
  assign _T_753 = io_banks_7_wdata_valid | _T_752; // @[SRAM.scala 148:15:@44049.4]
  assign _T_754 = io_banks_7_wdata_valid ? io_banks_7_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44051.6]
  assign _GEN_7 = _T_753 ? _T_754 : regs_7; // @[SRAM.scala 148:48:@44050.4]
  assign _T_760 = io_waddr == 6'h8; // @[SRAM.scala 148:37:@44058.4]
  assign _T_761 = io_wen & _T_760; // @[SRAM.scala 148:25:@44059.4]
  assign _T_762 = io_banks_8_wdata_valid | _T_761; // @[SRAM.scala 148:15:@44060.4]
  assign _T_763 = io_banks_8_wdata_valid ? io_banks_8_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44062.6]
  assign _GEN_8 = _T_762 ? _T_763 : regs_8; // @[SRAM.scala 148:48:@44061.4]
  assign _T_769 = io_waddr == 6'h9; // @[SRAM.scala 148:37:@44069.4]
  assign _T_770 = io_wen & _T_769; // @[SRAM.scala 148:25:@44070.4]
  assign _T_771 = io_banks_9_wdata_valid | _T_770; // @[SRAM.scala 148:15:@44071.4]
  assign _T_772 = io_banks_9_wdata_valid ? io_banks_9_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44073.6]
  assign _GEN_9 = _T_771 ? _T_772 : regs_9; // @[SRAM.scala 148:48:@44072.4]
  assign _T_778 = io_waddr == 6'ha; // @[SRAM.scala 148:37:@44080.4]
  assign _T_779 = io_wen & _T_778; // @[SRAM.scala 148:25:@44081.4]
  assign _T_780 = io_banks_10_wdata_valid | _T_779; // @[SRAM.scala 148:15:@44082.4]
  assign _T_781 = io_banks_10_wdata_valid ? io_banks_10_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44084.6]
  assign _GEN_10 = _T_780 ? _T_781 : regs_10; // @[SRAM.scala 148:48:@44083.4]
  assign _T_787 = io_waddr == 6'hb; // @[SRAM.scala 148:37:@44091.4]
  assign _T_788 = io_wen & _T_787; // @[SRAM.scala 148:25:@44092.4]
  assign _T_789 = io_banks_11_wdata_valid | _T_788; // @[SRAM.scala 148:15:@44093.4]
  assign _T_790 = io_banks_11_wdata_valid ? io_banks_11_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44095.6]
  assign _GEN_11 = _T_789 ? _T_790 : regs_11; // @[SRAM.scala 148:48:@44094.4]
  assign _T_796 = io_waddr == 6'hc; // @[SRAM.scala 148:37:@44102.4]
  assign _T_797 = io_wen & _T_796; // @[SRAM.scala 148:25:@44103.4]
  assign _T_798 = io_banks_12_wdata_valid | _T_797; // @[SRAM.scala 148:15:@44104.4]
  assign _T_799 = io_banks_12_wdata_valid ? io_banks_12_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44106.6]
  assign _GEN_12 = _T_798 ? _T_799 : regs_12; // @[SRAM.scala 148:48:@44105.4]
  assign _T_805 = io_waddr == 6'hd; // @[SRAM.scala 148:37:@44113.4]
  assign _T_806 = io_wen & _T_805; // @[SRAM.scala 148:25:@44114.4]
  assign _T_807 = io_banks_13_wdata_valid | _T_806; // @[SRAM.scala 148:15:@44115.4]
  assign _T_808 = io_banks_13_wdata_valid ? io_banks_13_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44117.6]
  assign _GEN_13 = _T_807 ? _T_808 : regs_13; // @[SRAM.scala 148:48:@44116.4]
  assign _T_814 = io_waddr == 6'he; // @[SRAM.scala 148:37:@44124.4]
  assign _T_815 = io_wen & _T_814; // @[SRAM.scala 148:25:@44125.4]
  assign _T_816 = io_banks_14_wdata_valid | _T_815; // @[SRAM.scala 148:15:@44126.4]
  assign _T_817 = io_banks_14_wdata_valid ? io_banks_14_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44128.6]
  assign _GEN_14 = _T_816 ? _T_817 : regs_14; // @[SRAM.scala 148:48:@44127.4]
  assign _T_823 = io_waddr == 6'hf; // @[SRAM.scala 148:37:@44135.4]
  assign _T_824 = io_wen & _T_823; // @[SRAM.scala 148:25:@44136.4]
  assign _T_825 = io_banks_15_wdata_valid | _T_824; // @[SRAM.scala 148:15:@44137.4]
  assign _T_826 = io_banks_15_wdata_valid ? io_banks_15_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44139.6]
  assign _GEN_15 = _T_825 ? _T_826 : regs_15; // @[SRAM.scala 148:48:@44138.4]
  assign _T_832 = io_waddr == 6'h10; // @[SRAM.scala 148:37:@44146.4]
  assign _T_833 = io_wen & _T_832; // @[SRAM.scala 148:25:@44147.4]
  assign _T_834 = io_banks_16_wdata_valid | _T_833; // @[SRAM.scala 148:15:@44148.4]
  assign _T_835 = io_banks_16_wdata_valid ? io_banks_16_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44150.6]
  assign _GEN_16 = _T_834 ? _T_835 : regs_16; // @[SRAM.scala 148:48:@44149.4]
  assign _T_841 = io_waddr == 6'h11; // @[SRAM.scala 148:37:@44157.4]
  assign _T_842 = io_wen & _T_841; // @[SRAM.scala 148:25:@44158.4]
  assign _T_843 = io_banks_17_wdata_valid | _T_842; // @[SRAM.scala 148:15:@44159.4]
  assign _T_844 = io_banks_17_wdata_valid ? io_banks_17_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44161.6]
  assign _GEN_17 = _T_843 ? _T_844 : regs_17; // @[SRAM.scala 148:48:@44160.4]
  assign _T_850 = io_waddr == 6'h12; // @[SRAM.scala 148:37:@44168.4]
  assign _T_851 = io_wen & _T_850; // @[SRAM.scala 148:25:@44169.4]
  assign _T_852 = io_banks_18_wdata_valid | _T_851; // @[SRAM.scala 148:15:@44170.4]
  assign _T_853 = io_banks_18_wdata_valid ? io_banks_18_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44172.6]
  assign _GEN_18 = _T_852 ? _T_853 : regs_18; // @[SRAM.scala 148:48:@44171.4]
  assign _T_859 = io_waddr == 6'h13; // @[SRAM.scala 148:37:@44179.4]
  assign _T_860 = io_wen & _T_859; // @[SRAM.scala 148:25:@44180.4]
  assign _T_861 = io_banks_19_wdata_valid | _T_860; // @[SRAM.scala 148:15:@44181.4]
  assign _T_862 = io_banks_19_wdata_valid ? io_banks_19_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44183.6]
  assign _GEN_19 = _T_861 ? _T_862 : regs_19; // @[SRAM.scala 148:48:@44182.4]
  assign _T_868 = io_waddr == 6'h14; // @[SRAM.scala 148:37:@44190.4]
  assign _T_869 = io_wen & _T_868; // @[SRAM.scala 148:25:@44191.4]
  assign _T_870 = io_banks_20_wdata_valid | _T_869; // @[SRAM.scala 148:15:@44192.4]
  assign _T_871 = io_banks_20_wdata_valid ? io_banks_20_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44194.6]
  assign _GEN_20 = _T_870 ? _T_871 : regs_20; // @[SRAM.scala 148:48:@44193.4]
  assign _T_877 = io_waddr == 6'h15; // @[SRAM.scala 148:37:@44201.4]
  assign _T_878 = io_wen & _T_877; // @[SRAM.scala 148:25:@44202.4]
  assign _T_879 = io_banks_21_wdata_valid | _T_878; // @[SRAM.scala 148:15:@44203.4]
  assign _T_880 = io_banks_21_wdata_valid ? io_banks_21_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44205.6]
  assign _GEN_21 = _T_879 ? _T_880 : regs_21; // @[SRAM.scala 148:48:@44204.4]
  assign _T_886 = io_waddr == 6'h16; // @[SRAM.scala 148:37:@44212.4]
  assign _T_887 = io_wen & _T_886; // @[SRAM.scala 148:25:@44213.4]
  assign _T_888 = io_banks_22_wdata_valid | _T_887; // @[SRAM.scala 148:15:@44214.4]
  assign _T_889 = io_banks_22_wdata_valid ? io_banks_22_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44216.6]
  assign _GEN_22 = _T_888 ? _T_889 : regs_22; // @[SRAM.scala 148:48:@44215.4]
  assign _T_895 = io_waddr == 6'h17; // @[SRAM.scala 148:37:@44223.4]
  assign _T_896 = io_wen & _T_895; // @[SRAM.scala 148:25:@44224.4]
  assign _T_897 = io_banks_23_wdata_valid | _T_896; // @[SRAM.scala 148:15:@44225.4]
  assign _T_898 = io_banks_23_wdata_valid ? io_banks_23_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44227.6]
  assign _GEN_23 = _T_897 ? _T_898 : regs_23; // @[SRAM.scala 148:48:@44226.4]
  assign _T_904 = io_waddr == 6'h18; // @[SRAM.scala 148:37:@44234.4]
  assign _T_905 = io_wen & _T_904; // @[SRAM.scala 148:25:@44235.4]
  assign _T_906 = io_banks_24_wdata_valid | _T_905; // @[SRAM.scala 148:15:@44236.4]
  assign _T_907 = io_banks_24_wdata_valid ? io_banks_24_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44238.6]
  assign _GEN_24 = _T_906 ? _T_907 : regs_24; // @[SRAM.scala 148:48:@44237.4]
  assign _T_913 = io_waddr == 6'h19; // @[SRAM.scala 148:37:@44245.4]
  assign _T_914 = io_wen & _T_913; // @[SRAM.scala 148:25:@44246.4]
  assign _T_915 = io_banks_25_wdata_valid | _T_914; // @[SRAM.scala 148:15:@44247.4]
  assign _T_916 = io_banks_25_wdata_valid ? io_banks_25_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44249.6]
  assign _GEN_25 = _T_915 ? _T_916 : regs_25; // @[SRAM.scala 148:48:@44248.4]
  assign _T_922 = io_waddr == 6'h1a; // @[SRAM.scala 148:37:@44256.4]
  assign _T_923 = io_wen & _T_922; // @[SRAM.scala 148:25:@44257.4]
  assign _T_924 = io_banks_26_wdata_valid | _T_923; // @[SRAM.scala 148:15:@44258.4]
  assign _T_925 = io_banks_26_wdata_valid ? io_banks_26_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44260.6]
  assign _GEN_26 = _T_924 ? _T_925 : regs_26; // @[SRAM.scala 148:48:@44259.4]
  assign _T_931 = io_waddr == 6'h1b; // @[SRAM.scala 148:37:@44267.4]
  assign _T_932 = io_wen & _T_931; // @[SRAM.scala 148:25:@44268.4]
  assign _T_933 = io_banks_27_wdata_valid | _T_932; // @[SRAM.scala 148:15:@44269.4]
  assign _T_934 = io_banks_27_wdata_valid ? io_banks_27_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44271.6]
  assign _GEN_27 = _T_933 ? _T_934 : regs_27; // @[SRAM.scala 148:48:@44270.4]
  assign _T_940 = io_waddr == 6'h1c; // @[SRAM.scala 148:37:@44278.4]
  assign _T_941 = io_wen & _T_940; // @[SRAM.scala 148:25:@44279.4]
  assign _T_942 = io_banks_28_wdata_valid | _T_941; // @[SRAM.scala 148:15:@44280.4]
  assign _T_943 = io_banks_28_wdata_valid ? io_banks_28_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44282.6]
  assign _GEN_28 = _T_942 ? _T_943 : regs_28; // @[SRAM.scala 148:48:@44281.4]
  assign _T_949 = io_waddr == 6'h1d; // @[SRAM.scala 148:37:@44289.4]
  assign _T_950 = io_wen & _T_949; // @[SRAM.scala 148:25:@44290.4]
  assign _T_951 = io_banks_29_wdata_valid | _T_950; // @[SRAM.scala 148:15:@44291.4]
  assign _T_952 = io_banks_29_wdata_valid ? io_banks_29_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44293.6]
  assign _GEN_29 = _T_951 ? _T_952 : regs_29; // @[SRAM.scala 148:48:@44292.4]
  assign _T_958 = io_waddr == 6'h1e; // @[SRAM.scala 148:37:@44300.4]
  assign _T_959 = io_wen & _T_958; // @[SRAM.scala 148:25:@44301.4]
  assign _T_960 = io_banks_30_wdata_valid | _T_959; // @[SRAM.scala 148:15:@44302.4]
  assign _T_961 = io_banks_30_wdata_valid ? io_banks_30_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44304.6]
  assign _GEN_30 = _T_960 ? _T_961 : regs_30; // @[SRAM.scala 148:48:@44303.4]
  assign _T_967 = io_waddr == 6'h1f; // @[SRAM.scala 148:37:@44311.4]
  assign _T_968 = io_wen & _T_967; // @[SRAM.scala 148:25:@44312.4]
  assign _T_969 = io_banks_31_wdata_valid | _T_968; // @[SRAM.scala 148:15:@44313.4]
  assign _T_970 = io_banks_31_wdata_valid ? io_banks_31_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44315.6]
  assign _GEN_31 = _T_969 ? _T_970 : regs_31; // @[SRAM.scala 148:48:@44314.4]
  assign _T_976 = io_waddr == 6'h20; // @[SRAM.scala 148:37:@44322.4]
  assign _T_977 = io_wen & _T_976; // @[SRAM.scala 148:25:@44323.4]
  assign _T_978 = io_banks_32_wdata_valid | _T_977; // @[SRAM.scala 148:15:@44324.4]
  assign _T_979 = io_banks_32_wdata_valid ? io_banks_32_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44326.6]
  assign _GEN_32 = _T_978 ? _T_979 : regs_32; // @[SRAM.scala 148:48:@44325.4]
  assign _T_985 = io_waddr == 6'h21; // @[SRAM.scala 148:37:@44333.4]
  assign _T_986 = io_wen & _T_985; // @[SRAM.scala 148:25:@44334.4]
  assign _T_987 = io_banks_33_wdata_valid | _T_986; // @[SRAM.scala 148:15:@44335.4]
  assign _T_988 = io_banks_33_wdata_valid ? io_banks_33_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44337.6]
  assign _GEN_33 = _T_987 ? _T_988 : regs_33; // @[SRAM.scala 148:48:@44336.4]
  assign _T_994 = io_waddr == 6'h22; // @[SRAM.scala 148:37:@44344.4]
  assign _T_995 = io_wen & _T_994; // @[SRAM.scala 148:25:@44345.4]
  assign _T_996 = io_banks_34_wdata_valid | _T_995; // @[SRAM.scala 148:15:@44346.4]
  assign _T_997 = io_banks_34_wdata_valid ? io_banks_34_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44348.6]
  assign _GEN_34 = _T_996 ? _T_997 : regs_34; // @[SRAM.scala 148:48:@44347.4]
  assign _T_1003 = io_waddr == 6'h23; // @[SRAM.scala 148:37:@44355.4]
  assign _T_1004 = io_wen & _T_1003; // @[SRAM.scala 148:25:@44356.4]
  assign _T_1005 = io_banks_35_wdata_valid | _T_1004; // @[SRAM.scala 148:15:@44357.4]
  assign _T_1006 = io_banks_35_wdata_valid ? io_banks_35_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44359.6]
  assign _GEN_35 = _T_1005 ? _T_1006 : regs_35; // @[SRAM.scala 148:48:@44358.4]
  assign _T_1012 = io_waddr == 6'h24; // @[SRAM.scala 148:37:@44366.4]
  assign _T_1013 = io_wen & _T_1012; // @[SRAM.scala 148:25:@44367.4]
  assign _T_1014 = io_banks_36_wdata_valid | _T_1013; // @[SRAM.scala 148:15:@44368.4]
  assign _T_1015 = io_banks_36_wdata_valid ? io_banks_36_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44370.6]
  assign _GEN_36 = _T_1014 ? _T_1015 : regs_36; // @[SRAM.scala 148:48:@44369.4]
  assign _T_1021 = io_waddr == 6'h25; // @[SRAM.scala 148:37:@44377.4]
  assign _T_1022 = io_wen & _T_1021; // @[SRAM.scala 148:25:@44378.4]
  assign _T_1023 = io_banks_37_wdata_valid | _T_1022; // @[SRAM.scala 148:15:@44379.4]
  assign _T_1024 = io_banks_37_wdata_valid ? io_banks_37_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44381.6]
  assign _GEN_37 = _T_1023 ? _T_1024 : regs_37; // @[SRAM.scala 148:48:@44380.4]
  assign _T_1030 = io_waddr == 6'h26; // @[SRAM.scala 148:37:@44388.4]
  assign _T_1031 = io_wen & _T_1030; // @[SRAM.scala 148:25:@44389.4]
  assign _T_1032 = io_banks_38_wdata_valid | _T_1031; // @[SRAM.scala 148:15:@44390.4]
  assign _T_1033 = io_banks_38_wdata_valid ? io_banks_38_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44392.6]
  assign _GEN_38 = _T_1032 ? _T_1033 : regs_38; // @[SRAM.scala 148:48:@44391.4]
  assign _T_1039 = io_waddr == 6'h27; // @[SRAM.scala 148:37:@44399.4]
  assign _T_1040 = io_wen & _T_1039; // @[SRAM.scala 148:25:@44400.4]
  assign _T_1041 = io_banks_39_wdata_valid | _T_1040; // @[SRAM.scala 148:15:@44401.4]
  assign _T_1042 = io_banks_39_wdata_valid ? io_banks_39_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44403.6]
  assign _GEN_39 = _T_1041 ? _T_1042 : regs_39; // @[SRAM.scala 148:48:@44402.4]
  assign _T_1048 = io_waddr == 6'h28; // @[SRAM.scala 148:37:@44410.4]
  assign _T_1049 = io_wen & _T_1048; // @[SRAM.scala 148:25:@44411.4]
  assign _T_1050 = io_banks_40_wdata_valid | _T_1049; // @[SRAM.scala 148:15:@44412.4]
  assign _T_1051 = io_banks_40_wdata_valid ? io_banks_40_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44414.6]
  assign _GEN_40 = _T_1050 ? _T_1051 : regs_40; // @[SRAM.scala 148:48:@44413.4]
  assign _T_1057 = io_waddr == 6'h29; // @[SRAM.scala 148:37:@44421.4]
  assign _T_1058 = io_wen & _T_1057; // @[SRAM.scala 148:25:@44422.4]
  assign _T_1059 = io_banks_41_wdata_valid | _T_1058; // @[SRAM.scala 148:15:@44423.4]
  assign _T_1060 = io_banks_41_wdata_valid ? io_banks_41_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44425.6]
  assign _GEN_41 = _T_1059 ? _T_1060 : regs_41; // @[SRAM.scala 148:48:@44424.4]
  assign _T_1066 = io_waddr == 6'h2a; // @[SRAM.scala 148:37:@44432.4]
  assign _T_1067 = io_wen & _T_1066; // @[SRAM.scala 148:25:@44433.4]
  assign _T_1068 = io_banks_42_wdata_valid | _T_1067; // @[SRAM.scala 148:15:@44434.4]
  assign _T_1069 = io_banks_42_wdata_valid ? io_banks_42_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44436.6]
  assign _GEN_42 = _T_1068 ? _T_1069 : regs_42; // @[SRAM.scala 148:48:@44435.4]
  assign _T_1075 = io_waddr == 6'h2b; // @[SRAM.scala 148:37:@44443.4]
  assign _T_1076 = io_wen & _T_1075; // @[SRAM.scala 148:25:@44444.4]
  assign _T_1077 = io_banks_43_wdata_valid | _T_1076; // @[SRAM.scala 148:15:@44445.4]
  assign _T_1078 = io_banks_43_wdata_valid ? io_banks_43_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44447.6]
  assign _GEN_43 = _T_1077 ? _T_1078 : regs_43; // @[SRAM.scala 148:48:@44446.4]
  assign _T_1084 = io_waddr == 6'h2c; // @[SRAM.scala 148:37:@44454.4]
  assign _T_1085 = io_wen & _T_1084; // @[SRAM.scala 148:25:@44455.4]
  assign _T_1086 = io_banks_44_wdata_valid | _T_1085; // @[SRAM.scala 148:15:@44456.4]
  assign _T_1087 = io_banks_44_wdata_valid ? io_banks_44_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44458.6]
  assign _GEN_44 = _T_1086 ? _T_1087 : regs_44; // @[SRAM.scala 148:48:@44457.4]
  assign _T_1093 = io_waddr == 6'h2d; // @[SRAM.scala 148:37:@44465.4]
  assign _T_1094 = io_wen & _T_1093; // @[SRAM.scala 148:25:@44466.4]
  assign _T_1095 = io_banks_45_wdata_valid | _T_1094; // @[SRAM.scala 148:15:@44467.4]
  assign _T_1096 = io_banks_45_wdata_valid ? io_banks_45_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44469.6]
  assign _GEN_45 = _T_1095 ? _T_1096 : regs_45; // @[SRAM.scala 148:48:@44468.4]
  assign _T_1102 = io_waddr == 6'h2e; // @[SRAM.scala 148:37:@44476.4]
  assign _T_1103 = io_wen & _T_1102; // @[SRAM.scala 148:25:@44477.4]
  assign _T_1104 = io_banks_46_wdata_valid | _T_1103; // @[SRAM.scala 148:15:@44478.4]
  assign _T_1105 = io_banks_46_wdata_valid ? io_banks_46_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44480.6]
  assign _GEN_46 = _T_1104 ? _T_1105 : regs_46; // @[SRAM.scala 148:48:@44479.4]
  assign _T_1111 = io_waddr == 6'h2f; // @[SRAM.scala 148:37:@44487.4]
  assign _T_1112 = io_wen & _T_1111; // @[SRAM.scala 148:25:@44488.4]
  assign _T_1113 = io_banks_47_wdata_valid | _T_1112; // @[SRAM.scala 148:15:@44489.4]
  assign _T_1114 = io_banks_47_wdata_valid ? io_banks_47_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44491.6]
  assign _GEN_47 = _T_1113 ? _T_1114 : regs_47; // @[SRAM.scala 148:48:@44490.4]
  assign _T_1120 = io_waddr == 6'h30; // @[SRAM.scala 148:37:@44498.4]
  assign _T_1121 = io_wen & _T_1120; // @[SRAM.scala 148:25:@44499.4]
  assign _T_1122 = io_banks_48_wdata_valid | _T_1121; // @[SRAM.scala 148:15:@44500.4]
  assign _T_1123 = io_banks_48_wdata_valid ? io_banks_48_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44502.6]
  assign _GEN_48 = _T_1122 ? _T_1123 : regs_48; // @[SRAM.scala 148:48:@44501.4]
  assign _T_1129 = io_waddr == 6'h31; // @[SRAM.scala 148:37:@44509.4]
  assign _T_1130 = io_wen & _T_1129; // @[SRAM.scala 148:25:@44510.4]
  assign _T_1131 = io_banks_49_wdata_valid | _T_1130; // @[SRAM.scala 148:15:@44511.4]
  assign _T_1132 = io_banks_49_wdata_valid ? io_banks_49_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44513.6]
  assign _GEN_49 = _T_1131 ? _T_1132 : regs_49; // @[SRAM.scala 148:48:@44512.4]
  assign _T_1138 = io_waddr == 6'h32; // @[SRAM.scala 148:37:@44520.4]
  assign _T_1139 = io_wen & _T_1138; // @[SRAM.scala 148:25:@44521.4]
  assign _T_1140 = io_banks_50_wdata_valid | _T_1139; // @[SRAM.scala 148:15:@44522.4]
  assign _T_1141 = io_banks_50_wdata_valid ? io_banks_50_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44524.6]
  assign _GEN_50 = _T_1140 ? _T_1141 : regs_50; // @[SRAM.scala 148:48:@44523.4]
  assign _T_1147 = io_waddr == 6'h33; // @[SRAM.scala 148:37:@44531.4]
  assign _T_1148 = io_wen & _T_1147; // @[SRAM.scala 148:25:@44532.4]
  assign _T_1149 = io_banks_51_wdata_valid | _T_1148; // @[SRAM.scala 148:15:@44533.4]
  assign _T_1150 = io_banks_51_wdata_valid ? io_banks_51_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44535.6]
  assign _GEN_51 = _T_1149 ? _T_1150 : regs_51; // @[SRAM.scala 148:48:@44534.4]
  assign _T_1156 = io_waddr == 6'h34; // @[SRAM.scala 148:37:@44542.4]
  assign _T_1157 = io_wen & _T_1156; // @[SRAM.scala 148:25:@44543.4]
  assign _T_1158 = io_banks_52_wdata_valid | _T_1157; // @[SRAM.scala 148:15:@44544.4]
  assign _T_1159 = io_banks_52_wdata_valid ? io_banks_52_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44546.6]
  assign _GEN_52 = _T_1158 ? _T_1159 : regs_52; // @[SRAM.scala 148:48:@44545.4]
  assign _T_1165 = io_waddr == 6'h35; // @[SRAM.scala 148:37:@44553.4]
  assign _T_1166 = io_wen & _T_1165; // @[SRAM.scala 148:25:@44554.4]
  assign _T_1167 = io_banks_53_wdata_valid | _T_1166; // @[SRAM.scala 148:15:@44555.4]
  assign _T_1168 = io_banks_53_wdata_valid ? io_banks_53_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44557.6]
  assign _GEN_53 = _T_1167 ? _T_1168 : regs_53; // @[SRAM.scala 148:48:@44556.4]
  assign _T_1174 = io_waddr == 6'h36; // @[SRAM.scala 148:37:@44564.4]
  assign _T_1175 = io_wen & _T_1174; // @[SRAM.scala 148:25:@44565.4]
  assign _T_1176 = io_banks_54_wdata_valid | _T_1175; // @[SRAM.scala 148:15:@44566.4]
  assign _T_1177 = io_banks_54_wdata_valid ? io_banks_54_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44568.6]
  assign _GEN_54 = _T_1176 ? _T_1177 : regs_54; // @[SRAM.scala 148:48:@44567.4]
  assign _T_1183 = io_waddr == 6'h37; // @[SRAM.scala 148:37:@44575.4]
  assign _T_1184 = io_wen & _T_1183; // @[SRAM.scala 148:25:@44576.4]
  assign _T_1185 = io_banks_55_wdata_valid | _T_1184; // @[SRAM.scala 148:15:@44577.4]
  assign _T_1186 = io_banks_55_wdata_valid ? io_banks_55_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44579.6]
  assign _GEN_55 = _T_1185 ? _T_1186 : regs_55; // @[SRAM.scala 148:48:@44578.4]
  assign _T_1192 = io_waddr == 6'h38; // @[SRAM.scala 148:37:@44586.4]
  assign _T_1193 = io_wen & _T_1192; // @[SRAM.scala 148:25:@44587.4]
  assign _T_1194 = io_banks_56_wdata_valid | _T_1193; // @[SRAM.scala 148:15:@44588.4]
  assign _T_1195 = io_banks_56_wdata_valid ? io_banks_56_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44590.6]
  assign _GEN_56 = _T_1194 ? _T_1195 : regs_56; // @[SRAM.scala 148:48:@44589.4]
  assign _T_1201 = io_waddr == 6'h39; // @[SRAM.scala 148:37:@44597.4]
  assign _T_1202 = io_wen & _T_1201; // @[SRAM.scala 148:25:@44598.4]
  assign _T_1203 = io_banks_57_wdata_valid | _T_1202; // @[SRAM.scala 148:15:@44599.4]
  assign _T_1204 = io_banks_57_wdata_valid ? io_banks_57_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44601.6]
  assign _GEN_57 = _T_1203 ? _T_1204 : regs_57; // @[SRAM.scala 148:48:@44600.4]
  assign _T_1210 = io_waddr == 6'h3a; // @[SRAM.scala 148:37:@44608.4]
  assign _T_1211 = io_wen & _T_1210; // @[SRAM.scala 148:25:@44609.4]
  assign _T_1212 = io_banks_58_wdata_valid | _T_1211; // @[SRAM.scala 148:15:@44610.4]
  assign _T_1213 = io_banks_58_wdata_valid ? io_banks_58_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44612.6]
  assign _GEN_58 = _T_1212 ? _T_1213 : regs_58; // @[SRAM.scala 148:48:@44611.4]
  assign _T_1219 = io_waddr == 6'h3b; // @[SRAM.scala 148:37:@44619.4]
  assign _T_1220 = io_wen & _T_1219; // @[SRAM.scala 148:25:@44620.4]
  assign _T_1221 = io_banks_59_wdata_valid | _T_1220; // @[SRAM.scala 148:15:@44621.4]
  assign _T_1222 = io_banks_59_wdata_valid ? io_banks_59_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44623.6]
  assign _GEN_59 = _T_1221 ? _T_1222 : regs_59; // @[SRAM.scala 148:48:@44622.4]
  assign _T_1228 = io_waddr == 6'h3c; // @[SRAM.scala 148:37:@44630.4]
  assign _T_1229 = io_wen & _T_1228; // @[SRAM.scala 148:25:@44631.4]
  assign _T_1230 = io_banks_60_wdata_valid | _T_1229; // @[SRAM.scala 148:15:@44632.4]
  assign _T_1231 = io_banks_60_wdata_valid ? io_banks_60_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44634.6]
  assign _GEN_60 = _T_1230 ? _T_1231 : regs_60; // @[SRAM.scala 148:48:@44633.4]
  assign _T_1237 = io_waddr == 6'h3d; // @[SRAM.scala 148:37:@44641.4]
  assign _T_1238 = io_wen & _T_1237; // @[SRAM.scala 148:25:@44642.4]
  assign _T_1239 = io_banks_61_wdata_valid | _T_1238; // @[SRAM.scala 148:15:@44643.4]
  assign _T_1240 = io_banks_61_wdata_valid ? io_banks_61_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44645.6]
  assign _GEN_61 = _T_1239 ? _T_1240 : regs_61; // @[SRAM.scala 148:48:@44644.4]
  assign _T_1246 = io_waddr == 6'h3e; // @[SRAM.scala 148:37:@44652.4]
  assign _T_1247 = io_wen & _T_1246; // @[SRAM.scala 148:25:@44653.4]
  assign _T_1248 = io_banks_62_wdata_valid | _T_1247; // @[SRAM.scala 148:15:@44654.4]
  assign _T_1249 = io_banks_62_wdata_valid ? io_banks_62_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44656.6]
  assign _GEN_62 = _T_1248 ? _T_1249 : regs_62; // @[SRAM.scala 148:48:@44655.4]
  assign _T_1255 = io_waddr == 6'h3f; // @[SRAM.scala 148:37:@44663.4]
  assign _T_1256 = io_wen & _T_1255; // @[SRAM.scala 148:25:@44664.4]
  assign _T_1257 = io_banks_63_wdata_valid | _T_1256; // @[SRAM.scala 148:15:@44665.4]
  assign _T_1258 = io_banks_63_wdata_valid ? io_banks_63_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@44667.6]
  assign _GEN_63 = _T_1257 ? _T_1258 : regs_63; // @[SRAM.scala 148:48:@44666.4]
  assign _GEN_65 = 6'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_66 = 6'h2 == io_raddr ? regs_2 : _GEN_65; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_67 = 6'h3 == io_raddr ? regs_3 : _GEN_66; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_68 = 6'h4 == io_raddr ? regs_4 : _GEN_67; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_69 = 6'h5 == io_raddr ? regs_5 : _GEN_68; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_70 = 6'h6 == io_raddr ? regs_6 : _GEN_69; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_71 = 6'h7 == io_raddr ? regs_7 : _GEN_70; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_72 = 6'h8 == io_raddr ? regs_8 : _GEN_71; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_73 = 6'h9 == io_raddr ? regs_9 : _GEN_72; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_74 = 6'ha == io_raddr ? regs_10 : _GEN_73; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_75 = 6'hb == io_raddr ? regs_11 : _GEN_74; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_76 = 6'hc == io_raddr ? regs_12 : _GEN_75; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_77 = 6'hd == io_raddr ? regs_13 : _GEN_76; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_78 = 6'he == io_raddr ? regs_14 : _GEN_77; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_79 = 6'hf == io_raddr ? regs_15 : _GEN_78; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_80 = 6'h10 == io_raddr ? regs_16 : _GEN_79; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_81 = 6'h11 == io_raddr ? regs_17 : _GEN_80; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_82 = 6'h12 == io_raddr ? regs_18 : _GEN_81; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_83 = 6'h13 == io_raddr ? regs_19 : _GEN_82; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_84 = 6'h14 == io_raddr ? regs_20 : _GEN_83; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_85 = 6'h15 == io_raddr ? regs_21 : _GEN_84; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_86 = 6'h16 == io_raddr ? regs_22 : _GEN_85; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_87 = 6'h17 == io_raddr ? regs_23 : _GEN_86; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_88 = 6'h18 == io_raddr ? regs_24 : _GEN_87; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_89 = 6'h19 == io_raddr ? regs_25 : _GEN_88; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_90 = 6'h1a == io_raddr ? regs_26 : _GEN_89; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_91 = 6'h1b == io_raddr ? regs_27 : _GEN_90; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_92 = 6'h1c == io_raddr ? regs_28 : _GEN_91; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_93 = 6'h1d == io_raddr ? regs_29 : _GEN_92; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_94 = 6'h1e == io_raddr ? regs_30 : _GEN_93; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_95 = 6'h1f == io_raddr ? regs_31 : _GEN_94; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_96 = 6'h20 == io_raddr ? regs_32 : _GEN_95; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_97 = 6'h21 == io_raddr ? regs_33 : _GEN_96; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_98 = 6'h22 == io_raddr ? regs_34 : _GEN_97; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_99 = 6'h23 == io_raddr ? regs_35 : _GEN_98; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_100 = 6'h24 == io_raddr ? regs_36 : _GEN_99; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_101 = 6'h25 == io_raddr ? regs_37 : _GEN_100; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_102 = 6'h26 == io_raddr ? regs_38 : _GEN_101; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_103 = 6'h27 == io_raddr ? regs_39 : _GEN_102; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_104 = 6'h28 == io_raddr ? regs_40 : _GEN_103; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_105 = 6'h29 == io_raddr ? regs_41 : _GEN_104; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_106 = 6'h2a == io_raddr ? regs_42 : _GEN_105; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_107 = 6'h2b == io_raddr ? regs_43 : _GEN_106; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_108 = 6'h2c == io_raddr ? regs_44 : _GEN_107; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_109 = 6'h2d == io_raddr ? regs_45 : _GEN_108; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_110 = 6'h2e == io_raddr ? regs_46 : _GEN_109; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_111 = 6'h2f == io_raddr ? regs_47 : _GEN_110; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_112 = 6'h30 == io_raddr ? regs_48 : _GEN_111; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_113 = 6'h31 == io_raddr ? regs_49 : _GEN_112; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_114 = 6'h32 == io_raddr ? regs_50 : _GEN_113; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_115 = 6'h33 == io_raddr ? regs_51 : _GEN_114; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_116 = 6'h34 == io_raddr ? regs_52 : _GEN_115; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_117 = 6'h35 == io_raddr ? regs_53 : _GEN_116; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_118 = 6'h36 == io_raddr ? regs_54 : _GEN_117; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_119 = 6'h37 == io_raddr ? regs_55 : _GEN_118; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_120 = 6'h38 == io_raddr ? regs_56 : _GEN_119; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_121 = 6'h39 == io_raddr ? regs_57 : _GEN_120; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_122 = 6'h3a == io_raddr ? regs_58 : _GEN_121; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_123 = 6'h3b == io_raddr ? regs_59 : _GEN_122; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_124 = 6'h3c == io_raddr ? regs_60 : _GEN_123; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_125 = 6'h3d == io_raddr ? regs_61 : _GEN_124; // @[SRAM.scala 155:12:@44736.4]
  assign _GEN_126 = 6'h3e == io_raddr ? regs_62 : _GEN_125; // @[SRAM.scala 155:12:@44736.4]
  assign io_rdata = 6'h3f == io_raddr ? regs_63 : _GEN_126; // @[SRAM.scala 155:12:@44736.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_690) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_699) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_708) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_717) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_4 <= 1'h0;
    end else begin
      if (_T_726) begin
        if (io_banks_4_wdata_valid) begin
          regs_4 <= io_banks_4_wdata_bits;
        end else begin
          regs_4 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_5 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (io_banks_5_wdata_valid) begin
          regs_5 <= io_banks_5_wdata_bits;
        end else begin
          regs_5 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_6 <= 1'h0;
    end else begin
      if (_T_744) begin
        if (io_banks_6_wdata_valid) begin
          regs_6 <= io_banks_6_wdata_bits;
        end else begin
          regs_6 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_7 <= 1'h0;
    end else begin
      if (_T_753) begin
        if (io_banks_7_wdata_valid) begin
          regs_7 <= io_banks_7_wdata_bits;
        end else begin
          regs_7 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_8 <= 1'h0;
    end else begin
      if (_T_762) begin
        if (io_banks_8_wdata_valid) begin
          regs_8 <= io_banks_8_wdata_bits;
        end else begin
          regs_8 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_9 <= 1'h0;
    end else begin
      if (_T_771) begin
        if (io_banks_9_wdata_valid) begin
          regs_9 <= io_banks_9_wdata_bits;
        end else begin
          regs_9 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_10 <= 1'h0;
    end else begin
      if (_T_780) begin
        if (io_banks_10_wdata_valid) begin
          regs_10 <= io_banks_10_wdata_bits;
        end else begin
          regs_10 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_11 <= 1'h0;
    end else begin
      if (_T_789) begin
        if (io_banks_11_wdata_valid) begin
          regs_11 <= io_banks_11_wdata_bits;
        end else begin
          regs_11 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_12 <= 1'h0;
    end else begin
      if (_T_798) begin
        if (io_banks_12_wdata_valid) begin
          regs_12 <= io_banks_12_wdata_bits;
        end else begin
          regs_12 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_13 <= 1'h0;
    end else begin
      if (_T_807) begin
        if (io_banks_13_wdata_valid) begin
          regs_13 <= io_banks_13_wdata_bits;
        end else begin
          regs_13 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_14 <= 1'h0;
    end else begin
      if (_T_816) begin
        if (io_banks_14_wdata_valid) begin
          regs_14 <= io_banks_14_wdata_bits;
        end else begin
          regs_14 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_15 <= 1'h0;
    end else begin
      if (_T_825) begin
        if (io_banks_15_wdata_valid) begin
          regs_15 <= io_banks_15_wdata_bits;
        end else begin
          regs_15 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_16 <= 1'h0;
    end else begin
      if (_T_834) begin
        if (io_banks_16_wdata_valid) begin
          regs_16 <= io_banks_16_wdata_bits;
        end else begin
          regs_16 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_17 <= 1'h0;
    end else begin
      if (_T_843) begin
        if (io_banks_17_wdata_valid) begin
          regs_17 <= io_banks_17_wdata_bits;
        end else begin
          regs_17 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_18 <= 1'h0;
    end else begin
      if (_T_852) begin
        if (io_banks_18_wdata_valid) begin
          regs_18 <= io_banks_18_wdata_bits;
        end else begin
          regs_18 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_19 <= 1'h0;
    end else begin
      if (_T_861) begin
        if (io_banks_19_wdata_valid) begin
          regs_19 <= io_banks_19_wdata_bits;
        end else begin
          regs_19 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_20 <= 1'h0;
    end else begin
      if (_T_870) begin
        if (io_banks_20_wdata_valid) begin
          regs_20 <= io_banks_20_wdata_bits;
        end else begin
          regs_20 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_21 <= 1'h0;
    end else begin
      if (_T_879) begin
        if (io_banks_21_wdata_valid) begin
          regs_21 <= io_banks_21_wdata_bits;
        end else begin
          regs_21 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_22 <= 1'h0;
    end else begin
      if (_T_888) begin
        if (io_banks_22_wdata_valid) begin
          regs_22 <= io_banks_22_wdata_bits;
        end else begin
          regs_22 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_23 <= 1'h0;
    end else begin
      if (_T_897) begin
        if (io_banks_23_wdata_valid) begin
          regs_23 <= io_banks_23_wdata_bits;
        end else begin
          regs_23 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_24 <= 1'h0;
    end else begin
      if (_T_906) begin
        if (io_banks_24_wdata_valid) begin
          regs_24 <= io_banks_24_wdata_bits;
        end else begin
          regs_24 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_25 <= 1'h0;
    end else begin
      if (_T_915) begin
        if (io_banks_25_wdata_valid) begin
          regs_25 <= io_banks_25_wdata_bits;
        end else begin
          regs_25 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_26 <= 1'h0;
    end else begin
      if (_T_924) begin
        if (io_banks_26_wdata_valid) begin
          regs_26 <= io_banks_26_wdata_bits;
        end else begin
          regs_26 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_27 <= 1'h0;
    end else begin
      if (_T_933) begin
        if (io_banks_27_wdata_valid) begin
          regs_27 <= io_banks_27_wdata_bits;
        end else begin
          regs_27 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_28 <= 1'h0;
    end else begin
      if (_T_942) begin
        if (io_banks_28_wdata_valid) begin
          regs_28 <= io_banks_28_wdata_bits;
        end else begin
          regs_28 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_29 <= 1'h0;
    end else begin
      if (_T_951) begin
        if (io_banks_29_wdata_valid) begin
          regs_29 <= io_banks_29_wdata_bits;
        end else begin
          regs_29 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_30 <= 1'h0;
    end else begin
      if (_T_960) begin
        if (io_banks_30_wdata_valid) begin
          regs_30 <= io_banks_30_wdata_bits;
        end else begin
          regs_30 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_31 <= 1'h0;
    end else begin
      if (_T_969) begin
        if (io_banks_31_wdata_valid) begin
          regs_31 <= io_banks_31_wdata_bits;
        end else begin
          regs_31 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_32 <= 1'h0;
    end else begin
      if (_T_978) begin
        if (io_banks_32_wdata_valid) begin
          regs_32 <= io_banks_32_wdata_bits;
        end else begin
          regs_32 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_33 <= 1'h0;
    end else begin
      if (_T_987) begin
        if (io_banks_33_wdata_valid) begin
          regs_33 <= io_banks_33_wdata_bits;
        end else begin
          regs_33 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_34 <= 1'h0;
    end else begin
      if (_T_996) begin
        if (io_banks_34_wdata_valid) begin
          regs_34 <= io_banks_34_wdata_bits;
        end else begin
          regs_34 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_35 <= 1'h0;
    end else begin
      if (_T_1005) begin
        if (io_banks_35_wdata_valid) begin
          regs_35 <= io_banks_35_wdata_bits;
        end else begin
          regs_35 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_36 <= 1'h0;
    end else begin
      if (_T_1014) begin
        if (io_banks_36_wdata_valid) begin
          regs_36 <= io_banks_36_wdata_bits;
        end else begin
          regs_36 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_37 <= 1'h0;
    end else begin
      if (_T_1023) begin
        if (io_banks_37_wdata_valid) begin
          regs_37 <= io_banks_37_wdata_bits;
        end else begin
          regs_37 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_38 <= 1'h0;
    end else begin
      if (_T_1032) begin
        if (io_banks_38_wdata_valid) begin
          regs_38 <= io_banks_38_wdata_bits;
        end else begin
          regs_38 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_39 <= 1'h0;
    end else begin
      if (_T_1041) begin
        if (io_banks_39_wdata_valid) begin
          regs_39 <= io_banks_39_wdata_bits;
        end else begin
          regs_39 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_40 <= 1'h0;
    end else begin
      if (_T_1050) begin
        if (io_banks_40_wdata_valid) begin
          regs_40 <= io_banks_40_wdata_bits;
        end else begin
          regs_40 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_41 <= 1'h0;
    end else begin
      if (_T_1059) begin
        if (io_banks_41_wdata_valid) begin
          regs_41 <= io_banks_41_wdata_bits;
        end else begin
          regs_41 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_42 <= 1'h0;
    end else begin
      if (_T_1068) begin
        if (io_banks_42_wdata_valid) begin
          regs_42 <= io_banks_42_wdata_bits;
        end else begin
          regs_42 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_43 <= 1'h0;
    end else begin
      if (_T_1077) begin
        if (io_banks_43_wdata_valid) begin
          regs_43 <= io_banks_43_wdata_bits;
        end else begin
          regs_43 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_44 <= 1'h0;
    end else begin
      if (_T_1086) begin
        if (io_banks_44_wdata_valid) begin
          regs_44 <= io_banks_44_wdata_bits;
        end else begin
          regs_44 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_45 <= 1'h0;
    end else begin
      if (_T_1095) begin
        if (io_banks_45_wdata_valid) begin
          regs_45 <= io_banks_45_wdata_bits;
        end else begin
          regs_45 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_46 <= 1'h0;
    end else begin
      if (_T_1104) begin
        if (io_banks_46_wdata_valid) begin
          regs_46 <= io_banks_46_wdata_bits;
        end else begin
          regs_46 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_47 <= 1'h0;
    end else begin
      if (_T_1113) begin
        if (io_banks_47_wdata_valid) begin
          regs_47 <= io_banks_47_wdata_bits;
        end else begin
          regs_47 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_48 <= 1'h0;
    end else begin
      if (_T_1122) begin
        if (io_banks_48_wdata_valid) begin
          regs_48 <= io_banks_48_wdata_bits;
        end else begin
          regs_48 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_49 <= 1'h0;
    end else begin
      if (_T_1131) begin
        if (io_banks_49_wdata_valid) begin
          regs_49 <= io_banks_49_wdata_bits;
        end else begin
          regs_49 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_50 <= 1'h0;
    end else begin
      if (_T_1140) begin
        if (io_banks_50_wdata_valid) begin
          regs_50 <= io_banks_50_wdata_bits;
        end else begin
          regs_50 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_51 <= 1'h0;
    end else begin
      if (_T_1149) begin
        if (io_banks_51_wdata_valid) begin
          regs_51 <= io_banks_51_wdata_bits;
        end else begin
          regs_51 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_52 <= 1'h0;
    end else begin
      if (_T_1158) begin
        if (io_banks_52_wdata_valid) begin
          regs_52 <= io_banks_52_wdata_bits;
        end else begin
          regs_52 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_53 <= 1'h0;
    end else begin
      if (_T_1167) begin
        if (io_banks_53_wdata_valid) begin
          regs_53 <= io_banks_53_wdata_bits;
        end else begin
          regs_53 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_54 <= 1'h0;
    end else begin
      if (_T_1176) begin
        if (io_banks_54_wdata_valid) begin
          regs_54 <= io_banks_54_wdata_bits;
        end else begin
          regs_54 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_55 <= 1'h0;
    end else begin
      if (_T_1185) begin
        if (io_banks_55_wdata_valid) begin
          regs_55 <= io_banks_55_wdata_bits;
        end else begin
          regs_55 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_56 <= 1'h0;
    end else begin
      if (_T_1194) begin
        if (io_banks_56_wdata_valid) begin
          regs_56 <= io_banks_56_wdata_bits;
        end else begin
          regs_56 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_57 <= 1'h0;
    end else begin
      if (_T_1203) begin
        if (io_banks_57_wdata_valid) begin
          regs_57 <= io_banks_57_wdata_bits;
        end else begin
          regs_57 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_58 <= 1'h0;
    end else begin
      if (_T_1212) begin
        if (io_banks_58_wdata_valid) begin
          regs_58 <= io_banks_58_wdata_bits;
        end else begin
          regs_58 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_59 <= 1'h0;
    end else begin
      if (_T_1221) begin
        if (io_banks_59_wdata_valid) begin
          regs_59 <= io_banks_59_wdata_bits;
        end else begin
          regs_59 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_60 <= 1'h0;
    end else begin
      if (_T_1230) begin
        if (io_banks_60_wdata_valid) begin
          regs_60 <= io_banks_60_wdata_bits;
        end else begin
          regs_60 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_61 <= 1'h0;
    end else begin
      if (_T_1239) begin
        if (io_banks_61_wdata_valid) begin
          regs_61 <= io_banks_61_wdata_bits;
        end else begin
          regs_61 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_62 <= 1'h0;
    end else begin
      if (_T_1248) begin
        if (io_banks_62_wdata_valid) begin
          regs_62 <= io_banks_62_wdata_bits;
        end else begin
          regs_62 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_63 <= 1'h0;
    end else begin
      if (_T_1257) begin
        if (io_banks_63_wdata_valid) begin
          regs_63 <= io_banks_63_wdata_bits;
        end else begin
          regs_63 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_33( // @[:@44738.2]
  input   clock, // @[:@44739.4]
  input   reset, // @[:@44740.4]
  output  io_in_ready, // @[:@44741.4]
  input   io_in_valid, // @[:@44741.4]
  input   io_in_bits, // @[:@44741.4]
  input   io_out_ready, // @[:@44741.4]
  output  io_out_valid, // @[:@44741.4]
  output  io_out_bits, // @[:@44741.4]
  input   io_banks_0_wdata_valid, // @[:@44741.4]
  input   io_banks_0_wdata_bits, // @[:@44741.4]
  input   io_banks_1_wdata_valid, // @[:@44741.4]
  input   io_banks_1_wdata_bits, // @[:@44741.4]
  input   io_banks_2_wdata_valid, // @[:@44741.4]
  input   io_banks_2_wdata_bits, // @[:@44741.4]
  input   io_banks_3_wdata_valid, // @[:@44741.4]
  input   io_banks_3_wdata_bits, // @[:@44741.4]
  input   io_banks_4_wdata_valid, // @[:@44741.4]
  input   io_banks_4_wdata_bits, // @[:@44741.4]
  input   io_banks_5_wdata_valid, // @[:@44741.4]
  input   io_banks_5_wdata_bits, // @[:@44741.4]
  input   io_banks_6_wdata_valid, // @[:@44741.4]
  input   io_banks_6_wdata_bits, // @[:@44741.4]
  input   io_banks_7_wdata_valid, // @[:@44741.4]
  input   io_banks_7_wdata_bits, // @[:@44741.4]
  input   io_banks_8_wdata_valid, // @[:@44741.4]
  input   io_banks_8_wdata_bits, // @[:@44741.4]
  input   io_banks_9_wdata_valid, // @[:@44741.4]
  input   io_banks_9_wdata_bits, // @[:@44741.4]
  input   io_banks_10_wdata_valid, // @[:@44741.4]
  input   io_banks_10_wdata_bits, // @[:@44741.4]
  input   io_banks_11_wdata_valid, // @[:@44741.4]
  input   io_banks_11_wdata_bits, // @[:@44741.4]
  input   io_banks_12_wdata_valid, // @[:@44741.4]
  input   io_banks_12_wdata_bits, // @[:@44741.4]
  input   io_banks_13_wdata_valid, // @[:@44741.4]
  input   io_banks_13_wdata_bits, // @[:@44741.4]
  input   io_banks_14_wdata_valid, // @[:@44741.4]
  input   io_banks_14_wdata_bits, // @[:@44741.4]
  input   io_banks_15_wdata_valid, // @[:@44741.4]
  input   io_banks_15_wdata_bits, // @[:@44741.4]
  input   io_banks_16_wdata_valid, // @[:@44741.4]
  input   io_banks_16_wdata_bits, // @[:@44741.4]
  input   io_banks_17_wdata_valid, // @[:@44741.4]
  input   io_banks_17_wdata_bits, // @[:@44741.4]
  input   io_banks_18_wdata_valid, // @[:@44741.4]
  input   io_banks_18_wdata_bits, // @[:@44741.4]
  input   io_banks_19_wdata_valid, // @[:@44741.4]
  input   io_banks_19_wdata_bits, // @[:@44741.4]
  input   io_banks_20_wdata_valid, // @[:@44741.4]
  input   io_banks_20_wdata_bits, // @[:@44741.4]
  input   io_banks_21_wdata_valid, // @[:@44741.4]
  input   io_banks_21_wdata_bits, // @[:@44741.4]
  input   io_banks_22_wdata_valid, // @[:@44741.4]
  input   io_banks_22_wdata_bits, // @[:@44741.4]
  input   io_banks_23_wdata_valid, // @[:@44741.4]
  input   io_banks_23_wdata_bits, // @[:@44741.4]
  input   io_banks_24_wdata_valid, // @[:@44741.4]
  input   io_banks_24_wdata_bits, // @[:@44741.4]
  input   io_banks_25_wdata_valid, // @[:@44741.4]
  input   io_banks_25_wdata_bits, // @[:@44741.4]
  input   io_banks_26_wdata_valid, // @[:@44741.4]
  input   io_banks_26_wdata_bits, // @[:@44741.4]
  input   io_banks_27_wdata_valid, // @[:@44741.4]
  input   io_banks_27_wdata_bits, // @[:@44741.4]
  input   io_banks_28_wdata_valid, // @[:@44741.4]
  input   io_banks_28_wdata_bits, // @[:@44741.4]
  input   io_banks_29_wdata_valid, // @[:@44741.4]
  input   io_banks_29_wdata_bits, // @[:@44741.4]
  input   io_banks_30_wdata_valid, // @[:@44741.4]
  input   io_banks_30_wdata_bits, // @[:@44741.4]
  input   io_banks_31_wdata_valid, // @[:@44741.4]
  input   io_banks_31_wdata_bits, // @[:@44741.4]
  input   io_banks_32_wdata_valid, // @[:@44741.4]
  input   io_banks_32_wdata_bits, // @[:@44741.4]
  input   io_banks_33_wdata_valid, // @[:@44741.4]
  input   io_banks_33_wdata_bits, // @[:@44741.4]
  input   io_banks_34_wdata_valid, // @[:@44741.4]
  input   io_banks_34_wdata_bits, // @[:@44741.4]
  input   io_banks_35_wdata_valid, // @[:@44741.4]
  input   io_banks_35_wdata_bits, // @[:@44741.4]
  input   io_banks_36_wdata_valid, // @[:@44741.4]
  input   io_banks_36_wdata_bits, // @[:@44741.4]
  input   io_banks_37_wdata_valid, // @[:@44741.4]
  input   io_banks_37_wdata_bits, // @[:@44741.4]
  input   io_banks_38_wdata_valid, // @[:@44741.4]
  input   io_banks_38_wdata_bits, // @[:@44741.4]
  input   io_banks_39_wdata_valid, // @[:@44741.4]
  input   io_banks_39_wdata_bits, // @[:@44741.4]
  input   io_banks_40_wdata_valid, // @[:@44741.4]
  input   io_banks_40_wdata_bits, // @[:@44741.4]
  input   io_banks_41_wdata_valid, // @[:@44741.4]
  input   io_banks_41_wdata_bits, // @[:@44741.4]
  input   io_banks_42_wdata_valid, // @[:@44741.4]
  input   io_banks_42_wdata_bits, // @[:@44741.4]
  input   io_banks_43_wdata_valid, // @[:@44741.4]
  input   io_banks_43_wdata_bits, // @[:@44741.4]
  input   io_banks_44_wdata_valid, // @[:@44741.4]
  input   io_banks_44_wdata_bits, // @[:@44741.4]
  input   io_banks_45_wdata_valid, // @[:@44741.4]
  input   io_banks_45_wdata_bits, // @[:@44741.4]
  input   io_banks_46_wdata_valid, // @[:@44741.4]
  input   io_banks_46_wdata_bits, // @[:@44741.4]
  input   io_banks_47_wdata_valid, // @[:@44741.4]
  input   io_banks_47_wdata_bits, // @[:@44741.4]
  input   io_banks_48_wdata_valid, // @[:@44741.4]
  input   io_banks_48_wdata_bits, // @[:@44741.4]
  input   io_banks_49_wdata_valid, // @[:@44741.4]
  input   io_banks_49_wdata_bits, // @[:@44741.4]
  input   io_banks_50_wdata_valid, // @[:@44741.4]
  input   io_banks_50_wdata_bits, // @[:@44741.4]
  input   io_banks_51_wdata_valid, // @[:@44741.4]
  input   io_banks_51_wdata_bits, // @[:@44741.4]
  input   io_banks_52_wdata_valid, // @[:@44741.4]
  input   io_banks_52_wdata_bits, // @[:@44741.4]
  input   io_banks_53_wdata_valid, // @[:@44741.4]
  input   io_banks_53_wdata_bits, // @[:@44741.4]
  input   io_banks_54_wdata_valid, // @[:@44741.4]
  input   io_banks_54_wdata_bits, // @[:@44741.4]
  input   io_banks_55_wdata_valid, // @[:@44741.4]
  input   io_banks_55_wdata_bits, // @[:@44741.4]
  input   io_banks_56_wdata_valid, // @[:@44741.4]
  input   io_banks_56_wdata_bits, // @[:@44741.4]
  input   io_banks_57_wdata_valid, // @[:@44741.4]
  input   io_banks_57_wdata_bits, // @[:@44741.4]
  input   io_banks_58_wdata_valid, // @[:@44741.4]
  input   io_banks_58_wdata_bits, // @[:@44741.4]
  input   io_banks_59_wdata_valid, // @[:@44741.4]
  input   io_banks_59_wdata_bits, // @[:@44741.4]
  input   io_banks_60_wdata_valid, // @[:@44741.4]
  input   io_banks_60_wdata_bits, // @[:@44741.4]
  input   io_banks_61_wdata_valid, // @[:@44741.4]
  input   io_banks_61_wdata_bits, // @[:@44741.4]
  input   io_banks_62_wdata_valid, // @[:@44741.4]
  input   io_banks_62_wdata_bits, // @[:@44741.4]
  input   io_banks_63_wdata_valid, // @[:@44741.4]
  input   io_banks_63_wdata_bits // @[:@44741.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@45007.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@45007.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@45007.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@45007.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@45007.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@45017.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@45017.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@45017.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@45017.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@45017.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@45032.4]
  wire [5:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@45032.4]
  wire [5:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_4_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_4_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_5_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_5_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_6_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_6_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_7_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_7_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_8_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_8_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_9_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_9_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_10_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_10_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_11_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_11_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_12_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_12_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_13_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_13_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_14_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_14_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_15_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_15_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_16_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_16_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_17_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_17_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_18_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_18_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_19_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_19_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_20_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_20_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_21_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_21_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_22_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_22_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_23_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_23_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_24_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_24_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_25_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_25_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_26_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_26_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_27_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_27_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_28_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_28_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_29_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_29_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_30_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_30_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_31_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_31_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_32_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_32_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_33_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_33_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_34_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_34_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_35_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_35_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_36_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_36_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_37_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_37_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_38_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_38_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_39_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_39_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_40_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_40_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_41_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_41_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_42_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_42_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_43_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_43_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_44_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_44_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_45_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_45_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_46_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_46_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_47_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_47_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_48_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_48_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_49_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_49_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_50_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_50_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_51_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_51_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_52_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_52_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_53_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_53_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_54_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_54_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_55_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_55_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_56_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_56_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_57_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_57_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_58_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_58_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_59_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_59_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_60_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_60_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_61_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_61_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_62_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_62_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_63_wdata_valid; // @[FIFO.scala 49:19:@45032.4]
  wire  FFRAM_io_banks_63_wdata_bits; // @[FIFO.scala 49:19:@45032.4]
  wire  writeEn; // @[FIFO.scala 30:29:@45005.4]
  wire  readEn; // @[FIFO.scala 31:29:@45006.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@45027.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@45028.4]
  wire  _T_824; // @[FIFO.scala 45:27:@45029.4]
  wire  empty; // @[FIFO.scala 45:24:@45030.4]
  wire  full; // @[FIFO.scala 46:23:@45031.4]
  wire  _T_1657; // @[FIFO.scala 83:17:@46198.4]
  wire  _GEN_64; // @[FIFO.scala 83:29:@46199.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@45007.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@45017.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM_16 FFRAM ( // @[FIFO.scala 49:19:@45032.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(FFRAM_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(FFRAM_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(FFRAM_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(FFRAM_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(FFRAM_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(FFRAM_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(FFRAM_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(FFRAM_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(FFRAM_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(FFRAM_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(FFRAM_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(FFRAM_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(FFRAM_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(FFRAM_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(FFRAM_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(FFRAM_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(FFRAM_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(FFRAM_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(FFRAM_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(FFRAM_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(FFRAM_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(FFRAM_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(FFRAM_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(FFRAM_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(FFRAM_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(FFRAM_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(FFRAM_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(FFRAM_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(FFRAM_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(FFRAM_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(FFRAM_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(FFRAM_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(FFRAM_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(FFRAM_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(FFRAM_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(FFRAM_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(FFRAM_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(FFRAM_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(FFRAM_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(FFRAM_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(FFRAM_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(FFRAM_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(FFRAM_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(FFRAM_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(FFRAM_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(FFRAM_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(FFRAM_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(FFRAM_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(FFRAM_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(FFRAM_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(FFRAM_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(FFRAM_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(FFRAM_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(FFRAM_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(FFRAM_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(FFRAM_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(FFRAM_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(FFRAM_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(FFRAM_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(FFRAM_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(FFRAM_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(FFRAM_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(FFRAM_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(FFRAM_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(FFRAM_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(FFRAM_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(FFRAM_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(FFRAM_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(FFRAM_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(FFRAM_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(FFRAM_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(FFRAM_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(FFRAM_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(FFRAM_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(FFRAM_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(FFRAM_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(FFRAM_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(FFRAM_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(FFRAM_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(FFRAM_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(FFRAM_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(FFRAM_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(FFRAM_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(FFRAM_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(FFRAM_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(FFRAM_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(FFRAM_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(FFRAM_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(FFRAM_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(FFRAM_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(FFRAM_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(FFRAM_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(FFRAM_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(FFRAM_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(FFRAM_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(FFRAM_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(FFRAM_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(FFRAM_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(FFRAM_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(FFRAM_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(FFRAM_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(FFRAM_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(FFRAM_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(FFRAM_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(FFRAM_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(FFRAM_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(FFRAM_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(FFRAM_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(FFRAM_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(FFRAM_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(FFRAM_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(FFRAM_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(FFRAM_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(FFRAM_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(FFRAM_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(FFRAM_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(FFRAM_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(FFRAM_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(FFRAM_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(FFRAM_io_banks_63_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@45005.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@45006.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@45028.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@45029.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@45030.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@45031.4]
  assign _T_1657 = writeEn != readEn; // @[FIFO.scala 83:17:@46198.4]
  assign _GEN_64 = _T_1657 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@46199.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@46205.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@46203.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@45237.4]
  assign enqCounter_clock = clock; // @[:@45008.4]
  assign enqCounter_reset = reset; // @[:@45009.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@45015.4]
  assign deqCounter_clock = clock; // @[:@45018.4]
  assign deqCounter_reset = reset; // @[:@45019.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@45025.4]
  assign FFRAM_clock = clock; // @[:@45033.4]
  assign FFRAM_reset = reset; // @[:@45034.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@45233.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@45234.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@45235.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@45236.4]
  assign FFRAM_io_banks_0_wdata_valid = io_banks_0_wdata_valid; // @[FIFO.scala 59:15:@45239.4]
  assign FFRAM_io_banks_0_wdata_bits = io_banks_0_wdata_bits; // @[FIFO.scala 59:15:@45238.4]
  assign FFRAM_io_banks_1_wdata_valid = io_banks_1_wdata_valid; // @[FIFO.scala 59:15:@45242.4]
  assign FFRAM_io_banks_1_wdata_bits = io_banks_1_wdata_bits; // @[FIFO.scala 59:15:@45241.4]
  assign FFRAM_io_banks_2_wdata_valid = io_banks_2_wdata_valid; // @[FIFO.scala 59:15:@45245.4]
  assign FFRAM_io_banks_2_wdata_bits = io_banks_2_wdata_bits; // @[FIFO.scala 59:15:@45244.4]
  assign FFRAM_io_banks_3_wdata_valid = io_banks_3_wdata_valid; // @[FIFO.scala 59:15:@45248.4]
  assign FFRAM_io_banks_3_wdata_bits = io_banks_3_wdata_bits; // @[FIFO.scala 59:15:@45247.4]
  assign FFRAM_io_banks_4_wdata_valid = io_banks_4_wdata_valid; // @[FIFO.scala 59:15:@45251.4]
  assign FFRAM_io_banks_4_wdata_bits = io_banks_4_wdata_bits; // @[FIFO.scala 59:15:@45250.4]
  assign FFRAM_io_banks_5_wdata_valid = io_banks_5_wdata_valid; // @[FIFO.scala 59:15:@45254.4]
  assign FFRAM_io_banks_5_wdata_bits = io_banks_5_wdata_bits; // @[FIFO.scala 59:15:@45253.4]
  assign FFRAM_io_banks_6_wdata_valid = io_banks_6_wdata_valid; // @[FIFO.scala 59:15:@45257.4]
  assign FFRAM_io_banks_6_wdata_bits = io_banks_6_wdata_bits; // @[FIFO.scala 59:15:@45256.4]
  assign FFRAM_io_banks_7_wdata_valid = io_banks_7_wdata_valid; // @[FIFO.scala 59:15:@45260.4]
  assign FFRAM_io_banks_7_wdata_bits = io_banks_7_wdata_bits; // @[FIFO.scala 59:15:@45259.4]
  assign FFRAM_io_banks_8_wdata_valid = io_banks_8_wdata_valid; // @[FIFO.scala 59:15:@45263.4]
  assign FFRAM_io_banks_8_wdata_bits = io_banks_8_wdata_bits; // @[FIFO.scala 59:15:@45262.4]
  assign FFRAM_io_banks_9_wdata_valid = io_banks_9_wdata_valid; // @[FIFO.scala 59:15:@45266.4]
  assign FFRAM_io_banks_9_wdata_bits = io_banks_9_wdata_bits; // @[FIFO.scala 59:15:@45265.4]
  assign FFRAM_io_banks_10_wdata_valid = io_banks_10_wdata_valid; // @[FIFO.scala 59:15:@45269.4]
  assign FFRAM_io_banks_10_wdata_bits = io_banks_10_wdata_bits; // @[FIFO.scala 59:15:@45268.4]
  assign FFRAM_io_banks_11_wdata_valid = io_banks_11_wdata_valid; // @[FIFO.scala 59:15:@45272.4]
  assign FFRAM_io_banks_11_wdata_bits = io_banks_11_wdata_bits; // @[FIFO.scala 59:15:@45271.4]
  assign FFRAM_io_banks_12_wdata_valid = io_banks_12_wdata_valid; // @[FIFO.scala 59:15:@45275.4]
  assign FFRAM_io_banks_12_wdata_bits = io_banks_12_wdata_bits; // @[FIFO.scala 59:15:@45274.4]
  assign FFRAM_io_banks_13_wdata_valid = io_banks_13_wdata_valid; // @[FIFO.scala 59:15:@45278.4]
  assign FFRAM_io_banks_13_wdata_bits = io_banks_13_wdata_bits; // @[FIFO.scala 59:15:@45277.4]
  assign FFRAM_io_banks_14_wdata_valid = io_banks_14_wdata_valid; // @[FIFO.scala 59:15:@45281.4]
  assign FFRAM_io_banks_14_wdata_bits = io_banks_14_wdata_bits; // @[FIFO.scala 59:15:@45280.4]
  assign FFRAM_io_banks_15_wdata_valid = io_banks_15_wdata_valid; // @[FIFO.scala 59:15:@45284.4]
  assign FFRAM_io_banks_15_wdata_bits = io_banks_15_wdata_bits; // @[FIFO.scala 59:15:@45283.4]
  assign FFRAM_io_banks_16_wdata_valid = io_banks_16_wdata_valid; // @[FIFO.scala 59:15:@45287.4]
  assign FFRAM_io_banks_16_wdata_bits = io_banks_16_wdata_bits; // @[FIFO.scala 59:15:@45286.4]
  assign FFRAM_io_banks_17_wdata_valid = io_banks_17_wdata_valid; // @[FIFO.scala 59:15:@45290.4]
  assign FFRAM_io_banks_17_wdata_bits = io_banks_17_wdata_bits; // @[FIFO.scala 59:15:@45289.4]
  assign FFRAM_io_banks_18_wdata_valid = io_banks_18_wdata_valid; // @[FIFO.scala 59:15:@45293.4]
  assign FFRAM_io_banks_18_wdata_bits = io_banks_18_wdata_bits; // @[FIFO.scala 59:15:@45292.4]
  assign FFRAM_io_banks_19_wdata_valid = io_banks_19_wdata_valid; // @[FIFO.scala 59:15:@45296.4]
  assign FFRAM_io_banks_19_wdata_bits = io_banks_19_wdata_bits; // @[FIFO.scala 59:15:@45295.4]
  assign FFRAM_io_banks_20_wdata_valid = io_banks_20_wdata_valid; // @[FIFO.scala 59:15:@45299.4]
  assign FFRAM_io_banks_20_wdata_bits = io_banks_20_wdata_bits; // @[FIFO.scala 59:15:@45298.4]
  assign FFRAM_io_banks_21_wdata_valid = io_banks_21_wdata_valid; // @[FIFO.scala 59:15:@45302.4]
  assign FFRAM_io_banks_21_wdata_bits = io_banks_21_wdata_bits; // @[FIFO.scala 59:15:@45301.4]
  assign FFRAM_io_banks_22_wdata_valid = io_banks_22_wdata_valid; // @[FIFO.scala 59:15:@45305.4]
  assign FFRAM_io_banks_22_wdata_bits = io_banks_22_wdata_bits; // @[FIFO.scala 59:15:@45304.4]
  assign FFRAM_io_banks_23_wdata_valid = io_banks_23_wdata_valid; // @[FIFO.scala 59:15:@45308.4]
  assign FFRAM_io_banks_23_wdata_bits = io_banks_23_wdata_bits; // @[FIFO.scala 59:15:@45307.4]
  assign FFRAM_io_banks_24_wdata_valid = io_banks_24_wdata_valid; // @[FIFO.scala 59:15:@45311.4]
  assign FFRAM_io_banks_24_wdata_bits = io_banks_24_wdata_bits; // @[FIFO.scala 59:15:@45310.4]
  assign FFRAM_io_banks_25_wdata_valid = io_banks_25_wdata_valid; // @[FIFO.scala 59:15:@45314.4]
  assign FFRAM_io_banks_25_wdata_bits = io_banks_25_wdata_bits; // @[FIFO.scala 59:15:@45313.4]
  assign FFRAM_io_banks_26_wdata_valid = io_banks_26_wdata_valid; // @[FIFO.scala 59:15:@45317.4]
  assign FFRAM_io_banks_26_wdata_bits = io_banks_26_wdata_bits; // @[FIFO.scala 59:15:@45316.4]
  assign FFRAM_io_banks_27_wdata_valid = io_banks_27_wdata_valid; // @[FIFO.scala 59:15:@45320.4]
  assign FFRAM_io_banks_27_wdata_bits = io_banks_27_wdata_bits; // @[FIFO.scala 59:15:@45319.4]
  assign FFRAM_io_banks_28_wdata_valid = io_banks_28_wdata_valid; // @[FIFO.scala 59:15:@45323.4]
  assign FFRAM_io_banks_28_wdata_bits = io_banks_28_wdata_bits; // @[FIFO.scala 59:15:@45322.4]
  assign FFRAM_io_banks_29_wdata_valid = io_banks_29_wdata_valid; // @[FIFO.scala 59:15:@45326.4]
  assign FFRAM_io_banks_29_wdata_bits = io_banks_29_wdata_bits; // @[FIFO.scala 59:15:@45325.4]
  assign FFRAM_io_banks_30_wdata_valid = io_banks_30_wdata_valid; // @[FIFO.scala 59:15:@45329.4]
  assign FFRAM_io_banks_30_wdata_bits = io_banks_30_wdata_bits; // @[FIFO.scala 59:15:@45328.4]
  assign FFRAM_io_banks_31_wdata_valid = io_banks_31_wdata_valid; // @[FIFO.scala 59:15:@45332.4]
  assign FFRAM_io_banks_31_wdata_bits = io_banks_31_wdata_bits; // @[FIFO.scala 59:15:@45331.4]
  assign FFRAM_io_banks_32_wdata_valid = io_banks_32_wdata_valid; // @[FIFO.scala 59:15:@45335.4]
  assign FFRAM_io_banks_32_wdata_bits = io_banks_32_wdata_bits; // @[FIFO.scala 59:15:@45334.4]
  assign FFRAM_io_banks_33_wdata_valid = io_banks_33_wdata_valid; // @[FIFO.scala 59:15:@45338.4]
  assign FFRAM_io_banks_33_wdata_bits = io_banks_33_wdata_bits; // @[FIFO.scala 59:15:@45337.4]
  assign FFRAM_io_banks_34_wdata_valid = io_banks_34_wdata_valid; // @[FIFO.scala 59:15:@45341.4]
  assign FFRAM_io_banks_34_wdata_bits = io_banks_34_wdata_bits; // @[FIFO.scala 59:15:@45340.4]
  assign FFRAM_io_banks_35_wdata_valid = io_banks_35_wdata_valid; // @[FIFO.scala 59:15:@45344.4]
  assign FFRAM_io_banks_35_wdata_bits = io_banks_35_wdata_bits; // @[FIFO.scala 59:15:@45343.4]
  assign FFRAM_io_banks_36_wdata_valid = io_banks_36_wdata_valid; // @[FIFO.scala 59:15:@45347.4]
  assign FFRAM_io_banks_36_wdata_bits = io_banks_36_wdata_bits; // @[FIFO.scala 59:15:@45346.4]
  assign FFRAM_io_banks_37_wdata_valid = io_banks_37_wdata_valid; // @[FIFO.scala 59:15:@45350.4]
  assign FFRAM_io_banks_37_wdata_bits = io_banks_37_wdata_bits; // @[FIFO.scala 59:15:@45349.4]
  assign FFRAM_io_banks_38_wdata_valid = io_banks_38_wdata_valid; // @[FIFO.scala 59:15:@45353.4]
  assign FFRAM_io_banks_38_wdata_bits = io_banks_38_wdata_bits; // @[FIFO.scala 59:15:@45352.4]
  assign FFRAM_io_banks_39_wdata_valid = io_banks_39_wdata_valid; // @[FIFO.scala 59:15:@45356.4]
  assign FFRAM_io_banks_39_wdata_bits = io_banks_39_wdata_bits; // @[FIFO.scala 59:15:@45355.4]
  assign FFRAM_io_banks_40_wdata_valid = io_banks_40_wdata_valid; // @[FIFO.scala 59:15:@45359.4]
  assign FFRAM_io_banks_40_wdata_bits = io_banks_40_wdata_bits; // @[FIFO.scala 59:15:@45358.4]
  assign FFRAM_io_banks_41_wdata_valid = io_banks_41_wdata_valid; // @[FIFO.scala 59:15:@45362.4]
  assign FFRAM_io_banks_41_wdata_bits = io_banks_41_wdata_bits; // @[FIFO.scala 59:15:@45361.4]
  assign FFRAM_io_banks_42_wdata_valid = io_banks_42_wdata_valid; // @[FIFO.scala 59:15:@45365.4]
  assign FFRAM_io_banks_42_wdata_bits = io_banks_42_wdata_bits; // @[FIFO.scala 59:15:@45364.4]
  assign FFRAM_io_banks_43_wdata_valid = io_banks_43_wdata_valid; // @[FIFO.scala 59:15:@45368.4]
  assign FFRAM_io_banks_43_wdata_bits = io_banks_43_wdata_bits; // @[FIFO.scala 59:15:@45367.4]
  assign FFRAM_io_banks_44_wdata_valid = io_banks_44_wdata_valid; // @[FIFO.scala 59:15:@45371.4]
  assign FFRAM_io_banks_44_wdata_bits = io_banks_44_wdata_bits; // @[FIFO.scala 59:15:@45370.4]
  assign FFRAM_io_banks_45_wdata_valid = io_banks_45_wdata_valid; // @[FIFO.scala 59:15:@45374.4]
  assign FFRAM_io_banks_45_wdata_bits = io_banks_45_wdata_bits; // @[FIFO.scala 59:15:@45373.4]
  assign FFRAM_io_banks_46_wdata_valid = io_banks_46_wdata_valid; // @[FIFO.scala 59:15:@45377.4]
  assign FFRAM_io_banks_46_wdata_bits = io_banks_46_wdata_bits; // @[FIFO.scala 59:15:@45376.4]
  assign FFRAM_io_banks_47_wdata_valid = io_banks_47_wdata_valid; // @[FIFO.scala 59:15:@45380.4]
  assign FFRAM_io_banks_47_wdata_bits = io_banks_47_wdata_bits; // @[FIFO.scala 59:15:@45379.4]
  assign FFRAM_io_banks_48_wdata_valid = io_banks_48_wdata_valid; // @[FIFO.scala 59:15:@45383.4]
  assign FFRAM_io_banks_48_wdata_bits = io_banks_48_wdata_bits; // @[FIFO.scala 59:15:@45382.4]
  assign FFRAM_io_banks_49_wdata_valid = io_banks_49_wdata_valid; // @[FIFO.scala 59:15:@45386.4]
  assign FFRAM_io_banks_49_wdata_bits = io_banks_49_wdata_bits; // @[FIFO.scala 59:15:@45385.4]
  assign FFRAM_io_banks_50_wdata_valid = io_banks_50_wdata_valid; // @[FIFO.scala 59:15:@45389.4]
  assign FFRAM_io_banks_50_wdata_bits = io_banks_50_wdata_bits; // @[FIFO.scala 59:15:@45388.4]
  assign FFRAM_io_banks_51_wdata_valid = io_banks_51_wdata_valid; // @[FIFO.scala 59:15:@45392.4]
  assign FFRAM_io_banks_51_wdata_bits = io_banks_51_wdata_bits; // @[FIFO.scala 59:15:@45391.4]
  assign FFRAM_io_banks_52_wdata_valid = io_banks_52_wdata_valid; // @[FIFO.scala 59:15:@45395.4]
  assign FFRAM_io_banks_52_wdata_bits = io_banks_52_wdata_bits; // @[FIFO.scala 59:15:@45394.4]
  assign FFRAM_io_banks_53_wdata_valid = io_banks_53_wdata_valid; // @[FIFO.scala 59:15:@45398.4]
  assign FFRAM_io_banks_53_wdata_bits = io_banks_53_wdata_bits; // @[FIFO.scala 59:15:@45397.4]
  assign FFRAM_io_banks_54_wdata_valid = io_banks_54_wdata_valid; // @[FIFO.scala 59:15:@45401.4]
  assign FFRAM_io_banks_54_wdata_bits = io_banks_54_wdata_bits; // @[FIFO.scala 59:15:@45400.4]
  assign FFRAM_io_banks_55_wdata_valid = io_banks_55_wdata_valid; // @[FIFO.scala 59:15:@45404.4]
  assign FFRAM_io_banks_55_wdata_bits = io_banks_55_wdata_bits; // @[FIFO.scala 59:15:@45403.4]
  assign FFRAM_io_banks_56_wdata_valid = io_banks_56_wdata_valid; // @[FIFO.scala 59:15:@45407.4]
  assign FFRAM_io_banks_56_wdata_bits = io_banks_56_wdata_bits; // @[FIFO.scala 59:15:@45406.4]
  assign FFRAM_io_banks_57_wdata_valid = io_banks_57_wdata_valid; // @[FIFO.scala 59:15:@45410.4]
  assign FFRAM_io_banks_57_wdata_bits = io_banks_57_wdata_bits; // @[FIFO.scala 59:15:@45409.4]
  assign FFRAM_io_banks_58_wdata_valid = io_banks_58_wdata_valid; // @[FIFO.scala 59:15:@45413.4]
  assign FFRAM_io_banks_58_wdata_bits = io_banks_58_wdata_bits; // @[FIFO.scala 59:15:@45412.4]
  assign FFRAM_io_banks_59_wdata_valid = io_banks_59_wdata_valid; // @[FIFO.scala 59:15:@45416.4]
  assign FFRAM_io_banks_59_wdata_bits = io_banks_59_wdata_bits; // @[FIFO.scala 59:15:@45415.4]
  assign FFRAM_io_banks_60_wdata_valid = io_banks_60_wdata_valid; // @[FIFO.scala 59:15:@45419.4]
  assign FFRAM_io_banks_60_wdata_bits = io_banks_60_wdata_bits; // @[FIFO.scala 59:15:@45418.4]
  assign FFRAM_io_banks_61_wdata_valid = io_banks_61_wdata_valid; // @[FIFO.scala 59:15:@45422.4]
  assign FFRAM_io_banks_61_wdata_bits = io_banks_61_wdata_bits; // @[FIFO.scala 59:15:@45421.4]
  assign FFRAM_io_banks_62_wdata_valid = io_banks_62_wdata_valid; // @[FIFO.scala 59:15:@45425.4]
  assign FFRAM_io_banks_62_wdata_bits = io_banks_62_wdata_bits; // @[FIFO.scala 59:15:@45424.4]
  assign FFRAM_io_banks_63_wdata_valid = io_banks_63_wdata_valid; // @[FIFO.scala 59:15:@45428.4]
  assign FFRAM_io_banks_63_wdata_bits = io_banks_63_wdata_bits; // @[FIFO.scala 59:15:@45427.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_1657) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module StreamControllerStore( // @[:@46207.2]
  input         clock, // @[:@46208.4]
  input         reset, // @[:@46209.4]
  input         io_dram_cmd_ready, // @[:@46210.4]
  output        io_dram_cmd_valid, // @[:@46210.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@46210.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@46210.4]
  input         io_dram_wdata_ready, // @[:@46210.4]
  output        io_dram_wdata_valid, // @[:@46210.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@46210.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@46210.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@46210.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@46210.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@46210.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@46210.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@46210.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@46210.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@46210.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@46210.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@46210.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@46210.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@46210.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@46210.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@46210.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@46210.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@46210.4]
  output        io_dram_wresp_ready, // @[:@46210.4]
  input         io_dram_wresp_valid, // @[:@46210.4]
  output        io_store_cmd_ready, // @[:@46210.4]
  input         io_store_cmd_valid, // @[:@46210.4]
  input  [63:0] io_store_cmd_bits_addr, // @[:@46210.4]
  input  [31:0] io_store_cmd_bits_size, // @[:@46210.4]
  output        io_store_data_ready, // @[:@46210.4]
  input         io_store_data_valid, // @[:@46210.4]
  input  [31:0] io_store_data_bits_wdata_0, // @[:@46210.4]
  input         io_store_data_bits_wstrb, // @[:@46210.4]
  input         io_store_wresp_ready, // @[:@46210.4]
  output        io_store_wresp_valid, // @[:@46210.4]
  output        io_store_wresp_bits // @[:@46210.4]
);
  wire  cmd_clock; // @[StreamController.scala 75:19:@46335.4]
  wire  cmd_reset; // @[StreamController.scala 75:19:@46335.4]
  wire  cmd_io_in_ready; // @[StreamController.scala 75:19:@46335.4]
  wire  cmd_io_in_valid; // @[StreamController.scala 75:19:@46335.4]
  wire [63:0] cmd_io_in_bits_addr; // @[StreamController.scala 75:19:@46335.4]
  wire [31:0] cmd_io_in_bits_size; // @[StreamController.scala 75:19:@46335.4]
  wire  cmd_io_out_ready; // @[StreamController.scala 75:19:@46335.4]
  wire  cmd_io_out_valid; // @[StreamController.scala 75:19:@46335.4]
  wire [63:0] cmd_io_out_bits_addr; // @[StreamController.scala 75:19:@46335.4]
  wire [31:0] cmd_io_out_bits_size; // @[StreamController.scala 75:19:@46335.4]
  wire  wdata_clock; // @[StreamController.scala 88:21:@46741.4]
  wire  wdata_reset; // @[StreamController.scala 88:21:@46741.4]
  wire  wdata_io_in_ready; // @[StreamController.scala 88:21:@46741.4]
  wire  wdata_io_in_valid; // @[StreamController.scala 88:21:@46741.4]
  wire [31:0] wdata_io_in_bits_data_0; // @[StreamController.scala 88:21:@46741.4]
  wire  wdata_io_in_bits_strobe; // @[StreamController.scala 88:21:@46741.4]
  wire  wdata_io_out_ready; // @[StreamController.scala 88:21:@46741.4]
  wire  wdata_io_out_valid; // @[StreamController.scala 88:21:@46741.4]
  wire [31:0] wdata_io_out_bits_data_0; // @[StreamController.scala 88:21:@46741.4]
  wire [31:0] wdata_io_out_bits_data_1; // @[StreamController.scala 88:21:@46741.4]
  wire [31:0] wdata_io_out_bits_data_2; // @[StreamController.scala 88:21:@46741.4]
  wire [31:0] wdata_io_out_bits_data_3; // @[StreamController.scala 88:21:@46741.4]
  wire [31:0] wdata_io_out_bits_data_4; // @[StreamController.scala 88:21:@46741.4]
  wire [31:0] wdata_io_out_bits_data_5; // @[StreamController.scala 88:21:@46741.4]
  wire [31:0] wdata_io_out_bits_data_6; // @[StreamController.scala 88:21:@46741.4]
  wire [31:0] wdata_io_out_bits_data_7; // @[StreamController.scala 88:21:@46741.4]
  wire [31:0] wdata_io_out_bits_data_8; // @[StreamController.scala 88:21:@46741.4]
  wire [31:0] wdata_io_out_bits_data_9; // @[StreamController.scala 88:21:@46741.4]
  wire [31:0] wdata_io_out_bits_data_10; // @[StreamController.scala 88:21:@46741.4]
  wire [31:0] wdata_io_out_bits_data_11; // @[StreamController.scala 88:21:@46741.4]
  wire [31:0] wdata_io_out_bits_data_12; // @[StreamController.scala 88:21:@46741.4]
  wire [31:0] wdata_io_out_bits_data_13; // @[StreamController.scala 88:21:@46741.4]
  wire [31:0] wdata_io_out_bits_data_14; // @[StreamController.scala 88:21:@46741.4]
  wire [31:0] wdata_io_out_bits_data_15; // @[StreamController.scala 88:21:@46741.4]
  wire [63:0] wdata_io_out_bits_strobe; // @[StreamController.scala 88:21:@46741.4]
  wire  wresp_clock; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_reset; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_in_ready; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_in_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_in_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_out_ready; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_out_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_out_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_0_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_0_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_1_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_1_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_2_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_2_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_3_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_3_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_4_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_4_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_5_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_5_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_6_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_6_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_7_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_7_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_8_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_8_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_9_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_9_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_10_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_10_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_11_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_11_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_12_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_12_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_13_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_13_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_14_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_14_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_15_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_15_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_16_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_16_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_17_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_17_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_18_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_18_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_19_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_19_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_20_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_20_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_21_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_21_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_22_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_22_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_23_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_23_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_24_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_24_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_25_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_25_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_26_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_26_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_27_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_27_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_28_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_28_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_29_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_29_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_30_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_30_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_31_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_31_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_32_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_32_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_33_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_33_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_34_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_34_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_35_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_35_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_36_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_36_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_37_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_37_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_38_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_38_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_39_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_39_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_40_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_40_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_41_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_41_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_42_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_42_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_43_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_43_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_44_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_44_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_45_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_45_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_46_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_46_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_47_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_47_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_48_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_48_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_49_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_49_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_50_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_50_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_51_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_51_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_52_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_52_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_53_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_53_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_54_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_54_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_55_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_55_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_56_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_56_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_57_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_57_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_58_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_58_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_59_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_59_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_60_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_60_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_61_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_61_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_62_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_62_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_63_wdata_valid; // @[StreamController.scala 100:21:@46982.4]
  wire  wresp_io_banks_63_wdata_bits; // @[StreamController.scala 100:21:@46982.4]
  wire [25:0] _T_111; // @[StreamController.scala 21:10:@46738.4]
  FIFO cmd ( // @[StreamController.scala 75:19:@46335.4]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_in_ready(cmd_io_in_ready),
    .io_in_valid(cmd_io_in_valid),
    .io_in_bits_addr(cmd_io_in_bits_addr),
    .io_in_bits_size(cmd_io_in_bits_size),
    .io_out_ready(cmd_io_out_ready),
    .io_out_valid(cmd_io_out_valid),
    .io_out_bits_addr(cmd_io_out_bits_addr),
    .io_out_bits_size(cmd_io_out_bits_size)
  );
  FIFOWidthConvert wdata ( // @[StreamController.scala 88:21:@46741.4]
    .clock(wdata_clock),
    .reset(wdata_reset),
    .io_in_ready(wdata_io_in_ready),
    .io_in_valid(wdata_io_in_valid),
    .io_in_bits_data_0(wdata_io_in_bits_data_0),
    .io_in_bits_strobe(wdata_io_in_bits_strobe),
    .io_out_ready(wdata_io_out_ready),
    .io_out_valid(wdata_io_out_valid),
    .io_out_bits_data_0(wdata_io_out_bits_data_0),
    .io_out_bits_data_1(wdata_io_out_bits_data_1),
    .io_out_bits_data_2(wdata_io_out_bits_data_2),
    .io_out_bits_data_3(wdata_io_out_bits_data_3),
    .io_out_bits_data_4(wdata_io_out_bits_data_4),
    .io_out_bits_data_5(wdata_io_out_bits_data_5),
    .io_out_bits_data_6(wdata_io_out_bits_data_6),
    .io_out_bits_data_7(wdata_io_out_bits_data_7),
    .io_out_bits_data_8(wdata_io_out_bits_data_8),
    .io_out_bits_data_9(wdata_io_out_bits_data_9),
    .io_out_bits_data_10(wdata_io_out_bits_data_10),
    .io_out_bits_data_11(wdata_io_out_bits_data_11),
    .io_out_bits_data_12(wdata_io_out_bits_data_12),
    .io_out_bits_data_13(wdata_io_out_bits_data_13),
    .io_out_bits_data_14(wdata_io_out_bits_data_14),
    .io_out_bits_data_15(wdata_io_out_bits_data_15),
    .io_out_bits_strobe(wdata_io_out_bits_strobe)
  );
  FIFO_33 wresp ( // @[StreamController.scala 100:21:@46982.4]
    .clock(wresp_clock),
    .reset(wresp_reset),
    .io_in_ready(wresp_io_in_ready),
    .io_in_valid(wresp_io_in_valid),
    .io_in_bits(wresp_io_in_bits),
    .io_out_ready(wresp_io_out_ready),
    .io_out_valid(wresp_io_out_valid),
    .io_out_bits(wresp_io_out_bits),
    .io_banks_0_wdata_valid(wresp_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(wresp_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(wresp_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(wresp_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(wresp_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(wresp_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(wresp_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(wresp_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(wresp_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(wresp_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(wresp_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(wresp_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(wresp_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(wresp_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(wresp_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(wresp_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(wresp_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(wresp_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(wresp_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(wresp_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(wresp_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(wresp_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(wresp_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(wresp_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(wresp_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(wresp_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(wresp_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(wresp_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(wresp_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(wresp_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(wresp_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(wresp_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(wresp_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(wresp_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(wresp_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(wresp_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(wresp_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(wresp_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(wresp_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(wresp_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(wresp_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(wresp_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(wresp_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(wresp_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(wresp_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(wresp_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(wresp_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(wresp_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(wresp_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(wresp_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(wresp_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(wresp_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(wresp_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(wresp_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(wresp_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(wresp_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(wresp_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(wresp_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(wresp_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(wresp_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(wresp_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(wresp_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(wresp_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(wresp_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(wresp_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(wresp_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(wresp_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(wresp_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(wresp_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(wresp_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(wresp_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(wresp_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(wresp_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(wresp_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(wresp_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(wresp_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(wresp_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(wresp_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(wresp_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(wresp_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(wresp_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(wresp_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(wresp_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(wresp_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(wresp_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(wresp_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(wresp_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(wresp_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(wresp_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(wresp_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(wresp_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(wresp_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(wresp_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(wresp_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(wresp_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(wresp_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(wresp_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(wresp_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(wresp_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(wresp_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(wresp_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(wresp_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(wresp_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(wresp_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(wresp_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(wresp_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(wresp_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(wresp_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(wresp_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(wresp_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(wresp_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(wresp_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(wresp_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(wresp_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(wresp_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(wresp_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(wresp_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(wresp_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(wresp_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(wresp_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(wresp_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(wresp_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(wresp_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(wresp_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(wresp_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(wresp_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(wresp_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(wresp_io_banks_63_wdata_bits)
  );
  assign _T_111 = cmd_io_out_bits_size[31:6]; // @[StreamController.scala 21:10:@46738.4]
  assign io_dram_cmd_valid = cmd_io_out_valid; // @[StreamController.scala 81:21:@46735.4]
  assign io_dram_cmd_bits_addr = cmd_io_out_bits_addr; // @[StreamController.scala 83:25:@46736.4]
  assign io_dram_cmd_bits_size = {{6'd0}, _T_111}; // @[StreamController.scala 85:25:@46739.4]
  assign io_dram_wdata_valid = wdata_io_out_valid; // @[StreamController.scala 95:23:@46771.4]
  assign io_dram_wdata_bits_wdata_0 = wdata_io_out_bits_data_0; // @[StreamController.scala 96:28:@46772.4]
  assign io_dram_wdata_bits_wdata_1 = wdata_io_out_bits_data_1; // @[StreamController.scala 96:28:@46773.4]
  assign io_dram_wdata_bits_wdata_2 = wdata_io_out_bits_data_2; // @[StreamController.scala 96:28:@46774.4]
  assign io_dram_wdata_bits_wdata_3 = wdata_io_out_bits_data_3; // @[StreamController.scala 96:28:@46775.4]
  assign io_dram_wdata_bits_wdata_4 = wdata_io_out_bits_data_4; // @[StreamController.scala 96:28:@46776.4]
  assign io_dram_wdata_bits_wdata_5 = wdata_io_out_bits_data_5; // @[StreamController.scala 96:28:@46777.4]
  assign io_dram_wdata_bits_wdata_6 = wdata_io_out_bits_data_6; // @[StreamController.scala 96:28:@46778.4]
  assign io_dram_wdata_bits_wdata_7 = wdata_io_out_bits_data_7; // @[StreamController.scala 96:28:@46779.4]
  assign io_dram_wdata_bits_wdata_8 = wdata_io_out_bits_data_8; // @[StreamController.scala 96:28:@46780.4]
  assign io_dram_wdata_bits_wdata_9 = wdata_io_out_bits_data_9; // @[StreamController.scala 96:28:@46781.4]
  assign io_dram_wdata_bits_wdata_10 = wdata_io_out_bits_data_10; // @[StreamController.scala 96:28:@46782.4]
  assign io_dram_wdata_bits_wdata_11 = wdata_io_out_bits_data_11; // @[StreamController.scala 96:28:@46783.4]
  assign io_dram_wdata_bits_wdata_12 = wdata_io_out_bits_data_12; // @[StreamController.scala 96:28:@46784.4]
  assign io_dram_wdata_bits_wdata_13 = wdata_io_out_bits_data_13; // @[StreamController.scala 96:28:@46785.4]
  assign io_dram_wdata_bits_wdata_14 = wdata_io_out_bits_data_14; // @[StreamController.scala 96:28:@46786.4]
  assign io_dram_wdata_bits_wdata_15 = wdata_io_out_bits_data_15; // @[StreamController.scala 96:28:@46787.4]
  assign io_dram_wdata_bits_wstrb_0 = wdata_io_out_bits_strobe[63]; // @[StreamController.scala 97:28:@46917.4]
  assign io_dram_wdata_bits_wstrb_1 = wdata_io_out_bits_strobe[62]; // @[StreamController.scala 97:28:@46918.4]
  assign io_dram_wdata_bits_wstrb_2 = wdata_io_out_bits_strobe[61]; // @[StreamController.scala 97:28:@46919.4]
  assign io_dram_wdata_bits_wstrb_3 = wdata_io_out_bits_strobe[60]; // @[StreamController.scala 97:28:@46920.4]
  assign io_dram_wdata_bits_wstrb_4 = wdata_io_out_bits_strobe[59]; // @[StreamController.scala 97:28:@46921.4]
  assign io_dram_wdata_bits_wstrb_5 = wdata_io_out_bits_strobe[58]; // @[StreamController.scala 97:28:@46922.4]
  assign io_dram_wdata_bits_wstrb_6 = wdata_io_out_bits_strobe[57]; // @[StreamController.scala 97:28:@46923.4]
  assign io_dram_wdata_bits_wstrb_7 = wdata_io_out_bits_strobe[56]; // @[StreamController.scala 97:28:@46924.4]
  assign io_dram_wdata_bits_wstrb_8 = wdata_io_out_bits_strobe[55]; // @[StreamController.scala 97:28:@46925.4]
  assign io_dram_wdata_bits_wstrb_9 = wdata_io_out_bits_strobe[54]; // @[StreamController.scala 97:28:@46926.4]
  assign io_dram_wdata_bits_wstrb_10 = wdata_io_out_bits_strobe[53]; // @[StreamController.scala 97:28:@46927.4]
  assign io_dram_wdata_bits_wstrb_11 = wdata_io_out_bits_strobe[52]; // @[StreamController.scala 97:28:@46928.4]
  assign io_dram_wdata_bits_wstrb_12 = wdata_io_out_bits_strobe[51]; // @[StreamController.scala 97:28:@46929.4]
  assign io_dram_wdata_bits_wstrb_13 = wdata_io_out_bits_strobe[50]; // @[StreamController.scala 97:28:@46930.4]
  assign io_dram_wdata_bits_wstrb_14 = wdata_io_out_bits_strobe[49]; // @[StreamController.scala 97:28:@46931.4]
  assign io_dram_wdata_bits_wstrb_15 = wdata_io_out_bits_strobe[48]; // @[StreamController.scala 97:28:@46932.4]
  assign io_dram_wdata_bits_wstrb_16 = wdata_io_out_bits_strobe[47]; // @[StreamController.scala 97:28:@46933.4]
  assign io_dram_wdata_bits_wstrb_17 = wdata_io_out_bits_strobe[46]; // @[StreamController.scala 97:28:@46934.4]
  assign io_dram_wdata_bits_wstrb_18 = wdata_io_out_bits_strobe[45]; // @[StreamController.scala 97:28:@46935.4]
  assign io_dram_wdata_bits_wstrb_19 = wdata_io_out_bits_strobe[44]; // @[StreamController.scala 97:28:@46936.4]
  assign io_dram_wdata_bits_wstrb_20 = wdata_io_out_bits_strobe[43]; // @[StreamController.scala 97:28:@46937.4]
  assign io_dram_wdata_bits_wstrb_21 = wdata_io_out_bits_strobe[42]; // @[StreamController.scala 97:28:@46938.4]
  assign io_dram_wdata_bits_wstrb_22 = wdata_io_out_bits_strobe[41]; // @[StreamController.scala 97:28:@46939.4]
  assign io_dram_wdata_bits_wstrb_23 = wdata_io_out_bits_strobe[40]; // @[StreamController.scala 97:28:@46940.4]
  assign io_dram_wdata_bits_wstrb_24 = wdata_io_out_bits_strobe[39]; // @[StreamController.scala 97:28:@46941.4]
  assign io_dram_wdata_bits_wstrb_25 = wdata_io_out_bits_strobe[38]; // @[StreamController.scala 97:28:@46942.4]
  assign io_dram_wdata_bits_wstrb_26 = wdata_io_out_bits_strobe[37]; // @[StreamController.scala 97:28:@46943.4]
  assign io_dram_wdata_bits_wstrb_27 = wdata_io_out_bits_strobe[36]; // @[StreamController.scala 97:28:@46944.4]
  assign io_dram_wdata_bits_wstrb_28 = wdata_io_out_bits_strobe[35]; // @[StreamController.scala 97:28:@46945.4]
  assign io_dram_wdata_bits_wstrb_29 = wdata_io_out_bits_strobe[34]; // @[StreamController.scala 97:28:@46946.4]
  assign io_dram_wdata_bits_wstrb_30 = wdata_io_out_bits_strobe[33]; // @[StreamController.scala 97:28:@46947.4]
  assign io_dram_wdata_bits_wstrb_31 = wdata_io_out_bits_strobe[32]; // @[StreamController.scala 97:28:@46948.4]
  assign io_dram_wdata_bits_wstrb_32 = wdata_io_out_bits_strobe[31]; // @[StreamController.scala 97:28:@46949.4]
  assign io_dram_wdata_bits_wstrb_33 = wdata_io_out_bits_strobe[30]; // @[StreamController.scala 97:28:@46950.4]
  assign io_dram_wdata_bits_wstrb_34 = wdata_io_out_bits_strobe[29]; // @[StreamController.scala 97:28:@46951.4]
  assign io_dram_wdata_bits_wstrb_35 = wdata_io_out_bits_strobe[28]; // @[StreamController.scala 97:28:@46952.4]
  assign io_dram_wdata_bits_wstrb_36 = wdata_io_out_bits_strobe[27]; // @[StreamController.scala 97:28:@46953.4]
  assign io_dram_wdata_bits_wstrb_37 = wdata_io_out_bits_strobe[26]; // @[StreamController.scala 97:28:@46954.4]
  assign io_dram_wdata_bits_wstrb_38 = wdata_io_out_bits_strobe[25]; // @[StreamController.scala 97:28:@46955.4]
  assign io_dram_wdata_bits_wstrb_39 = wdata_io_out_bits_strobe[24]; // @[StreamController.scala 97:28:@46956.4]
  assign io_dram_wdata_bits_wstrb_40 = wdata_io_out_bits_strobe[23]; // @[StreamController.scala 97:28:@46957.4]
  assign io_dram_wdata_bits_wstrb_41 = wdata_io_out_bits_strobe[22]; // @[StreamController.scala 97:28:@46958.4]
  assign io_dram_wdata_bits_wstrb_42 = wdata_io_out_bits_strobe[21]; // @[StreamController.scala 97:28:@46959.4]
  assign io_dram_wdata_bits_wstrb_43 = wdata_io_out_bits_strobe[20]; // @[StreamController.scala 97:28:@46960.4]
  assign io_dram_wdata_bits_wstrb_44 = wdata_io_out_bits_strobe[19]; // @[StreamController.scala 97:28:@46961.4]
  assign io_dram_wdata_bits_wstrb_45 = wdata_io_out_bits_strobe[18]; // @[StreamController.scala 97:28:@46962.4]
  assign io_dram_wdata_bits_wstrb_46 = wdata_io_out_bits_strobe[17]; // @[StreamController.scala 97:28:@46963.4]
  assign io_dram_wdata_bits_wstrb_47 = wdata_io_out_bits_strobe[16]; // @[StreamController.scala 97:28:@46964.4]
  assign io_dram_wdata_bits_wstrb_48 = wdata_io_out_bits_strobe[15]; // @[StreamController.scala 97:28:@46965.4]
  assign io_dram_wdata_bits_wstrb_49 = wdata_io_out_bits_strobe[14]; // @[StreamController.scala 97:28:@46966.4]
  assign io_dram_wdata_bits_wstrb_50 = wdata_io_out_bits_strobe[13]; // @[StreamController.scala 97:28:@46967.4]
  assign io_dram_wdata_bits_wstrb_51 = wdata_io_out_bits_strobe[12]; // @[StreamController.scala 97:28:@46968.4]
  assign io_dram_wdata_bits_wstrb_52 = wdata_io_out_bits_strobe[11]; // @[StreamController.scala 97:28:@46969.4]
  assign io_dram_wdata_bits_wstrb_53 = wdata_io_out_bits_strobe[10]; // @[StreamController.scala 97:28:@46970.4]
  assign io_dram_wdata_bits_wstrb_54 = wdata_io_out_bits_strobe[9]; // @[StreamController.scala 97:28:@46971.4]
  assign io_dram_wdata_bits_wstrb_55 = wdata_io_out_bits_strobe[8]; // @[StreamController.scala 97:28:@46972.4]
  assign io_dram_wdata_bits_wstrb_56 = wdata_io_out_bits_strobe[7]; // @[StreamController.scala 97:28:@46973.4]
  assign io_dram_wdata_bits_wstrb_57 = wdata_io_out_bits_strobe[6]; // @[StreamController.scala 97:28:@46974.4]
  assign io_dram_wdata_bits_wstrb_58 = wdata_io_out_bits_strobe[5]; // @[StreamController.scala 97:28:@46975.4]
  assign io_dram_wdata_bits_wstrb_59 = wdata_io_out_bits_strobe[4]; // @[StreamController.scala 97:28:@46976.4]
  assign io_dram_wdata_bits_wstrb_60 = wdata_io_out_bits_strobe[3]; // @[StreamController.scala 97:28:@46977.4]
  assign io_dram_wdata_bits_wstrb_61 = wdata_io_out_bits_strobe[2]; // @[StreamController.scala 97:28:@46978.4]
  assign io_dram_wdata_bits_wstrb_62 = wdata_io_out_bits_strobe[1]; // @[StreamController.scala 97:28:@46979.4]
  assign io_dram_wdata_bits_wstrb_63 = wdata_io_out_bits_strobe[0]; // @[StreamController.scala 97:28:@46980.4]
  assign io_dram_wresp_ready = wresp_io_in_ready; // @[StreamController.scala 104:23:@47249.4]
  assign io_store_cmd_ready = cmd_io_in_ready; // @[StreamController.scala 79:22:@46733.4]
  assign io_store_data_ready = wdata_io_in_ready; // @[StreamController.scala 93:23:@46770.4]
  assign io_store_wresp_valid = wresp_io_out_valid; // @[StreamController.scala 106:24:@47250.4]
  assign io_store_wresp_bits = wresp_io_out_bits; // @[StreamController.scala 107:23:@47251.4]
  assign cmd_clock = clock; // @[:@46336.4]
  assign cmd_reset = reset; // @[:@46337.4]
  assign cmd_io_in_valid = io_store_cmd_valid; // @[StreamController.scala 77:19:@46730.4]
  assign cmd_io_in_bits_addr = io_store_cmd_bits_addr; // @[StreamController.scala 78:18:@46732.4]
  assign cmd_io_in_bits_size = io_store_cmd_bits_size; // @[StreamController.scala 78:18:@46731.4]
  assign cmd_io_out_ready = io_dram_cmd_ready; // @[StreamController.scala 80:20:@46734.4]
  assign wdata_clock = clock; // @[:@46742.4]
  assign wdata_reset = reset; // @[:@46743.4]
  assign wdata_io_in_valid = io_store_data_valid; // @[StreamController.scala 90:21:@46767.4]
  assign wdata_io_in_bits_data_0 = io_store_data_bits_wdata_0; // @[StreamController.scala 91:25:@46768.4]
  assign wdata_io_in_bits_strobe = io_store_data_bits_wstrb; // @[StreamController.scala 92:27:@46769.4]
  assign wdata_io_out_ready = io_dram_wdata_ready; // @[StreamController.scala 98:22:@46981.4]
  assign wresp_clock = clock; // @[:@46983.4]
  assign wresp_reset = reset; // @[:@46984.4]
  assign wresp_io_in_valid = io_dram_wresp_valid; // @[StreamController.scala 102:21:@47247.4]
  assign wresp_io_in_bits = 1'h1; // @[StreamController.scala 103:20:@47248.4]
  assign wresp_io_out_ready = io_store_wresp_ready; // @[StreamController.scala 108:22:@47252.4]
  assign wresp_io_banks_0_wdata_valid = 1'h0;
  assign wresp_io_banks_0_wdata_bits = 1'h0;
  assign wresp_io_banks_1_wdata_valid = 1'h0;
  assign wresp_io_banks_1_wdata_bits = 1'h0;
  assign wresp_io_banks_2_wdata_valid = 1'h0;
  assign wresp_io_banks_2_wdata_bits = 1'h0;
  assign wresp_io_banks_3_wdata_valid = 1'h0;
  assign wresp_io_banks_3_wdata_bits = 1'h0;
  assign wresp_io_banks_4_wdata_valid = 1'h0;
  assign wresp_io_banks_4_wdata_bits = 1'h0;
  assign wresp_io_banks_5_wdata_valid = 1'h0;
  assign wresp_io_banks_5_wdata_bits = 1'h0;
  assign wresp_io_banks_6_wdata_valid = 1'h0;
  assign wresp_io_banks_6_wdata_bits = 1'h0;
  assign wresp_io_banks_7_wdata_valid = 1'h0;
  assign wresp_io_banks_7_wdata_bits = 1'h0;
  assign wresp_io_banks_8_wdata_valid = 1'h0;
  assign wresp_io_banks_8_wdata_bits = 1'h0;
  assign wresp_io_banks_9_wdata_valid = 1'h0;
  assign wresp_io_banks_9_wdata_bits = 1'h0;
  assign wresp_io_banks_10_wdata_valid = 1'h0;
  assign wresp_io_banks_10_wdata_bits = 1'h0;
  assign wresp_io_banks_11_wdata_valid = 1'h0;
  assign wresp_io_banks_11_wdata_bits = 1'h0;
  assign wresp_io_banks_12_wdata_valid = 1'h0;
  assign wresp_io_banks_12_wdata_bits = 1'h0;
  assign wresp_io_banks_13_wdata_valid = 1'h0;
  assign wresp_io_banks_13_wdata_bits = 1'h0;
  assign wresp_io_banks_14_wdata_valid = 1'h0;
  assign wresp_io_banks_14_wdata_bits = 1'h0;
  assign wresp_io_banks_15_wdata_valid = 1'h0;
  assign wresp_io_banks_15_wdata_bits = 1'h0;
  assign wresp_io_banks_16_wdata_valid = 1'h0;
  assign wresp_io_banks_16_wdata_bits = 1'h0;
  assign wresp_io_banks_17_wdata_valid = 1'h0;
  assign wresp_io_banks_17_wdata_bits = 1'h0;
  assign wresp_io_banks_18_wdata_valid = 1'h0;
  assign wresp_io_banks_18_wdata_bits = 1'h0;
  assign wresp_io_banks_19_wdata_valid = 1'h0;
  assign wresp_io_banks_19_wdata_bits = 1'h0;
  assign wresp_io_banks_20_wdata_valid = 1'h0;
  assign wresp_io_banks_20_wdata_bits = 1'h0;
  assign wresp_io_banks_21_wdata_valid = 1'h0;
  assign wresp_io_banks_21_wdata_bits = 1'h0;
  assign wresp_io_banks_22_wdata_valid = 1'h0;
  assign wresp_io_banks_22_wdata_bits = 1'h0;
  assign wresp_io_banks_23_wdata_valid = 1'h0;
  assign wresp_io_banks_23_wdata_bits = 1'h0;
  assign wresp_io_banks_24_wdata_valid = 1'h0;
  assign wresp_io_banks_24_wdata_bits = 1'h0;
  assign wresp_io_banks_25_wdata_valid = 1'h0;
  assign wresp_io_banks_25_wdata_bits = 1'h0;
  assign wresp_io_banks_26_wdata_valid = 1'h0;
  assign wresp_io_banks_26_wdata_bits = 1'h0;
  assign wresp_io_banks_27_wdata_valid = 1'h0;
  assign wresp_io_banks_27_wdata_bits = 1'h0;
  assign wresp_io_banks_28_wdata_valid = 1'h0;
  assign wresp_io_banks_28_wdata_bits = 1'h0;
  assign wresp_io_banks_29_wdata_valid = 1'h0;
  assign wresp_io_banks_29_wdata_bits = 1'h0;
  assign wresp_io_banks_30_wdata_valid = 1'h0;
  assign wresp_io_banks_30_wdata_bits = 1'h0;
  assign wresp_io_banks_31_wdata_valid = 1'h0;
  assign wresp_io_banks_31_wdata_bits = 1'h0;
  assign wresp_io_banks_32_wdata_valid = 1'h0;
  assign wresp_io_banks_32_wdata_bits = 1'h0;
  assign wresp_io_banks_33_wdata_valid = 1'h0;
  assign wresp_io_banks_33_wdata_bits = 1'h0;
  assign wresp_io_banks_34_wdata_valid = 1'h0;
  assign wresp_io_banks_34_wdata_bits = 1'h0;
  assign wresp_io_banks_35_wdata_valid = 1'h0;
  assign wresp_io_banks_35_wdata_bits = 1'h0;
  assign wresp_io_banks_36_wdata_valid = 1'h0;
  assign wresp_io_banks_36_wdata_bits = 1'h0;
  assign wresp_io_banks_37_wdata_valid = 1'h0;
  assign wresp_io_banks_37_wdata_bits = 1'h0;
  assign wresp_io_banks_38_wdata_valid = 1'h0;
  assign wresp_io_banks_38_wdata_bits = 1'h0;
  assign wresp_io_banks_39_wdata_valid = 1'h0;
  assign wresp_io_banks_39_wdata_bits = 1'h0;
  assign wresp_io_banks_40_wdata_valid = 1'h0;
  assign wresp_io_banks_40_wdata_bits = 1'h0;
  assign wresp_io_banks_41_wdata_valid = 1'h0;
  assign wresp_io_banks_41_wdata_bits = 1'h0;
  assign wresp_io_banks_42_wdata_valid = 1'h0;
  assign wresp_io_banks_42_wdata_bits = 1'h0;
  assign wresp_io_banks_43_wdata_valid = 1'h0;
  assign wresp_io_banks_43_wdata_bits = 1'h0;
  assign wresp_io_banks_44_wdata_valid = 1'h0;
  assign wresp_io_banks_44_wdata_bits = 1'h0;
  assign wresp_io_banks_45_wdata_valid = 1'h0;
  assign wresp_io_banks_45_wdata_bits = 1'h0;
  assign wresp_io_banks_46_wdata_valid = 1'h0;
  assign wresp_io_banks_46_wdata_bits = 1'h0;
  assign wresp_io_banks_47_wdata_valid = 1'h0;
  assign wresp_io_banks_47_wdata_bits = 1'h0;
  assign wresp_io_banks_48_wdata_valid = 1'h0;
  assign wresp_io_banks_48_wdata_bits = 1'h0;
  assign wresp_io_banks_49_wdata_valid = 1'h0;
  assign wresp_io_banks_49_wdata_bits = 1'h0;
  assign wresp_io_banks_50_wdata_valid = 1'h0;
  assign wresp_io_banks_50_wdata_bits = 1'h0;
  assign wresp_io_banks_51_wdata_valid = 1'h0;
  assign wresp_io_banks_51_wdata_bits = 1'h0;
  assign wresp_io_banks_52_wdata_valid = 1'h0;
  assign wresp_io_banks_52_wdata_bits = 1'h0;
  assign wresp_io_banks_53_wdata_valid = 1'h0;
  assign wresp_io_banks_53_wdata_bits = 1'h0;
  assign wresp_io_banks_54_wdata_valid = 1'h0;
  assign wresp_io_banks_54_wdata_bits = 1'h0;
  assign wresp_io_banks_55_wdata_valid = 1'h0;
  assign wresp_io_banks_55_wdata_bits = 1'h0;
  assign wresp_io_banks_56_wdata_valid = 1'h0;
  assign wresp_io_banks_56_wdata_bits = 1'h0;
  assign wresp_io_banks_57_wdata_valid = 1'h0;
  assign wresp_io_banks_57_wdata_bits = 1'h0;
  assign wresp_io_banks_58_wdata_valid = 1'h0;
  assign wresp_io_banks_58_wdata_bits = 1'h0;
  assign wresp_io_banks_59_wdata_valid = 1'h0;
  assign wresp_io_banks_59_wdata_bits = 1'h0;
  assign wresp_io_banks_60_wdata_valid = 1'h0;
  assign wresp_io_banks_60_wdata_bits = 1'h0;
  assign wresp_io_banks_61_wdata_valid = 1'h0;
  assign wresp_io_banks_61_wdata_bits = 1'h0;
  assign wresp_io_banks_62_wdata_valid = 1'h0;
  assign wresp_io_banks_62_wdata_bits = 1'h0;
  assign wresp_io_banks_63_wdata_valid = 1'h0;
  assign wresp_io_banks_63_wdata_bits = 1'h0;
endmodule
module MuxPipe( // @[:@47318.2]
  output        io_in_ready, // @[:@47321.4]
  input         io_in_valid, // @[:@47321.4]
  input  [63:0] io_in_bits_0_addr, // @[:@47321.4]
  input  [31:0] io_in_bits_0_size, // @[:@47321.4]
  input         io_in_bits_0_isWr, // @[:@47321.4]
  input  [31:0] io_in_bits_0_tag, // @[:@47321.4]
  input         io_out_ready, // @[:@47321.4]
  output        io_out_valid, // @[:@47321.4]
  output [63:0] io_out_bits_addr, // @[:@47321.4]
  output [31:0] io_out_bits_size, // @[:@47321.4]
  output        io_out_bits_isWr, // @[:@47321.4]
  output [31:0] io_out_bits_tag // @[:@47321.4]
);
  wire  _T_42; // @[MuxN.scala 28:31:@47323.4]
  assign _T_42 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@47323.4]
  assign io_in_ready = io_out_ready | _T_42; // @[MuxN.scala 71:15:@47332.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@47331.4]
  assign io_out_bits_addr = io_in_bits_0_addr; // @[MuxN.scala 72:15:@47337.4]
  assign io_out_bits_size = io_in_bits_0_size; // @[MuxN.scala 72:15:@47336.4]
  assign io_out_bits_isWr = io_in_bits_0_isWr; // @[MuxN.scala 72:15:@47334.4]
  assign io_out_bits_tag = io_in_bits_0_tag; // @[MuxN.scala 72:15:@47333.4]
endmodule
module MuxPipe_1( // @[:@47339.2]
  output        io_in_ready, // @[:@47342.4]
  input         io_in_valid, // @[:@47342.4]
  input  [31:0] io_in_bits_0_wdata_0, // @[:@47342.4]
  input  [31:0] io_in_bits_0_wdata_1, // @[:@47342.4]
  input  [31:0] io_in_bits_0_wdata_2, // @[:@47342.4]
  input  [31:0] io_in_bits_0_wdata_3, // @[:@47342.4]
  input  [31:0] io_in_bits_0_wdata_4, // @[:@47342.4]
  input  [31:0] io_in_bits_0_wdata_5, // @[:@47342.4]
  input  [31:0] io_in_bits_0_wdata_6, // @[:@47342.4]
  input  [31:0] io_in_bits_0_wdata_7, // @[:@47342.4]
  input  [31:0] io_in_bits_0_wdata_8, // @[:@47342.4]
  input  [31:0] io_in_bits_0_wdata_9, // @[:@47342.4]
  input  [31:0] io_in_bits_0_wdata_10, // @[:@47342.4]
  input  [31:0] io_in_bits_0_wdata_11, // @[:@47342.4]
  input  [31:0] io_in_bits_0_wdata_12, // @[:@47342.4]
  input  [31:0] io_in_bits_0_wdata_13, // @[:@47342.4]
  input  [31:0] io_in_bits_0_wdata_14, // @[:@47342.4]
  input  [31:0] io_in_bits_0_wdata_15, // @[:@47342.4]
  input         io_in_bits_0_wstrb_0, // @[:@47342.4]
  input         io_in_bits_0_wstrb_1, // @[:@47342.4]
  input         io_in_bits_0_wstrb_2, // @[:@47342.4]
  input         io_in_bits_0_wstrb_3, // @[:@47342.4]
  input         io_in_bits_0_wstrb_4, // @[:@47342.4]
  input         io_in_bits_0_wstrb_5, // @[:@47342.4]
  input         io_in_bits_0_wstrb_6, // @[:@47342.4]
  input         io_in_bits_0_wstrb_7, // @[:@47342.4]
  input         io_in_bits_0_wstrb_8, // @[:@47342.4]
  input         io_in_bits_0_wstrb_9, // @[:@47342.4]
  input         io_in_bits_0_wstrb_10, // @[:@47342.4]
  input         io_in_bits_0_wstrb_11, // @[:@47342.4]
  input         io_in_bits_0_wstrb_12, // @[:@47342.4]
  input         io_in_bits_0_wstrb_13, // @[:@47342.4]
  input         io_in_bits_0_wstrb_14, // @[:@47342.4]
  input         io_in_bits_0_wstrb_15, // @[:@47342.4]
  input         io_in_bits_0_wstrb_16, // @[:@47342.4]
  input         io_in_bits_0_wstrb_17, // @[:@47342.4]
  input         io_in_bits_0_wstrb_18, // @[:@47342.4]
  input         io_in_bits_0_wstrb_19, // @[:@47342.4]
  input         io_in_bits_0_wstrb_20, // @[:@47342.4]
  input         io_in_bits_0_wstrb_21, // @[:@47342.4]
  input         io_in_bits_0_wstrb_22, // @[:@47342.4]
  input         io_in_bits_0_wstrb_23, // @[:@47342.4]
  input         io_in_bits_0_wstrb_24, // @[:@47342.4]
  input         io_in_bits_0_wstrb_25, // @[:@47342.4]
  input         io_in_bits_0_wstrb_26, // @[:@47342.4]
  input         io_in_bits_0_wstrb_27, // @[:@47342.4]
  input         io_in_bits_0_wstrb_28, // @[:@47342.4]
  input         io_in_bits_0_wstrb_29, // @[:@47342.4]
  input         io_in_bits_0_wstrb_30, // @[:@47342.4]
  input         io_in_bits_0_wstrb_31, // @[:@47342.4]
  input         io_in_bits_0_wstrb_32, // @[:@47342.4]
  input         io_in_bits_0_wstrb_33, // @[:@47342.4]
  input         io_in_bits_0_wstrb_34, // @[:@47342.4]
  input         io_in_bits_0_wstrb_35, // @[:@47342.4]
  input         io_in_bits_0_wstrb_36, // @[:@47342.4]
  input         io_in_bits_0_wstrb_37, // @[:@47342.4]
  input         io_in_bits_0_wstrb_38, // @[:@47342.4]
  input         io_in_bits_0_wstrb_39, // @[:@47342.4]
  input         io_in_bits_0_wstrb_40, // @[:@47342.4]
  input         io_in_bits_0_wstrb_41, // @[:@47342.4]
  input         io_in_bits_0_wstrb_42, // @[:@47342.4]
  input         io_in_bits_0_wstrb_43, // @[:@47342.4]
  input         io_in_bits_0_wstrb_44, // @[:@47342.4]
  input         io_in_bits_0_wstrb_45, // @[:@47342.4]
  input         io_in_bits_0_wstrb_46, // @[:@47342.4]
  input         io_in_bits_0_wstrb_47, // @[:@47342.4]
  input         io_in_bits_0_wstrb_48, // @[:@47342.4]
  input         io_in_bits_0_wstrb_49, // @[:@47342.4]
  input         io_in_bits_0_wstrb_50, // @[:@47342.4]
  input         io_in_bits_0_wstrb_51, // @[:@47342.4]
  input         io_in_bits_0_wstrb_52, // @[:@47342.4]
  input         io_in_bits_0_wstrb_53, // @[:@47342.4]
  input         io_in_bits_0_wstrb_54, // @[:@47342.4]
  input         io_in_bits_0_wstrb_55, // @[:@47342.4]
  input         io_in_bits_0_wstrb_56, // @[:@47342.4]
  input         io_in_bits_0_wstrb_57, // @[:@47342.4]
  input         io_in_bits_0_wstrb_58, // @[:@47342.4]
  input         io_in_bits_0_wstrb_59, // @[:@47342.4]
  input         io_in_bits_0_wstrb_60, // @[:@47342.4]
  input         io_in_bits_0_wstrb_61, // @[:@47342.4]
  input         io_in_bits_0_wstrb_62, // @[:@47342.4]
  input         io_in_bits_0_wstrb_63, // @[:@47342.4]
  input         io_out_ready, // @[:@47342.4]
  output        io_out_valid, // @[:@47342.4]
  output [31:0] io_out_bits_wdata_0, // @[:@47342.4]
  output [31:0] io_out_bits_wdata_1, // @[:@47342.4]
  output [31:0] io_out_bits_wdata_2, // @[:@47342.4]
  output [31:0] io_out_bits_wdata_3, // @[:@47342.4]
  output [31:0] io_out_bits_wdata_4, // @[:@47342.4]
  output [31:0] io_out_bits_wdata_5, // @[:@47342.4]
  output [31:0] io_out_bits_wdata_6, // @[:@47342.4]
  output [31:0] io_out_bits_wdata_7, // @[:@47342.4]
  output [31:0] io_out_bits_wdata_8, // @[:@47342.4]
  output [31:0] io_out_bits_wdata_9, // @[:@47342.4]
  output [31:0] io_out_bits_wdata_10, // @[:@47342.4]
  output [31:0] io_out_bits_wdata_11, // @[:@47342.4]
  output [31:0] io_out_bits_wdata_12, // @[:@47342.4]
  output [31:0] io_out_bits_wdata_13, // @[:@47342.4]
  output [31:0] io_out_bits_wdata_14, // @[:@47342.4]
  output [31:0] io_out_bits_wdata_15, // @[:@47342.4]
  output        io_out_bits_wstrb_0, // @[:@47342.4]
  output        io_out_bits_wstrb_1, // @[:@47342.4]
  output        io_out_bits_wstrb_2, // @[:@47342.4]
  output        io_out_bits_wstrb_3, // @[:@47342.4]
  output        io_out_bits_wstrb_4, // @[:@47342.4]
  output        io_out_bits_wstrb_5, // @[:@47342.4]
  output        io_out_bits_wstrb_6, // @[:@47342.4]
  output        io_out_bits_wstrb_7, // @[:@47342.4]
  output        io_out_bits_wstrb_8, // @[:@47342.4]
  output        io_out_bits_wstrb_9, // @[:@47342.4]
  output        io_out_bits_wstrb_10, // @[:@47342.4]
  output        io_out_bits_wstrb_11, // @[:@47342.4]
  output        io_out_bits_wstrb_12, // @[:@47342.4]
  output        io_out_bits_wstrb_13, // @[:@47342.4]
  output        io_out_bits_wstrb_14, // @[:@47342.4]
  output        io_out_bits_wstrb_15, // @[:@47342.4]
  output        io_out_bits_wstrb_16, // @[:@47342.4]
  output        io_out_bits_wstrb_17, // @[:@47342.4]
  output        io_out_bits_wstrb_18, // @[:@47342.4]
  output        io_out_bits_wstrb_19, // @[:@47342.4]
  output        io_out_bits_wstrb_20, // @[:@47342.4]
  output        io_out_bits_wstrb_21, // @[:@47342.4]
  output        io_out_bits_wstrb_22, // @[:@47342.4]
  output        io_out_bits_wstrb_23, // @[:@47342.4]
  output        io_out_bits_wstrb_24, // @[:@47342.4]
  output        io_out_bits_wstrb_25, // @[:@47342.4]
  output        io_out_bits_wstrb_26, // @[:@47342.4]
  output        io_out_bits_wstrb_27, // @[:@47342.4]
  output        io_out_bits_wstrb_28, // @[:@47342.4]
  output        io_out_bits_wstrb_29, // @[:@47342.4]
  output        io_out_bits_wstrb_30, // @[:@47342.4]
  output        io_out_bits_wstrb_31, // @[:@47342.4]
  output        io_out_bits_wstrb_32, // @[:@47342.4]
  output        io_out_bits_wstrb_33, // @[:@47342.4]
  output        io_out_bits_wstrb_34, // @[:@47342.4]
  output        io_out_bits_wstrb_35, // @[:@47342.4]
  output        io_out_bits_wstrb_36, // @[:@47342.4]
  output        io_out_bits_wstrb_37, // @[:@47342.4]
  output        io_out_bits_wstrb_38, // @[:@47342.4]
  output        io_out_bits_wstrb_39, // @[:@47342.4]
  output        io_out_bits_wstrb_40, // @[:@47342.4]
  output        io_out_bits_wstrb_41, // @[:@47342.4]
  output        io_out_bits_wstrb_42, // @[:@47342.4]
  output        io_out_bits_wstrb_43, // @[:@47342.4]
  output        io_out_bits_wstrb_44, // @[:@47342.4]
  output        io_out_bits_wstrb_45, // @[:@47342.4]
  output        io_out_bits_wstrb_46, // @[:@47342.4]
  output        io_out_bits_wstrb_47, // @[:@47342.4]
  output        io_out_bits_wstrb_48, // @[:@47342.4]
  output        io_out_bits_wstrb_49, // @[:@47342.4]
  output        io_out_bits_wstrb_50, // @[:@47342.4]
  output        io_out_bits_wstrb_51, // @[:@47342.4]
  output        io_out_bits_wstrb_52, // @[:@47342.4]
  output        io_out_bits_wstrb_53, // @[:@47342.4]
  output        io_out_bits_wstrb_54, // @[:@47342.4]
  output        io_out_bits_wstrb_55, // @[:@47342.4]
  output        io_out_bits_wstrb_56, // @[:@47342.4]
  output        io_out_bits_wstrb_57, // @[:@47342.4]
  output        io_out_bits_wstrb_58, // @[:@47342.4]
  output        io_out_bits_wstrb_59, // @[:@47342.4]
  output        io_out_bits_wstrb_60, // @[:@47342.4]
  output        io_out_bits_wstrb_61, // @[:@47342.4]
  output        io_out_bits_wstrb_62, // @[:@47342.4]
  output        io_out_bits_wstrb_63 // @[:@47342.4]
);
  wire  _T_146; // @[MuxN.scala 28:31:@47344.4]
  assign _T_146 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@47344.4]
  assign io_in_ready = io_out_ready | _T_146; // @[MuxN.scala 71:15:@47429.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@47428.4]
  assign io_out_bits_wdata_0 = io_in_bits_0_wdata_0; // @[MuxN.scala 72:15:@47495.4]
  assign io_out_bits_wdata_1 = io_in_bits_0_wdata_1; // @[MuxN.scala 72:15:@47496.4]
  assign io_out_bits_wdata_2 = io_in_bits_0_wdata_2; // @[MuxN.scala 72:15:@47497.4]
  assign io_out_bits_wdata_3 = io_in_bits_0_wdata_3; // @[MuxN.scala 72:15:@47498.4]
  assign io_out_bits_wdata_4 = io_in_bits_0_wdata_4; // @[MuxN.scala 72:15:@47499.4]
  assign io_out_bits_wdata_5 = io_in_bits_0_wdata_5; // @[MuxN.scala 72:15:@47500.4]
  assign io_out_bits_wdata_6 = io_in_bits_0_wdata_6; // @[MuxN.scala 72:15:@47501.4]
  assign io_out_bits_wdata_7 = io_in_bits_0_wdata_7; // @[MuxN.scala 72:15:@47502.4]
  assign io_out_bits_wdata_8 = io_in_bits_0_wdata_8; // @[MuxN.scala 72:15:@47503.4]
  assign io_out_bits_wdata_9 = io_in_bits_0_wdata_9; // @[MuxN.scala 72:15:@47504.4]
  assign io_out_bits_wdata_10 = io_in_bits_0_wdata_10; // @[MuxN.scala 72:15:@47505.4]
  assign io_out_bits_wdata_11 = io_in_bits_0_wdata_11; // @[MuxN.scala 72:15:@47506.4]
  assign io_out_bits_wdata_12 = io_in_bits_0_wdata_12; // @[MuxN.scala 72:15:@47507.4]
  assign io_out_bits_wdata_13 = io_in_bits_0_wdata_13; // @[MuxN.scala 72:15:@47508.4]
  assign io_out_bits_wdata_14 = io_in_bits_0_wdata_14; // @[MuxN.scala 72:15:@47509.4]
  assign io_out_bits_wdata_15 = io_in_bits_0_wdata_15; // @[MuxN.scala 72:15:@47510.4]
  assign io_out_bits_wstrb_0 = io_in_bits_0_wstrb_0; // @[MuxN.scala 72:15:@47431.4]
  assign io_out_bits_wstrb_1 = io_in_bits_0_wstrb_1; // @[MuxN.scala 72:15:@47432.4]
  assign io_out_bits_wstrb_2 = io_in_bits_0_wstrb_2; // @[MuxN.scala 72:15:@47433.4]
  assign io_out_bits_wstrb_3 = io_in_bits_0_wstrb_3; // @[MuxN.scala 72:15:@47434.4]
  assign io_out_bits_wstrb_4 = io_in_bits_0_wstrb_4; // @[MuxN.scala 72:15:@47435.4]
  assign io_out_bits_wstrb_5 = io_in_bits_0_wstrb_5; // @[MuxN.scala 72:15:@47436.4]
  assign io_out_bits_wstrb_6 = io_in_bits_0_wstrb_6; // @[MuxN.scala 72:15:@47437.4]
  assign io_out_bits_wstrb_7 = io_in_bits_0_wstrb_7; // @[MuxN.scala 72:15:@47438.4]
  assign io_out_bits_wstrb_8 = io_in_bits_0_wstrb_8; // @[MuxN.scala 72:15:@47439.4]
  assign io_out_bits_wstrb_9 = io_in_bits_0_wstrb_9; // @[MuxN.scala 72:15:@47440.4]
  assign io_out_bits_wstrb_10 = io_in_bits_0_wstrb_10; // @[MuxN.scala 72:15:@47441.4]
  assign io_out_bits_wstrb_11 = io_in_bits_0_wstrb_11; // @[MuxN.scala 72:15:@47442.4]
  assign io_out_bits_wstrb_12 = io_in_bits_0_wstrb_12; // @[MuxN.scala 72:15:@47443.4]
  assign io_out_bits_wstrb_13 = io_in_bits_0_wstrb_13; // @[MuxN.scala 72:15:@47444.4]
  assign io_out_bits_wstrb_14 = io_in_bits_0_wstrb_14; // @[MuxN.scala 72:15:@47445.4]
  assign io_out_bits_wstrb_15 = io_in_bits_0_wstrb_15; // @[MuxN.scala 72:15:@47446.4]
  assign io_out_bits_wstrb_16 = io_in_bits_0_wstrb_16; // @[MuxN.scala 72:15:@47447.4]
  assign io_out_bits_wstrb_17 = io_in_bits_0_wstrb_17; // @[MuxN.scala 72:15:@47448.4]
  assign io_out_bits_wstrb_18 = io_in_bits_0_wstrb_18; // @[MuxN.scala 72:15:@47449.4]
  assign io_out_bits_wstrb_19 = io_in_bits_0_wstrb_19; // @[MuxN.scala 72:15:@47450.4]
  assign io_out_bits_wstrb_20 = io_in_bits_0_wstrb_20; // @[MuxN.scala 72:15:@47451.4]
  assign io_out_bits_wstrb_21 = io_in_bits_0_wstrb_21; // @[MuxN.scala 72:15:@47452.4]
  assign io_out_bits_wstrb_22 = io_in_bits_0_wstrb_22; // @[MuxN.scala 72:15:@47453.4]
  assign io_out_bits_wstrb_23 = io_in_bits_0_wstrb_23; // @[MuxN.scala 72:15:@47454.4]
  assign io_out_bits_wstrb_24 = io_in_bits_0_wstrb_24; // @[MuxN.scala 72:15:@47455.4]
  assign io_out_bits_wstrb_25 = io_in_bits_0_wstrb_25; // @[MuxN.scala 72:15:@47456.4]
  assign io_out_bits_wstrb_26 = io_in_bits_0_wstrb_26; // @[MuxN.scala 72:15:@47457.4]
  assign io_out_bits_wstrb_27 = io_in_bits_0_wstrb_27; // @[MuxN.scala 72:15:@47458.4]
  assign io_out_bits_wstrb_28 = io_in_bits_0_wstrb_28; // @[MuxN.scala 72:15:@47459.4]
  assign io_out_bits_wstrb_29 = io_in_bits_0_wstrb_29; // @[MuxN.scala 72:15:@47460.4]
  assign io_out_bits_wstrb_30 = io_in_bits_0_wstrb_30; // @[MuxN.scala 72:15:@47461.4]
  assign io_out_bits_wstrb_31 = io_in_bits_0_wstrb_31; // @[MuxN.scala 72:15:@47462.4]
  assign io_out_bits_wstrb_32 = io_in_bits_0_wstrb_32; // @[MuxN.scala 72:15:@47463.4]
  assign io_out_bits_wstrb_33 = io_in_bits_0_wstrb_33; // @[MuxN.scala 72:15:@47464.4]
  assign io_out_bits_wstrb_34 = io_in_bits_0_wstrb_34; // @[MuxN.scala 72:15:@47465.4]
  assign io_out_bits_wstrb_35 = io_in_bits_0_wstrb_35; // @[MuxN.scala 72:15:@47466.4]
  assign io_out_bits_wstrb_36 = io_in_bits_0_wstrb_36; // @[MuxN.scala 72:15:@47467.4]
  assign io_out_bits_wstrb_37 = io_in_bits_0_wstrb_37; // @[MuxN.scala 72:15:@47468.4]
  assign io_out_bits_wstrb_38 = io_in_bits_0_wstrb_38; // @[MuxN.scala 72:15:@47469.4]
  assign io_out_bits_wstrb_39 = io_in_bits_0_wstrb_39; // @[MuxN.scala 72:15:@47470.4]
  assign io_out_bits_wstrb_40 = io_in_bits_0_wstrb_40; // @[MuxN.scala 72:15:@47471.4]
  assign io_out_bits_wstrb_41 = io_in_bits_0_wstrb_41; // @[MuxN.scala 72:15:@47472.4]
  assign io_out_bits_wstrb_42 = io_in_bits_0_wstrb_42; // @[MuxN.scala 72:15:@47473.4]
  assign io_out_bits_wstrb_43 = io_in_bits_0_wstrb_43; // @[MuxN.scala 72:15:@47474.4]
  assign io_out_bits_wstrb_44 = io_in_bits_0_wstrb_44; // @[MuxN.scala 72:15:@47475.4]
  assign io_out_bits_wstrb_45 = io_in_bits_0_wstrb_45; // @[MuxN.scala 72:15:@47476.4]
  assign io_out_bits_wstrb_46 = io_in_bits_0_wstrb_46; // @[MuxN.scala 72:15:@47477.4]
  assign io_out_bits_wstrb_47 = io_in_bits_0_wstrb_47; // @[MuxN.scala 72:15:@47478.4]
  assign io_out_bits_wstrb_48 = io_in_bits_0_wstrb_48; // @[MuxN.scala 72:15:@47479.4]
  assign io_out_bits_wstrb_49 = io_in_bits_0_wstrb_49; // @[MuxN.scala 72:15:@47480.4]
  assign io_out_bits_wstrb_50 = io_in_bits_0_wstrb_50; // @[MuxN.scala 72:15:@47481.4]
  assign io_out_bits_wstrb_51 = io_in_bits_0_wstrb_51; // @[MuxN.scala 72:15:@47482.4]
  assign io_out_bits_wstrb_52 = io_in_bits_0_wstrb_52; // @[MuxN.scala 72:15:@47483.4]
  assign io_out_bits_wstrb_53 = io_in_bits_0_wstrb_53; // @[MuxN.scala 72:15:@47484.4]
  assign io_out_bits_wstrb_54 = io_in_bits_0_wstrb_54; // @[MuxN.scala 72:15:@47485.4]
  assign io_out_bits_wstrb_55 = io_in_bits_0_wstrb_55; // @[MuxN.scala 72:15:@47486.4]
  assign io_out_bits_wstrb_56 = io_in_bits_0_wstrb_56; // @[MuxN.scala 72:15:@47487.4]
  assign io_out_bits_wstrb_57 = io_in_bits_0_wstrb_57; // @[MuxN.scala 72:15:@47488.4]
  assign io_out_bits_wstrb_58 = io_in_bits_0_wstrb_58; // @[MuxN.scala 72:15:@47489.4]
  assign io_out_bits_wstrb_59 = io_in_bits_0_wstrb_59; // @[MuxN.scala 72:15:@47490.4]
  assign io_out_bits_wstrb_60 = io_in_bits_0_wstrb_60; // @[MuxN.scala 72:15:@47491.4]
  assign io_out_bits_wstrb_61 = io_in_bits_0_wstrb_61; // @[MuxN.scala 72:15:@47492.4]
  assign io_out_bits_wstrb_62 = io_in_bits_0_wstrb_62; // @[MuxN.scala 72:15:@47493.4]
  assign io_out_bits_wstrb_63 = io_in_bits_0_wstrb_63; // @[MuxN.scala 72:15:@47494.4]
endmodule
module ElementCounter( // @[:@47512.2]
  input         clock, // @[:@47513.4]
  input         reset, // @[:@47514.4]
  input         io_reset, // @[:@47515.4]
  input         io_enable, // @[:@47515.4]
  output [31:0] io_out // @[:@47515.4]
);
  reg [31:0] count; // @[Counter.scala 37:22:@47517.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_14; // @[Counter.scala 39:24:@47518.4]
  wire [31:0] newCount; // @[Counter.scala 39:24:@47519.4]
  wire [31:0] _GEN_0; // @[Counter.scala 43:26:@47524.6]
  wire [31:0] _GEN_1; // @[Counter.scala 41:18:@47520.4]
  assign _T_14 = count + 32'h1; // @[Counter.scala 39:24:@47518.4]
  assign newCount = count + 32'h1; // @[Counter.scala 39:24:@47519.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 43:26:@47524.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 41:18:@47520.4]
  assign io_out = count; // @[Counter.scala 47:10:@47527.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module StreamArbiter( // @[:@47529.2]
  input         clock, // @[:@47530.4]
  input         reset, // @[:@47531.4]
  output        io_app_0_cmd_ready, // @[:@47532.4]
  input         io_app_0_cmd_valid, // @[:@47532.4]
  input  [63:0] io_app_0_cmd_bits_addr, // @[:@47532.4]
  input  [31:0] io_app_0_cmd_bits_size, // @[:@47532.4]
  input         io_app_0_cmd_bits_isWr, // @[:@47532.4]
  input  [31:0] io_app_0_cmd_bits_tag, // @[:@47532.4]
  output        io_app_0_wdata_ready, // @[:@47532.4]
  input         io_app_0_wdata_valid, // @[:@47532.4]
  input  [31:0] io_app_0_wdata_bits_wdata_0, // @[:@47532.4]
  input  [31:0] io_app_0_wdata_bits_wdata_1, // @[:@47532.4]
  input  [31:0] io_app_0_wdata_bits_wdata_2, // @[:@47532.4]
  input  [31:0] io_app_0_wdata_bits_wdata_3, // @[:@47532.4]
  input  [31:0] io_app_0_wdata_bits_wdata_4, // @[:@47532.4]
  input  [31:0] io_app_0_wdata_bits_wdata_5, // @[:@47532.4]
  input  [31:0] io_app_0_wdata_bits_wdata_6, // @[:@47532.4]
  input  [31:0] io_app_0_wdata_bits_wdata_7, // @[:@47532.4]
  input  [31:0] io_app_0_wdata_bits_wdata_8, // @[:@47532.4]
  input  [31:0] io_app_0_wdata_bits_wdata_9, // @[:@47532.4]
  input  [31:0] io_app_0_wdata_bits_wdata_10, // @[:@47532.4]
  input  [31:0] io_app_0_wdata_bits_wdata_11, // @[:@47532.4]
  input  [31:0] io_app_0_wdata_bits_wdata_12, // @[:@47532.4]
  input  [31:0] io_app_0_wdata_bits_wdata_13, // @[:@47532.4]
  input  [31:0] io_app_0_wdata_bits_wdata_14, // @[:@47532.4]
  input  [31:0] io_app_0_wdata_bits_wdata_15, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_0, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_1, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_2, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_3, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_4, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_5, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_6, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_7, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_8, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_9, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_10, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_11, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_12, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_13, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_14, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_15, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_16, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_17, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_18, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_19, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_20, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_21, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_22, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_23, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_24, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_25, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_26, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_27, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_28, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_29, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_30, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_31, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_32, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_33, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_34, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_35, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_36, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_37, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_38, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_39, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_40, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_41, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_42, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_43, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_44, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_45, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_46, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_47, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_48, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_49, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_50, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_51, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_52, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_53, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_54, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_55, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_56, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_57, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_58, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_59, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_60, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_61, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_62, // @[:@47532.4]
  input         io_app_0_wdata_bits_wstrb_63, // @[:@47532.4]
  input         io_app_0_rresp_ready, // @[:@47532.4]
  input         io_app_0_wresp_ready, // @[:@47532.4]
  output        io_app_0_wresp_valid, // @[:@47532.4]
  input         io_dram_cmd_ready, // @[:@47532.4]
  output        io_dram_cmd_valid, // @[:@47532.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@47532.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@47532.4]
  output        io_dram_cmd_bits_isWr, // @[:@47532.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@47532.4]
  input         io_dram_wdata_ready, // @[:@47532.4]
  output        io_dram_wdata_valid, // @[:@47532.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@47532.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@47532.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@47532.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@47532.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@47532.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@47532.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@47532.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@47532.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@47532.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@47532.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@47532.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@47532.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@47532.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@47532.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@47532.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@47532.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@47532.4]
  output        io_dram_rresp_ready, // @[:@47532.4]
  output        io_dram_wresp_ready, // @[:@47532.4]
  input         io_dram_wresp_valid, // @[:@47532.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@47532.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@47761.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@47761.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@47761.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@47761.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@47761.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@47768.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@47768.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@47768.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@47768.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@47768.4]
  wire  cmdMux_io_in_ready; // @[StreamArbiter.scala 25:22:@47778.4]
  wire  cmdMux_io_in_valid; // @[StreamArbiter.scala 25:22:@47778.4]
  wire [63:0] cmdMux_io_in_bits_0_addr; // @[StreamArbiter.scala 25:22:@47778.4]
  wire [31:0] cmdMux_io_in_bits_0_size; // @[StreamArbiter.scala 25:22:@47778.4]
  wire  cmdMux_io_in_bits_0_isWr; // @[StreamArbiter.scala 25:22:@47778.4]
  wire [31:0] cmdMux_io_in_bits_0_tag; // @[StreamArbiter.scala 25:22:@47778.4]
  wire  cmdMux_io_out_ready; // @[StreamArbiter.scala 25:22:@47778.4]
  wire  cmdMux_io_out_valid; // @[StreamArbiter.scala 25:22:@47778.4]
  wire [63:0] cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 25:22:@47778.4]
  wire [31:0] cmdMux_io_out_bits_size; // @[StreamArbiter.scala 25:22:@47778.4]
  wire  cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 25:22:@47778.4]
  wire [31:0] cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 25:22:@47778.4]
  wire  wdataMux_io_in_ready; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_valid; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_0; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_1; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_2; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_3; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_4; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_5; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_6; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_7; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_8; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_9; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_10; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_11; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_12; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_13; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_14; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_15; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_0; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_1; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_2; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_3; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_4; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_5; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_6; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_7; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_8; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_9; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_10; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_11; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_12; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_13; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_14; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_15; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_16; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_17; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_18; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_19; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_20; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_21; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_22; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_23; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_24; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_25; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_26; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_27; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_28; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_29; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_30; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_31; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_32; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_33; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_34; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_35; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_36; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_37; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_38; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_39; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_40; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_41; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_42; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_43; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_44; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_45; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_46; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_47; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_48; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_49; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_50; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_51; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_52; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_53; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_54; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_55; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_56; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_57; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_58; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_59; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_60; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_61; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_62; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_in_bits_0_wstrb_63; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_ready; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_valid; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 35:24:@47801.4]
  wire [31:0] wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 35:24:@47801.4]
  wire  elementCtr_clock; // @[StreamArbiter.scala 36:26:@47804.4]
  wire  elementCtr_reset; // @[StreamArbiter.scala 36:26:@47804.4]
  wire  elementCtr_io_reset; // @[StreamArbiter.scala 36:26:@47804.4]
  wire  elementCtr_io_enable; // @[StreamArbiter.scala 36:26:@47804.4]
  wire [31:0] elementCtr_io_out; // @[StreamArbiter.scala 36:26:@47804.4]
  wire  _T_346; // @[package.scala 96:25:@47773.4 package.scala 96:25:@47774.4]
  wire  cmdIdx; // @[StreamArbiter.scala 21:16:@47775.4]
  wire [1:0] cmdInDecoder; // @[OneHot.scala 45:35:@47777.4]
  wire  _T_355; // @[FringeBundles.scala 114:28:@47793.4]
  wire [22:0] _T_356; // @[FringeBundles.scala 114:28:@47795.4]
  wire [23:0] _T_358; // @[FringeBundles.scala 115:37:@47798.4]
  wire  _T_360; // @[StreamArbiter.scala 37:49:@47807.4]
  wire [31:0] _T_365; // @[:@47811.4 :@47812.4]
  wire [7:0] _T_366; // @[FringeBundles.scala 114:28:@47813.4]
  wire [255:0] cmdOutDecoder; // @[OneHot.scala 45:35:@47819.4]
  wire  _T_379; // @[StreamArbiter.scala 42:78:@47822.4]
  wire  _T_380; // @[StreamArbiter.scala 42:121:@47823.4]
  wire [7:0] _T_395; // @[FringeBundles.scala 140:28:@48010.4]
  wire [255:0] wrespDecoder; // @[OneHot.scala 45:35:@48017.4]
  wire  _T_400; // @[StreamArbiter.scala 61:55:@48022.4]
  wire  _T_403; // @[StreamArbiter.scala 62:85:@48026.4]
  wire  _T_404; // @[StreamArbiter.scala 62:70:@48027.4]
  wire  _T_409; // @[StreamArbiter.scala 67:58:@48051.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@47761.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@47768.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  MuxPipe cmdMux ( // @[StreamArbiter.scala 25:22:@47778.4]
    .io_in_ready(cmdMux_io_in_ready),
    .io_in_valid(cmdMux_io_in_valid),
    .io_in_bits_0_addr(cmdMux_io_in_bits_0_addr),
    .io_in_bits_0_size(cmdMux_io_in_bits_0_size),
    .io_in_bits_0_isWr(cmdMux_io_in_bits_0_isWr),
    .io_in_bits_0_tag(cmdMux_io_in_bits_0_tag),
    .io_out_ready(cmdMux_io_out_ready),
    .io_out_valid(cmdMux_io_out_valid),
    .io_out_bits_addr(cmdMux_io_out_bits_addr),
    .io_out_bits_size(cmdMux_io_out_bits_size),
    .io_out_bits_isWr(cmdMux_io_out_bits_isWr),
    .io_out_bits_tag(cmdMux_io_out_bits_tag)
  );
  MuxPipe_1 wdataMux ( // @[StreamArbiter.scala 35:24:@47801.4]
    .io_in_ready(wdataMux_io_in_ready),
    .io_in_valid(wdataMux_io_in_valid),
    .io_in_bits_0_wdata_0(wdataMux_io_in_bits_0_wdata_0),
    .io_in_bits_0_wdata_1(wdataMux_io_in_bits_0_wdata_1),
    .io_in_bits_0_wdata_2(wdataMux_io_in_bits_0_wdata_2),
    .io_in_bits_0_wdata_3(wdataMux_io_in_bits_0_wdata_3),
    .io_in_bits_0_wdata_4(wdataMux_io_in_bits_0_wdata_4),
    .io_in_bits_0_wdata_5(wdataMux_io_in_bits_0_wdata_5),
    .io_in_bits_0_wdata_6(wdataMux_io_in_bits_0_wdata_6),
    .io_in_bits_0_wdata_7(wdataMux_io_in_bits_0_wdata_7),
    .io_in_bits_0_wdata_8(wdataMux_io_in_bits_0_wdata_8),
    .io_in_bits_0_wdata_9(wdataMux_io_in_bits_0_wdata_9),
    .io_in_bits_0_wdata_10(wdataMux_io_in_bits_0_wdata_10),
    .io_in_bits_0_wdata_11(wdataMux_io_in_bits_0_wdata_11),
    .io_in_bits_0_wdata_12(wdataMux_io_in_bits_0_wdata_12),
    .io_in_bits_0_wdata_13(wdataMux_io_in_bits_0_wdata_13),
    .io_in_bits_0_wdata_14(wdataMux_io_in_bits_0_wdata_14),
    .io_in_bits_0_wdata_15(wdataMux_io_in_bits_0_wdata_15),
    .io_in_bits_0_wstrb_0(wdataMux_io_in_bits_0_wstrb_0),
    .io_in_bits_0_wstrb_1(wdataMux_io_in_bits_0_wstrb_1),
    .io_in_bits_0_wstrb_2(wdataMux_io_in_bits_0_wstrb_2),
    .io_in_bits_0_wstrb_3(wdataMux_io_in_bits_0_wstrb_3),
    .io_in_bits_0_wstrb_4(wdataMux_io_in_bits_0_wstrb_4),
    .io_in_bits_0_wstrb_5(wdataMux_io_in_bits_0_wstrb_5),
    .io_in_bits_0_wstrb_6(wdataMux_io_in_bits_0_wstrb_6),
    .io_in_bits_0_wstrb_7(wdataMux_io_in_bits_0_wstrb_7),
    .io_in_bits_0_wstrb_8(wdataMux_io_in_bits_0_wstrb_8),
    .io_in_bits_0_wstrb_9(wdataMux_io_in_bits_0_wstrb_9),
    .io_in_bits_0_wstrb_10(wdataMux_io_in_bits_0_wstrb_10),
    .io_in_bits_0_wstrb_11(wdataMux_io_in_bits_0_wstrb_11),
    .io_in_bits_0_wstrb_12(wdataMux_io_in_bits_0_wstrb_12),
    .io_in_bits_0_wstrb_13(wdataMux_io_in_bits_0_wstrb_13),
    .io_in_bits_0_wstrb_14(wdataMux_io_in_bits_0_wstrb_14),
    .io_in_bits_0_wstrb_15(wdataMux_io_in_bits_0_wstrb_15),
    .io_in_bits_0_wstrb_16(wdataMux_io_in_bits_0_wstrb_16),
    .io_in_bits_0_wstrb_17(wdataMux_io_in_bits_0_wstrb_17),
    .io_in_bits_0_wstrb_18(wdataMux_io_in_bits_0_wstrb_18),
    .io_in_bits_0_wstrb_19(wdataMux_io_in_bits_0_wstrb_19),
    .io_in_bits_0_wstrb_20(wdataMux_io_in_bits_0_wstrb_20),
    .io_in_bits_0_wstrb_21(wdataMux_io_in_bits_0_wstrb_21),
    .io_in_bits_0_wstrb_22(wdataMux_io_in_bits_0_wstrb_22),
    .io_in_bits_0_wstrb_23(wdataMux_io_in_bits_0_wstrb_23),
    .io_in_bits_0_wstrb_24(wdataMux_io_in_bits_0_wstrb_24),
    .io_in_bits_0_wstrb_25(wdataMux_io_in_bits_0_wstrb_25),
    .io_in_bits_0_wstrb_26(wdataMux_io_in_bits_0_wstrb_26),
    .io_in_bits_0_wstrb_27(wdataMux_io_in_bits_0_wstrb_27),
    .io_in_bits_0_wstrb_28(wdataMux_io_in_bits_0_wstrb_28),
    .io_in_bits_0_wstrb_29(wdataMux_io_in_bits_0_wstrb_29),
    .io_in_bits_0_wstrb_30(wdataMux_io_in_bits_0_wstrb_30),
    .io_in_bits_0_wstrb_31(wdataMux_io_in_bits_0_wstrb_31),
    .io_in_bits_0_wstrb_32(wdataMux_io_in_bits_0_wstrb_32),
    .io_in_bits_0_wstrb_33(wdataMux_io_in_bits_0_wstrb_33),
    .io_in_bits_0_wstrb_34(wdataMux_io_in_bits_0_wstrb_34),
    .io_in_bits_0_wstrb_35(wdataMux_io_in_bits_0_wstrb_35),
    .io_in_bits_0_wstrb_36(wdataMux_io_in_bits_0_wstrb_36),
    .io_in_bits_0_wstrb_37(wdataMux_io_in_bits_0_wstrb_37),
    .io_in_bits_0_wstrb_38(wdataMux_io_in_bits_0_wstrb_38),
    .io_in_bits_0_wstrb_39(wdataMux_io_in_bits_0_wstrb_39),
    .io_in_bits_0_wstrb_40(wdataMux_io_in_bits_0_wstrb_40),
    .io_in_bits_0_wstrb_41(wdataMux_io_in_bits_0_wstrb_41),
    .io_in_bits_0_wstrb_42(wdataMux_io_in_bits_0_wstrb_42),
    .io_in_bits_0_wstrb_43(wdataMux_io_in_bits_0_wstrb_43),
    .io_in_bits_0_wstrb_44(wdataMux_io_in_bits_0_wstrb_44),
    .io_in_bits_0_wstrb_45(wdataMux_io_in_bits_0_wstrb_45),
    .io_in_bits_0_wstrb_46(wdataMux_io_in_bits_0_wstrb_46),
    .io_in_bits_0_wstrb_47(wdataMux_io_in_bits_0_wstrb_47),
    .io_in_bits_0_wstrb_48(wdataMux_io_in_bits_0_wstrb_48),
    .io_in_bits_0_wstrb_49(wdataMux_io_in_bits_0_wstrb_49),
    .io_in_bits_0_wstrb_50(wdataMux_io_in_bits_0_wstrb_50),
    .io_in_bits_0_wstrb_51(wdataMux_io_in_bits_0_wstrb_51),
    .io_in_bits_0_wstrb_52(wdataMux_io_in_bits_0_wstrb_52),
    .io_in_bits_0_wstrb_53(wdataMux_io_in_bits_0_wstrb_53),
    .io_in_bits_0_wstrb_54(wdataMux_io_in_bits_0_wstrb_54),
    .io_in_bits_0_wstrb_55(wdataMux_io_in_bits_0_wstrb_55),
    .io_in_bits_0_wstrb_56(wdataMux_io_in_bits_0_wstrb_56),
    .io_in_bits_0_wstrb_57(wdataMux_io_in_bits_0_wstrb_57),
    .io_in_bits_0_wstrb_58(wdataMux_io_in_bits_0_wstrb_58),
    .io_in_bits_0_wstrb_59(wdataMux_io_in_bits_0_wstrb_59),
    .io_in_bits_0_wstrb_60(wdataMux_io_in_bits_0_wstrb_60),
    .io_in_bits_0_wstrb_61(wdataMux_io_in_bits_0_wstrb_61),
    .io_in_bits_0_wstrb_62(wdataMux_io_in_bits_0_wstrb_62),
    .io_in_bits_0_wstrb_63(wdataMux_io_in_bits_0_wstrb_63),
    .io_out_ready(wdataMux_io_out_ready),
    .io_out_valid(wdataMux_io_out_valid),
    .io_out_bits_wdata_0(wdataMux_io_out_bits_wdata_0),
    .io_out_bits_wdata_1(wdataMux_io_out_bits_wdata_1),
    .io_out_bits_wdata_2(wdataMux_io_out_bits_wdata_2),
    .io_out_bits_wdata_3(wdataMux_io_out_bits_wdata_3),
    .io_out_bits_wdata_4(wdataMux_io_out_bits_wdata_4),
    .io_out_bits_wdata_5(wdataMux_io_out_bits_wdata_5),
    .io_out_bits_wdata_6(wdataMux_io_out_bits_wdata_6),
    .io_out_bits_wdata_7(wdataMux_io_out_bits_wdata_7),
    .io_out_bits_wdata_8(wdataMux_io_out_bits_wdata_8),
    .io_out_bits_wdata_9(wdataMux_io_out_bits_wdata_9),
    .io_out_bits_wdata_10(wdataMux_io_out_bits_wdata_10),
    .io_out_bits_wdata_11(wdataMux_io_out_bits_wdata_11),
    .io_out_bits_wdata_12(wdataMux_io_out_bits_wdata_12),
    .io_out_bits_wdata_13(wdataMux_io_out_bits_wdata_13),
    .io_out_bits_wdata_14(wdataMux_io_out_bits_wdata_14),
    .io_out_bits_wdata_15(wdataMux_io_out_bits_wdata_15),
    .io_out_bits_wstrb_0(wdataMux_io_out_bits_wstrb_0),
    .io_out_bits_wstrb_1(wdataMux_io_out_bits_wstrb_1),
    .io_out_bits_wstrb_2(wdataMux_io_out_bits_wstrb_2),
    .io_out_bits_wstrb_3(wdataMux_io_out_bits_wstrb_3),
    .io_out_bits_wstrb_4(wdataMux_io_out_bits_wstrb_4),
    .io_out_bits_wstrb_5(wdataMux_io_out_bits_wstrb_5),
    .io_out_bits_wstrb_6(wdataMux_io_out_bits_wstrb_6),
    .io_out_bits_wstrb_7(wdataMux_io_out_bits_wstrb_7),
    .io_out_bits_wstrb_8(wdataMux_io_out_bits_wstrb_8),
    .io_out_bits_wstrb_9(wdataMux_io_out_bits_wstrb_9),
    .io_out_bits_wstrb_10(wdataMux_io_out_bits_wstrb_10),
    .io_out_bits_wstrb_11(wdataMux_io_out_bits_wstrb_11),
    .io_out_bits_wstrb_12(wdataMux_io_out_bits_wstrb_12),
    .io_out_bits_wstrb_13(wdataMux_io_out_bits_wstrb_13),
    .io_out_bits_wstrb_14(wdataMux_io_out_bits_wstrb_14),
    .io_out_bits_wstrb_15(wdataMux_io_out_bits_wstrb_15),
    .io_out_bits_wstrb_16(wdataMux_io_out_bits_wstrb_16),
    .io_out_bits_wstrb_17(wdataMux_io_out_bits_wstrb_17),
    .io_out_bits_wstrb_18(wdataMux_io_out_bits_wstrb_18),
    .io_out_bits_wstrb_19(wdataMux_io_out_bits_wstrb_19),
    .io_out_bits_wstrb_20(wdataMux_io_out_bits_wstrb_20),
    .io_out_bits_wstrb_21(wdataMux_io_out_bits_wstrb_21),
    .io_out_bits_wstrb_22(wdataMux_io_out_bits_wstrb_22),
    .io_out_bits_wstrb_23(wdataMux_io_out_bits_wstrb_23),
    .io_out_bits_wstrb_24(wdataMux_io_out_bits_wstrb_24),
    .io_out_bits_wstrb_25(wdataMux_io_out_bits_wstrb_25),
    .io_out_bits_wstrb_26(wdataMux_io_out_bits_wstrb_26),
    .io_out_bits_wstrb_27(wdataMux_io_out_bits_wstrb_27),
    .io_out_bits_wstrb_28(wdataMux_io_out_bits_wstrb_28),
    .io_out_bits_wstrb_29(wdataMux_io_out_bits_wstrb_29),
    .io_out_bits_wstrb_30(wdataMux_io_out_bits_wstrb_30),
    .io_out_bits_wstrb_31(wdataMux_io_out_bits_wstrb_31),
    .io_out_bits_wstrb_32(wdataMux_io_out_bits_wstrb_32),
    .io_out_bits_wstrb_33(wdataMux_io_out_bits_wstrb_33),
    .io_out_bits_wstrb_34(wdataMux_io_out_bits_wstrb_34),
    .io_out_bits_wstrb_35(wdataMux_io_out_bits_wstrb_35),
    .io_out_bits_wstrb_36(wdataMux_io_out_bits_wstrb_36),
    .io_out_bits_wstrb_37(wdataMux_io_out_bits_wstrb_37),
    .io_out_bits_wstrb_38(wdataMux_io_out_bits_wstrb_38),
    .io_out_bits_wstrb_39(wdataMux_io_out_bits_wstrb_39),
    .io_out_bits_wstrb_40(wdataMux_io_out_bits_wstrb_40),
    .io_out_bits_wstrb_41(wdataMux_io_out_bits_wstrb_41),
    .io_out_bits_wstrb_42(wdataMux_io_out_bits_wstrb_42),
    .io_out_bits_wstrb_43(wdataMux_io_out_bits_wstrb_43),
    .io_out_bits_wstrb_44(wdataMux_io_out_bits_wstrb_44),
    .io_out_bits_wstrb_45(wdataMux_io_out_bits_wstrb_45),
    .io_out_bits_wstrb_46(wdataMux_io_out_bits_wstrb_46),
    .io_out_bits_wstrb_47(wdataMux_io_out_bits_wstrb_47),
    .io_out_bits_wstrb_48(wdataMux_io_out_bits_wstrb_48),
    .io_out_bits_wstrb_49(wdataMux_io_out_bits_wstrb_49),
    .io_out_bits_wstrb_50(wdataMux_io_out_bits_wstrb_50),
    .io_out_bits_wstrb_51(wdataMux_io_out_bits_wstrb_51),
    .io_out_bits_wstrb_52(wdataMux_io_out_bits_wstrb_52),
    .io_out_bits_wstrb_53(wdataMux_io_out_bits_wstrb_53),
    .io_out_bits_wstrb_54(wdataMux_io_out_bits_wstrb_54),
    .io_out_bits_wstrb_55(wdataMux_io_out_bits_wstrb_55),
    .io_out_bits_wstrb_56(wdataMux_io_out_bits_wstrb_56),
    .io_out_bits_wstrb_57(wdataMux_io_out_bits_wstrb_57),
    .io_out_bits_wstrb_58(wdataMux_io_out_bits_wstrb_58),
    .io_out_bits_wstrb_59(wdataMux_io_out_bits_wstrb_59),
    .io_out_bits_wstrb_60(wdataMux_io_out_bits_wstrb_60),
    .io_out_bits_wstrb_61(wdataMux_io_out_bits_wstrb_61),
    .io_out_bits_wstrb_62(wdataMux_io_out_bits_wstrb_62),
    .io_out_bits_wstrb_63(wdataMux_io_out_bits_wstrb_63)
  );
  ElementCounter elementCtr ( // @[StreamArbiter.scala 36:26:@47804.4]
    .clock(elementCtr_clock),
    .reset(elementCtr_reset),
    .io_reset(elementCtr_io_reset),
    .io_enable(elementCtr_io_enable),
    .io_out(elementCtr_io_out)
  );
  assign _T_346 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@47773.4 package.scala 96:25:@47774.4]
  assign cmdIdx = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[StreamArbiter.scala 21:16:@47775.4]
  assign cmdInDecoder = 2'h1 << cmdIdx; // @[OneHot.scala 45:35:@47777.4]
  assign _T_355 = io_app_0_cmd_bits_tag[8]; // @[FringeBundles.scala 114:28:@47793.4]
  assign _T_356 = io_app_0_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@47795.4]
  assign _T_358 = {_T_356,_T_355}; // @[FringeBundles.scala 115:37:@47798.4]
  assign _T_360 = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:49:@47807.4]
  assign _T_365 = cmdMux_io_out_bits_tag; // @[:@47811.4 :@47812.4]
  assign _T_366 = _T_365[7:0]; // @[FringeBundles.scala 114:28:@47813.4]
  assign cmdOutDecoder = 256'h1 << _T_366; // @[OneHot.scala 45:35:@47819.4]
  assign _T_379 = io_app_0_wdata_valid & cmdMux_io_out_valid; // @[StreamArbiter.scala 42:78:@47822.4]
  assign _T_380 = elementCtr_io_out < cmdMux_io_out_bits_size; // @[StreamArbiter.scala 42:121:@47823.4]
  assign _T_395 = io_dram_wresp_bits_tag[7:0]; // @[FringeBundles.scala 140:28:@48010.4]
  assign wrespDecoder = 256'h1 << _T_395; // @[OneHot.scala 45:35:@48017.4]
  assign _T_400 = cmdInDecoder[0]; // @[StreamArbiter.scala 61:55:@48022.4]
  assign _T_403 = cmdOutDecoder[0]; // @[StreamArbiter.scala 62:85:@48026.4]
  assign _T_404 = _T_360 & _T_403; // @[StreamArbiter.scala 62:70:@48027.4]
  assign _T_409 = wrespDecoder[0]; // @[StreamArbiter.scala 67:58:@48051.4]
  assign io_app_0_cmd_ready = cmdMux_io_in_ready & _T_400; // @[StreamArbiter.scala 61:19:@48024.4]
  assign io_app_0_wdata_ready = _T_404 & _T_380; // @[StreamArbiter.scala 62:21:@48030.4]
  assign io_app_0_wresp_valid = io_dram_wresp_valid & _T_409; // @[StreamArbiter.scala 67:21:@48053.4]
  assign io_dram_cmd_valid = cmdMux_io_out_valid; // @[StreamArbiter.scala 46:15:@47913.4]
  assign io_dram_cmd_bits_addr = cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 46:15:@47912.4]
  assign io_dram_cmd_bits_size = cmdMux_io_out_bits_size; // @[StreamArbiter.scala 46:15:@47911.4]
  assign io_dram_cmd_bits_isWr = cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 46:15:@47909.4]
  assign io_dram_cmd_bits_tag = cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 46:15:@47908.4]
  assign io_dram_wdata_valid = wdataMux_io_out_valid; // @[StreamArbiter.scala 47:17:@47996.4]
  assign io_dram_wdata_bits_wdata_0 = wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 47:17:@47980.4]
  assign io_dram_wdata_bits_wdata_1 = wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 47:17:@47981.4]
  assign io_dram_wdata_bits_wdata_2 = wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 47:17:@47982.4]
  assign io_dram_wdata_bits_wdata_3 = wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 47:17:@47983.4]
  assign io_dram_wdata_bits_wdata_4 = wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 47:17:@47984.4]
  assign io_dram_wdata_bits_wdata_5 = wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 47:17:@47985.4]
  assign io_dram_wdata_bits_wdata_6 = wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 47:17:@47986.4]
  assign io_dram_wdata_bits_wdata_7 = wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 47:17:@47987.4]
  assign io_dram_wdata_bits_wdata_8 = wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 47:17:@47988.4]
  assign io_dram_wdata_bits_wdata_9 = wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 47:17:@47989.4]
  assign io_dram_wdata_bits_wdata_10 = wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 47:17:@47990.4]
  assign io_dram_wdata_bits_wdata_11 = wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 47:17:@47991.4]
  assign io_dram_wdata_bits_wdata_12 = wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 47:17:@47992.4]
  assign io_dram_wdata_bits_wdata_13 = wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 47:17:@47993.4]
  assign io_dram_wdata_bits_wdata_14 = wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 47:17:@47994.4]
  assign io_dram_wdata_bits_wdata_15 = wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 47:17:@47995.4]
  assign io_dram_wdata_bits_wstrb_0 = wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 47:17:@47916.4]
  assign io_dram_wdata_bits_wstrb_1 = wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 47:17:@47917.4]
  assign io_dram_wdata_bits_wstrb_2 = wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 47:17:@47918.4]
  assign io_dram_wdata_bits_wstrb_3 = wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 47:17:@47919.4]
  assign io_dram_wdata_bits_wstrb_4 = wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 47:17:@47920.4]
  assign io_dram_wdata_bits_wstrb_5 = wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 47:17:@47921.4]
  assign io_dram_wdata_bits_wstrb_6 = wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 47:17:@47922.4]
  assign io_dram_wdata_bits_wstrb_7 = wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 47:17:@47923.4]
  assign io_dram_wdata_bits_wstrb_8 = wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 47:17:@47924.4]
  assign io_dram_wdata_bits_wstrb_9 = wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 47:17:@47925.4]
  assign io_dram_wdata_bits_wstrb_10 = wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 47:17:@47926.4]
  assign io_dram_wdata_bits_wstrb_11 = wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 47:17:@47927.4]
  assign io_dram_wdata_bits_wstrb_12 = wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 47:17:@47928.4]
  assign io_dram_wdata_bits_wstrb_13 = wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 47:17:@47929.4]
  assign io_dram_wdata_bits_wstrb_14 = wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 47:17:@47930.4]
  assign io_dram_wdata_bits_wstrb_15 = wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 47:17:@47931.4]
  assign io_dram_wdata_bits_wstrb_16 = wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 47:17:@47932.4]
  assign io_dram_wdata_bits_wstrb_17 = wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 47:17:@47933.4]
  assign io_dram_wdata_bits_wstrb_18 = wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 47:17:@47934.4]
  assign io_dram_wdata_bits_wstrb_19 = wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 47:17:@47935.4]
  assign io_dram_wdata_bits_wstrb_20 = wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 47:17:@47936.4]
  assign io_dram_wdata_bits_wstrb_21 = wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 47:17:@47937.4]
  assign io_dram_wdata_bits_wstrb_22 = wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 47:17:@47938.4]
  assign io_dram_wdata_bits_wstrb_23 = wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 47:17:@47939.4]
  assign io_dram_wdata_bits_wstrb_24 = wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 47:17:@47940.4]
  assign io_dram_wdata_bits_wstrb_25 = wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 47:17:@47941.4]
  assign io_dram_wdata_bits_wstrb_26 = wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 47:17:@47942.4]
  assign io_dram_wdata_bits_wstrb_27 = wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 47:17:@47943.4]
  assign io_dram_wdata_bits_wstrb_28 = wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 47:17:@47944.4]
  assign io_dram_wdata_bits_wstrb_29 = wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 47:17:@47945.4]
  assign io_dram_wdata_bits_wstrb_30 = wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 47:17:@47946.4]
  assign io_dram_wdata_bits_wstrb_31 = wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 47:17:@47947.4]
  assign io_dram_wdata_bits_wstrb_32 = wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 47:17:@47948.4]
  assign io_dram_wdata_bits_wstrb_33 = wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 47:17:@47949.4]
  assign io_dram_wdata_bits_wstrb_34 = wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 47:17:@47950.4]
  assign io_dram_wdata_bits_wstrb_35 = wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 47:17:@47951.4]
  assign io_dram_wdata_bits_wstrb_36 = wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 47:17:@47952.4]
  assign io_dram_wdata_bits_wstrb_37 = wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 47:17:@47953.4]
  assign io_dram_wdata_bits_wstrb_38 = wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 47:17:@47954.4]
  assign io_dram_wdata_bits_wstrb_39 = wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 47:17:@47955.4]
  assign io_dram_wdata_bits_wstrb_40 = wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 47:17:@47956.4]
  assign io_dram_wdata_bits_wstrb_41 = wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 47:17:@47957.4]
  assign io_dram_wdata_bits_wstrb_42 = wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 47:17:@47958.4]
  assign io_dram_wdata_bits_wstrb_43 = wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 47:17:@47959.4]
  assign io_dram_wdata_bits_wstrb_44 = wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 47:17:@47960.4]
  assign io_dram_wdata_bits_wstrb_45 = wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 47:17:@47961.4]
  assign io_dram_wdata_bits_wstrb_46 = wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 47:17:@47962.4]
  assign io_dram_wdata_bits_wstrb_47 = wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 47:17:@47963.4]
  assign io_dram_wdata_bits_wstrb_48 = wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 47:17:@47964.4]
  assign io_dram_wdata_bits_wstrb_49 = wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 47:17:@47965.4]
  assign io_dram_wdata_bits_wstrb_50 = wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 47:17:@47966.4]
  assign io_dram_wdata_bits_wstrb_51 = wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 47:17:@47967.4]
  assign io_dram_wdata_bits_wstrb_52 = wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 47:17:@47968.4]
  assign io_dram_wdata_bits_wstrb_53 = wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 47:17:@47969.4]
  assign io_dram_wdata_bits_wstrb_54 = wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 47:17:@47970.4]
  assign io_dram_wdata_bits_wstrb_55 = wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 47:17:@47971.4]
  assign io_dram_wdata_bits_wstrb_56 = wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 47:17:@47972.4]
  assign io_dram_wdata_bits_wstrb_57 = wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 47:17:@47973.4]
  assign io_dram_wdata_bits_wstrb_58 = wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 47:17:@47974.4]
  assign io_dram_wdata_bits_wstrb_59 = wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 47:17:@47975.4]
  assign io_dram_wdata_bits_wstrb_60 = wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 47:17:@47976.4]
  assign io_dram_wdata_bits_wstrb_61 = wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 47:17:@47977.4]
  assign io_dram_wdata_bits_wstrb_62 = wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 47:17:@47978.4]
  assign io_dram_wdata_bits_wstrb_63 = wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 47:17:@47979.4]
  assign io_dram_rresp_ready = io_app_0_rresp_ready; // @[StreamArbiter.scala 72:23:@48057.4]
  assign io_dram_wresp_ready = io_app_0_wresp_ready; // @[StreamArbiter.scala 73:23:@48060.4]
  assign RetimeWrapper_clock = clock; // @[:@47762.4]
  assign RetimeWrapper_reset = reset; // @[:@47763.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@47765.4]
  assign RetimeWrapper_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@47764.4]
  assign RetimeWrapper_1_clock = clock; // @[:@47769.4]
  assign RetimeWrapper_1_reset = reset; // @[:@47770.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@47772.4]
  assign RetimeWrapper_1_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@47771.4]
  assign cmdMux_io_in_valid = io_app_0_cmd_valid; // @[StreamArbiter.scala 26:22:@47781.4]
  assign cmdMux_io_in_bits_0_addr = io_app_0_cmd_bits_addr; // @[StreamArbiter.scala 29:9:@47787.4]
  assign cmdMux_io_in_bits_0_size = io_app_0_cmd_bits_size; // @[StreamArbiter.scala 29:9:@47786.4]
  assign cmdMux_io_in_bits_0_isWr = io_app_0_cmd_bits_isWr; // @[StreamArbiter.scala 29:9:@47784.4]
  assign cmdMux_io_in_bits_0_tag = {_T_358,8'h0}; // @[StreamArbiter.scala 29:9:@47783.4 FringeBundles.scala 115:32:@47800.4]
  assign cmdMux_io_out_ready = io_dram_cmd_valid & io_dram_cmd_ready; // @[StreamArbiter.scala 46:15:@47914.4 StreamArbiter.scala 57:23:@48020.4]
  assign wdataMux_io_in_valid = _T_379 & _T_380; // @[StreamArbiter.scala 42:24:@47825.4]
  assign wdataMux_io_in_bits_0_wdata_0 = io_app_0_wdata_bits_wdata_0; // @[StreamArbiter.scala 44:23:@47892.4]
  assign wdataMux_io_in_bits_0_wdata_1 = io_app_0_wdata_bits_wdata_1; // @[StreamArbiter.scala 44:23:@47893.4]
  assign wdataMux_io_in_bits_0_wdata_2 = io_app_0_wdata_bits_wdata_2; // @[StreamArbiter.scala 44:23:@47894.4]
  assign wdataMux_io_in_bits_0_wdata_3 = io_app_0_wdata_bits_wdata_3; // @[StreamArbiter.scala 44:23:@47895.4]
  assign wdataMux_io_in_bits_0_wdata_4 = io_app_0_wdata_bits_wdata_4; // @[StreamArbiter.scala 44:23:@47896.4]
  assign wdataMux_io_in_bits_0_wdata_5 = io_app_0_wdata_bits_wdata_5; // @[StreamArbiter.scala 44:23:@47897.4]
  assign wdataMux_io_in_bits_0_wdata_6 = io_app_0_wdata_bits_wdata_6; // @[StreamArbiter.scala 44:23:@47898.4]
  assign wdataMux_io_in_bits_0_wdata_7 = io_app_0_wdata_bits_wdata_7; // @[StreamArbiter.scala 44:23:@47899.4]
  assign wdataMux_io_in_bits_0_wdata_8 = io_app_0_wdata_bits_wdata_8; // @[StreamArbiter.scala 44:23:@47900.4]
  assign wdataMux_io_in_bits_0_wdata_9 = io_app_0_wdata_bits_wdata_9; // @[StreamArbiter.scala 44:23:@47901.4]
  assign wdataMux_io_in_bits_0_wdata_10 = io_app_0_wdata_bits_wdata_10; // @[StreamArbiter.scala 44:23:@47902.4]
  assign wdataMux_io_in_bits_0_wdata_11 = io_app_0_wdata_bits_wdata_11; // @[StreamArbiter.scala 44:23:@47903.4]
  assign wdataMux_io_in_bits_0_wdata_12 = io_app_0_wdata_bits_wdata_12; // @[StreamArbiter.scala 44:23:@47904.4]
  assign wdataMux_io_in_bits_0_wdata_13 = io_app_0_wdata_bits_wdata_13; // @[StreamArbiter.scala 44:23:@47905.4]
  assign wdataMux_io_in_bits_0_wdata_14 = io_app_0_wdata_bits_wdata_14; // @[StreamArbiter.scala 44:23:@47906.4]
  assign wdataMux_io_in_bits_0_wdata_15 = io_app_0_wdata_bits_wdata_15; // @[StreamArbiter.scala 44:23:@47907.4]
  assign wdataMux_io_in_bits_0_wstrb_0 = io_app_0_wdata_bits_wstrb_0; // @[StreamArbiter.scala 44:23:@47828.4]
  assign wdataMux_io_in_bits_0_wstrb_1 = io_app_0_wdata_bits_wstrb_1; // @[StreamArbiter.scala 44:23:@47829.4]
  assign wdataMux_io_in_bits_0_wstrb_2 = io_app_0_wdata_bits_wstrb_2; // @[StreamArbiter.scala 44:23:@47830.4]
  assign wdataMux_io_in_bits_0_wstrb_3 = io_app_0_wdata_bits_wstrb_3; // @[StreamArbiter.scala 44:23:@47831.4]
  assign wdataMux_io_in_bits_0_wstrb_4 = io_app_0_wdata_bits_wstrb_4; // @[StreamArbiter.scala 44:23:@47832.4]
  assign wdataMux_io_in_bits_0_wstrb_5 = io_app_0_wdata_bits_wstrb_5; // @[StreamArbiter.scala 44:23:@47833.4]
  assign wdataMux_io_in_bits_0_wstrb_6 = io_app_0_wdata_bits_wstrb_6; // @[StreamArbiter.scala 44:23:@47834.4]
  assign wdataMux_io_in_bits_0_wstrb_7 = io_app_0_wdata_bits_wstrb_7; // @[StreamArbiter.scala 44:23:@47835.4]
  assign wdataMux_io_in_bits_0_wstrb_8 = io_app_0_wdata_bits_wstrb_8; // @[StreamArbiter.scala 44:23:@47836.4]
  assign wdataMux_io_in_bits_0_wstrb_9 = io_app_0_wdata_bits_wstrb_9; // @[StreamArbiter.scala 44:23:@47837.4]
  assign wdataMux_io_in_bits_0_wstrb_10 = io_app_0_wdata_bits_wstrb_10; // @[StreamArbiter.scala 44:23:@47838.4]
  assign wdataMux_io_in_bits_0_wstrb_11 = io_app_0_wdata_bits_wstrb_11; // @[StreamArbiter.scala 44:23:@47839.4]
  assign wdataMux_io_in_bits_0_wstrb_12 = io_app_0_wdata_bits_wstrb_12; // @[StreamArbiter.scala 44:23:@47840.4]
  assign wdataMux_io_in_bits_0_wstrb_13 = io_app_0_wdata_bits_wstrb_13; // @[StreamArbiter.scala 44:23:@47841.4]
  assign wdataMux_io_in_bits_0_wstrb_14 = io_app_0_wdata_bits_wstrb_14; // @[StreamArbiter.scala 44:23:@47842.4]
  assign wdataMux_io_in_bits_0_wstrb_15 = io_app_0_wdata_bits_wstrb_15; // @[StreamArbiter.scala 44:23:@47843.4]
  assign wdataMux_io_in_bits_0_wstrb_16 = io_app_0_wdata_bits_wstrb_16; // @[StreamArbiter.scala 44:23:@47844.4]
  assign wdataMux_io_in_bits_0_wstrb_17 = io_app_0_wdata_bits_wstrb_17; // @[StreamArbiter.scala 44:23:@47845.4]
  assign wdataMux_io_in_bits_0_wstrb_18 = io_app_0_wdata_bits_wstrb_18; // @[StreamArbiter.scala 44:23:@47846.4]
  assign wdataMux_io_in_bits_0_wstrb_19 = io_app_0_wdata_bits_wstrb_19; // @[StreamArbiter.scala 44:23:@47847.4]
  assign wdataMux_io_in_bits_0_wstrb_20 = io_app_0_wdata_bits_wstrb_20; // @[StreamArbiter.scala 44:23:@47848.4]
  assign wdataMux_io_in_bits_0_wstrb_21 = io_app_0_wdata_bits_wstrb_21; // @[StreamArbiter.scala 44:23:@47849.4]
  assign wdataMux_io_in_bits_0_wstrb_22 = io_app_0_wdata_bits_wstrb_22; // @[StreamArbiter.scala 44:23:@47850.4]
  assign wdataMux_io_in_bits_0_wstrb_23 = io_app_0_wdata_bits_wstrb_23; // @[StreamArbiter.scala 44:23:@47851.4]
  assign wdataMux_io_in_bits_0_wstrb_24 = io_app_0_wdata_bits_wstrb_24; // @[StreamArbiter.scala 44:23:@47852.4]
  assign wdataMux_io_in_bits_0_wstrb_25 = io_app_0_wdata_bits_wstrb_25; // @[StreamArbiter.scala 44:23:@47853.4]
  assign wdataMux_io_in_bits_0_wstrb_26 = io_app_0_wdata_bits_wstrb_26; // @[StreamArbiter.scala 44:23:@47854.4]
  assign wdataMux_io_in_bits_0_wstrb_27 = io_app_0_wdata_bits_wstrb_27; // @[StreamArbiter.scala 44:23:@47855.4]
  assign wdataMux_io_in_bits_0_wstrb_28 = io_app_0_wdata_bits_wstrb_28; // @[StreamArbiter.scala 44:23:@47856.4]
  assign wdataMux_io_in_bits_0_wstrb_29 = io_app_0_wdata_bits_wstrb_29; // @[StreamArbiter.scala 44:23:@47857.4]
  assign wdataMux_io_in_bits_0_wstrb_30 = io_app_0_wdata_bits_wstrb_30; // @[StreamArbiter.scala 44:23:@47858.4]
  assign wdataMux_io_in_bits_0_wstrb_31 = io_app_0_wdata_bits_wstrb_31; // @[StreamArbiter.scala 44:23:@47859.4]
  assign wdataMux_io_in_bits_0_wstrb_32 = io_app_0_wdata_bits_wstrb_32; // @[StreamArbiter.scala 44:23:@47860.4]
  assign wdataMux_io_in_bits_0_wstrb_33 = io_app_0_wdata_bits_wstrb_33; // @[StreamArbiter.scala 44:23:@47861.4]
  assign wdataMux_io_in_bits_0_wstrb_34 = io_app_0_wdata_bits_wstrb_34; // @[StreamArbiter.scala 44:23:@47862.4]
  assign wdataMux_io_in_bits_0_wstrb_35 = io_app_0_wdata_bits_wstrb_35; // @[StreamArbiter.scala 44:23:@47863.4]
  assign wdataMux_io_in_bits_0_wstrb_36 = io_app_0_wdata_bits_wstrb_36; // @[StreamArbiter.scala 44:23:@47864.4]
  assign wdataMux_io_in_bits_0_wstrb_37 = io_app_0_wdata_bits_wstrb_37; // @[StreamArbiter.scala 44:23:@47865.4]
  assign wdataMux_io_in_bits_0_wstrb_38 = io_app_0_wdata_bits_wstrb_38; // @[StreamArbiter.scala 44:23:@47866.4]
  assign wdataMux_io_in_bits_0_wstrb_39 = io_app_0_wdata_bits_wstrb_39; // @[StreamArbiter.scala 44:23:@47867.4]
  assign wdataMux_io_in_bits_0_wstrb_40 = io_app_0_wdata_bits_wstrb_40; // @[StreamArbiter.scala 44:23:@47868.4]
  assign wdataMux_io_in_bits_0_wstrb_41 = io_app_0_wdata_bits_wstrb_41; // @[StreamArbiter.scala 44:23:@47869.4]
  assign wdataMux_io_in_bits_0_wstrb_42 = io_app_0_wdata_bits_wstrb_42; // @[StreamArbiter.scala 44:23:@47870.4]
  assign wdataMux_io_in_bits_0_wstrb_43 = io_app_0_wdata_bits_wstrb_43; // @[StreamArbiter.scala 44:23:@47871.4]
  assign wdataMux_io_in_bits_0_wstrb_44 = io_app_0_wdata_bits_wstrb_44; // @[StreamArbiter.scala 44:23:@47872.4]
  assign wdataMux_io_in_bits_0_wstrb_45 = io_app_0_wdata_bits_wstrb_45; // @[StreamArbiter.scala 44:23:@47873.4]
  assign wdataMux_io_in_bits_0_wstrb_46 = io_app_0_wdata_bits_wstrb_46; // @[StreamArbiter.scala 44:23:@47874.4]
  assign wdataMux_io_in_bits_0_wstrb_47 = io_app_0_wdata_bits_wstrb_47; // @[StreamArbiter.scala 44:23:@47875.4]
  assign wdataMux_io_in_bits_0_wstrb_48 = io_app_0_wdata_bits_wstrb_48; // @[StreamArbiter.scala 44:23:@47876.4]
  assign wdataMux_io_in_bits_0_wstrb_49 = io_app_0_wdata_bits_wstrb_49; // @[StreamArbiter.scala 44:23:@47877.4]
  assign wdataMux_io_in_bits_0_wstrb_50 = io_app_0_wdata_bits_wstrb_50; // @[StreamArbiter.scala 44:23:@47878.4]
  assign wdataMux_io_in_bits_0_wstrb_51 = io_app_0_wdata_bits_wstrb_51; // @[StreamArbiter.scala 44:23:@47879.4]
  assign wdataMux_io_in_bits_0_wstrb_52 = io_app_0_wdata_bits_wstrb_52; // @[StreamArbiter.scala 44:23:@47880.4]
  assign wdataMux_io_in_bits_0_wstrb_53 = io_app_0_wdata_bits_wstrb_53; // @[StreamArbiter.scala 44:23:@47881.4]
  assign wdataMux_io_in_bits_0_wstrb_54 = io_app_0_wdata_bits_wstrb_54; // @[StreamArbiter.scala 44:23:@47882.4]
  assign wdataMux_io_in_bits_0_wstrb_55 = io_app_0_wdata_bits_wstrb_55; // @[StreamArbiter.scala 44:23:@47883.4]
  assign wdataMux_io_in_bits_0_wstrb_56 = io_app_0_wdata_bits_wstrb_56; // @[StreamArbiter.scala 44:23:@47884.4]
  assign wdataMux_io_in_bits_0_wstrb_57 = io_app_0_wdata_bits_wstrb_57; // @[StreamArbiter.scala 44:23:@47885.4]
  assign wdataMux_io_in_bits_0_wstrb_58 = io_app_0_wdata_bits_wstrb_58; // @[StreamArbiter.scala 44:23:@47886.4]
  assign wdataMux_io_in_bits_0_wstrb_59 = io_app_0_wdata_bits_wstrb_59; // @[StreamArbiter.scala 44:23:@47887.4]
  assign wdataMux_io_in_bits_0_wstrb_60 = io_app_0_wdata_bits_wstrb_60; // @[StreamArbiter.scala 44:23:@47888.4]
  assign wdataMux_io_in_bits_0_wstrb_61 = io_app_0_wdata_bits_wstrb_61; // @[StreamArbiter.scala 44:23:@47889.4]
  assign wdataMux_io_in_bits_0_wstrb_62 = io_app_0_wdata_bits_wstrb_62; // @[StreamArbiter.scala 44:23:@47890.4]
  assign wdataMux_io_in_bits_0_wstrb_63 = io_app_0_wdata_bits_wstrb_63; // @[StreamArbiter.scala 44:23:@47891.4]
  assign wdataMux_io_out_ready = io_dram_wdata_valid & io_dram_wdata_ready; // @[StreamArbiter.scala 47:17:@47997.4 StreamArbiter.scala 58:25:@48021.4]
  assign elementCtr_clock = clock; // @[:@47805.4]
  assign elementCtr_reset = reset; // @[:@47806.4]
  assign elementCtr_io_reset = cmdMux_io_out_ready; // @[StreamArbiter.scala 38:23:@47809.4]
  assign elementCtr_io_enable = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:24:@47808.4]
endmodule
module Counter_72( // @[:@48062.2]
  input         clock, // @[:@48063.4]
  input         reset, // @[:@48064.4]
  input         io_reset, // @[:@48065.4]
  input         io_enable, // @[:@48065.4]
  input  [31:0] io_stride, // @[:@48065.4]
  output [31:0] io_out, // @[:@48065.4]
  output [31:0] io_next // @[:@48065.4]
);
  reg [31:0] count; // @[Counter.scala 15:22:@48067.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_17; // @[Counter.scala 17:24:@48068.4]
  wire [31:0] newCount; // @[Counter.scala 17:24:@48069.4]
  wire [31:0] _GEN_0; // @[Counter.scala 21:26:@48074.6]
  wire [31:0] _GEN_1; // @[Counter.scala 19:18:@48070.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@48068.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@48069.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@48074.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 19:18:@48070.4]
  assign io_out = count; // @[Counter.scala 25:10:@48077.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@48078.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module AXICmdSplit( // @[:@48080.2]
  input         clock, // @[:@48081.4]
  input         reset, // @[:@48082.4]
  output        io_in_cmd_ready, // @[:@48083.4]
  input         io_in_cmd_valid, // @[:@48083.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@48083.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@48083.4]
  input         io_in_cmd_bits_isWr, // @[:@48083.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@48083.4]
  output        io_in_wdata_ready, // @[:@48083.4]
  input         io_in_wdata_valid, // @[:@48083.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@48083.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@48083.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@48083.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@48083.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@48083.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@48083.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@48083.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@48083.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@48083.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@48083.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@48083.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@48083.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@48083.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@48083.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@48083.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@48083.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@48083.4]
  input         io_in_rresp_ready, // @[:@48083.4]
  input         io_in_wresp_ready, // @[:@48083.4]
  output        io_in_wresp_valid, // @[:@48083.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@48083.4]
  input         io_out_cmd_ready, // @[:@48083.4]
  output        io_out_cmd_valid, // @[:@48083.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@48083.4]
  output [31:0] io_out_cmd_bits_size, // @[:@48083.4]
  output        io_out_cmd_bits_isWr, // @[:@48083.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@48083.4]
  input         io_out_wdata_ready, // @[:@48083.4]
  output        io_out_wdata_valid, // @[:@48083.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@48083.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@48083.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@48083.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@48083.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@48083.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@48083.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@48083.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@48083.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@48083.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@48083.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@48083.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@48083.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@48083.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@48083.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@48083.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@48083.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@48083.4]
  output        io_out_rresp_ready, // @[:@48083.4]
  output        io_out_wresp_ready, // @[:@48083.4]
  input         io_out_wresp_valid, // @[:@48083.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@48083.4]
);
  wire  cmdSizeCounter_clock; // @[AXIProtocol.scala 18:30:@48197.4]
  wire  cmdSizeCounter_reset; // @[AXIProtocol.scala 18:30:@48197.4]
  wire  cmdSizeCounter_io_reset; // @[AXIProtocol.scala 18:30:@48197.4]
  wire  cmdSizeCounter_io_enable; // @[AXIProtocol.scala 18:30:@48197.4]
  wire [31:0] cmdSizeCounter_io_stride; // @[AXIProtocol.scala 18:30:@48197.4]
  wire [31:0] cmdSizeCounter_io_out; // @[AXIProtocol.scala 18:30:@48197.4]
  wire [31:0] cmdSizeCounter_io_next; // @[AXIProtocol.scala 18:30:@48197.4]
  wire [32:0] _T_199; // @[AXIProtocol.scala 20:46:@48200.4]
  wire [32:0] _T_200; // @[AXIProtocol.scala 20:46:@48201.4]
  wire [31:0] cmdSizeRemaining; // @[AXIProtocol.scala 20:46:@48202.4]
  wire  lastCmd; // @[AXIProtocol.scala 23:35:@48203.4]
  wire [37:0] _GEN_0; // @[AXIProtocol.scala 27:47:@48206.4]
  wire [37:0] addrOffsetBytes; // @[AXIProtocol.scala 27:47:@48206.4]
  wire [63:0] _GEN_1; // @[AXIProtocol.scala 28:49:@48207.4]
  wire [64:0] _T_201; // @[AXIProtocol.scala 28:49:@48207.4]
  wire [63:0] cmdAddr_bits; // @[AXIProtocol.scala 28:49:@48208.4]
  wire [57:0] _T_204; // @[FringeBundles.scala 158:22:@48211.4]
  wire [7:0] cmdTag_streamID; // @[FringeBundles.scala 114:28:@48218.4]
  wire [22:0] cmdTag_uid; // @[FringeBundles.scala 114:28:@48222.4]
  wire [23:0] _T_214; // @[FringeBundles.scala 115:37:@48225.4]
  wire  cmdIssue; // @[AXIProtocol.scala 36:35:@48228.4]
  wire  _T_223; // @[FringeBundles.scala 140:28:@48239.4]
  Counter_72 cmdSizeCounter ( // @[AXIProtocol.scala 18:30:@48197.4]
    .clock(cmdSizeCounter_clock),
    .reset(cmdSizeCounter_reset),
    .io_reset(cmdSizeCounter_io_reset),
    .io_enable(cmdSizeCounter_io_enable),
    .io_stride(cmdSizeCounter_io_stride),
    .io_out(cmdSizeCounter_io_out),
    .io_next(cmdSizeCounter_io_next)
  );
  assign _T_199 = io_in_cmd_bits_size - cmdSizeCounter_io_out; // @[AXIProtocol.scala 20:46:@48200.4]
  assign _T_200 = $unsigned(_T_199); // @[AXIProtocol.scala 20:46:@48201.4]
  assign cmdSizeRemaining = _T_200[31:0]; // @[AXIProtocol.scala 20:46:@48202.4]
  assign lastCmd = cmdSizeRemaining <= 32'h100; // @[AXIProtocol.scala 23:35:@48203.4]
  assign _GEN_0 = {{6'd0}, cmdSizeCounter_io_out}; // @[AXIProtocol.scala 27:47:@48206.4]
  assign addrOffsetBytes = _GEN_0 << 6; // @[AXIProtocol.scala 27:47:@48206.4]
  assign _GEN_1 = {{26'd0}, addrOffsetBytes}; // @[AXIProtocol.scala 28:49:@48207.4]
  assign _T_201 = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@48207.4]
  assign cmdAddr_bits = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@48208.4]
  assign _T_204 = cmdAddr_bits[63:6]; // @[FringeBundles.scala 158:22:@48211.4]
  assign cmdTag_streamID = io_in_cmd_bits_tag[7:0]; // @[FringeBundles.scala 114:28:@48218.4]
  assign cmdTag_uid = io_in_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@48222.4]
  assign _T_214 = {cmdTag_uid,lastCmd}; // @[FringeBundles.scala 115:37:@48225.4]
  assign cmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 36:35:@48228.4]
  assign _T_223 = io_out_wresp_bits_tag[8]; // @[FringeBundles.scala 140:28:@48239.4]
  assign io_in_cmd_ready = lastCmd & cmdIssue; // @[AXIProtocol.scala 15:10:@48196.4 AXIProtocol.scala 38:19:@48230.4]
  assign io_in_wdata_ready = io_out_wdata_ready; // @[AXIProtocol.scala 15:10:@48189.4]
  assign io_in_wresp_valid = io_out_wresp_valid & _T_223; // @[AXIProtocol.scala 15:10:@48086.4 AXIProtocol.scala 46:21:@48244.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 15:10:@48085.4]
  assign io_out_cmd_valid = io_in_cmd_valid; // @[AXIProtocol.scala 15:10:@48195.4]
  assign io_out_cmd_bits_addr = {_T_204,6'h0}; // @[AXIProtocol.scala 15:10:@48194.4 AXIProtocol.scala 29:24:@48213.4]
  assign io_out_cmd_bits_size = lastCmd ? cmdSizeRemaining : 32'h100; // @[AXIProtocol.scala 15:10:@48193.4 AXIProtocol.scala 25:24:@48205.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 15:10:@48191.4]
  assign io_out_cmd_bits_tag = {_T_214,cmdTag_streamID}; // @[AXIProtocol.scala 15:10:@48190.4 FringeBundles.scala 115:32:@48227.4]
  assign io_out_wdata_valid = io_in_wdata_valid; // @[AXIProtocol.scala 15:10:@48188.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 15:10:@48172.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 15:10:@48173.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 15:10:@48174.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 15:10:@48175.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 15:10:@48176.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 15:10:@48177.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 15:10:@48178.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 15:10:@48179.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 15:10:@48180.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 15:10:@48181.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 15:10:@48182.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 15:10:@48183.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 15:10:@48184.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 15:10:@48185.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 15:10:@48186.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 15:10:@48187.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 15:10:@48108.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 15:10:@48109.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 15:10:@48110.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 15:10:@48111.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 15:10:@48112.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 15:10:@48113.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 15:10:@48114.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 15:10:@48115.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 15:10:@48116.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 15:10:@48117.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 15:10:@48118.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 15:10:@48119.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 15:10:@48120.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 15:10:@48121.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 15:10:@48122.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 15:10:@48123.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 15:10:@48124.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 15:10:@48125.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 15:10:@48126.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 15:10:@48127.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 15:10:@48128.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 15:10:@48129.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 15:10:@48130.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 15:10:@48131.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 15:10:@48132.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 15:10:@48133.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 15:10:@48134.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 15:10:@48135.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 15:10:@48136.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 15:10:@48137.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 15:10:@48138.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 15:10:@48139.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 15:10:@48140.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 15:10:@48141.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 15:10:@48142.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 15:10:@48143.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 15:10:@48144.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 15:10:@48145.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 15:10:@48146.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 15:10:@48147.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 15:10:@48148.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 15:10:@48149.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 15:10:@48150.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 15:10:@48151.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 15:10:@48152.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 15:10:@48153.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 15:10:@48154.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 15:10:@48155.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 15:10:@48156.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 15:10:@48157.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 15:10:@48158.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 15:10:@48159.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 15:10:@48160.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 15:10:@48161.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 15:10:@48162.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 15:10:@48163.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 15:10:@48164.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 15:10:@48165.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 15:10:@48166.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 15:10:@48167.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 15:10:@48168.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 15:10:@48169.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 15:10:@48170.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 15:10:@48171.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 15:10:@48106.4]
  assign io_out_wresp_ready = _T_223 ? io_in_wresp_ready : 1'h1; // @[AXIProtocol.scala 15:10:@48087.4 AXIProtocol.scala 47:22:@48246.4]
  assign cmdSizeCounter_clock = clock; // @[:@48198.4]
  assign cmdSizeCounter_reset = reset; // @[:@48199.4]
  assign cmdSizeCounter_io_reset = lastCmd & cmdIssue; // @[AXIProtocol.scala 40:27:@48231.4]
  assign cmdSizeCounter_io_enable = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 41:28:@48232.4]
  assign cmdSizeCounter_io_stride = 32'h100; // @[AXIProtocol.scala 42:28:@48233.4]
endmodule
module AXICmdIssue( // @[:@48266.2]
  input         clock, // @[:@48267.4]
  input         reset, // @[:@48268.4]
  output        io_in_cmd_ready, // @[:@48269.4]
  input         io_in_cmd_valid, // @[:@48269.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@48269.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@48269.4]
  input         io_in_cmd_bits_isWr, // @[:@48269.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@48269.4]
  output        io_in_wdata_ready, // @[:@48269.4]
  input         io_in_wdata_valid, // @[:@48269.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@48269.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@48269.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@48269.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@48269.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@48269.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@48269.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@48269.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@48269.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@48269.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@48269.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@48269.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@48269.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@48269.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@48269.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@48269.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@48269.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@48269.4]
  input         io_in_rresp_ready, // @[:@48269.4]
  input         io_in_wresp_ready, // @[:@48269.4]
  output        io_in_wresp_valid, // @[:@48269.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@48269.4]
  input         io_out_cmd_ready, // @[:@48269.4]
  output        io_out_cmd_valid, // @[:@48269.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@48269.4]
  output [31:0] io_out_cmd_bits_size, // @[:@48269.4]
  output        io_out_cmd_bits_isWr, // @[:@48269.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@48269.4]
  input         io_out_wdata_ready, // @[:@48269.4]
  output        io_out_wdata_valid, // @[:@48269.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@48269.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@48269.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@48269.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@48269.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@48269.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@48269.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@48269.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@48269.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@48269.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@48269.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@48269.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@48269.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@48269.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@48269.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@48269.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@48269.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@48269.4]
  output        io_out_wdata_bits_wlast, // @[:@48269.4]
  output        io_out_rresp_ready, // @[:@48269.4]
  output        io_out_wresp_ready, // @[:@48269.4]
  input         io_out_wresp_valid, // @[:@48269.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@48269.4]
);
  wire  wdataCounter_clock; // @[AXIProtocol.scala 59:28:@48383.4]
  wire  wdataCounter_reset; // @[AXIProtocol.scala 59:28:@48383.4]
  wire  wdataCounter_io_reset; // @[AXIProtocol.scala 59:28:@48383.4]
  wire  wdataCounter_io_enable; // @[AXIProtocol.scala 59:28:@48383.4]
  wire [31:0] wdataCounter_io_stride; // @[AXIProtocol.scala 59:28:@48383.4]
  wire [31:0] wdataCounter_io_out; // @[AXIProtocol.scala 59:28:@48383.4]
  wire [31:0] wdataCounter_io_next; // @[AXIProtocol.scala 59:28:@48383.4]
  reg  writeIssued; // @[AXIProtocol.scala 61:28:@48386.4]
  reg [31:0] _RAND_0;
  wire  dramCmdIssue; // @[AXIProtocol.scala 63:39:@48387.4]
  wire  dramWriteIssue; // @[AXIProtocol.scala 64:43:@48388.4]
  wire  _T_201; // @[AXIProtocol.scala 68:54:@48389.4]
  wire  wlast; // @[AXIProtocol.scala 68:30:@48390.4]
  wire  _T_203; // @[AXIProtocol.scala 72:28:@48396.6]
  wire  _GEN_0; // @[AXIProtocol.scala 72:40:@48397.6]
  wire  _GEN_1; // @[AXIProtocol.scala 70:15:@48392.4]
  wire  _T_208; // @[AXIProtocol.scala 84:55:@48406.4]
  wire  _T_210; // @[AXIProtocol.scala 84:44:@48407.4]
  Counter_72 wdataCounter ( // @[AXIProtocol.scala 59:28:@48383.4]
    .clock(wdataCounter_clock),
    .reset(wdataCounter_reset),
    .io_reset(wdataCounter_io_reset),
    .io_enable(wdataCounter_io_enable),
    .io_stride(wdataCounter_io_stride),
    .io_out(wdataCounter_io_out),
    .io_next(wdataCounter_io_next)
  );
  assign dramCmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 63:39:@48387.4]
  assign dramWriteIssue = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 64:43:@48388.4]
  assign _T_201 = wdataCounter_io_next == io_in_cmd_bits_size; // @[AXIProtocol.scala 68:54:@48389.4]
  assign wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 68:30:@48390.4]
  assign _T_203 = dramCmdIssue & io_in_cmd_bits_isWr; // @[AXIProtocol.scala 72:28:@48396.6]
  assign _GEN_0 = _T_203 ? 1'h1 : writeIssued; // @[AXIProtocol.scala 72:40:@48397.6]
  assign _GEN_1 = wlast ? 1'h0 : _GEN_0; // @[AXIProtocol.scala 70:15:@48392.4]
  assign _T_208 = writeIssued == 1'h0; // @[AXIProtocol.scala 84:55:@48406.4]
  assign _T_210 = io_in_cmd_bits_isWr ? _T_208 : 1'h1; // @[AXIProtocol.scala 84:44:@48407.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? wlast : dramCmdIssue; // @[AXIProtocol.scala 56:10:@48382.4 AXIProtocol.scala 81:19:@48404.4]
  assign io_in_wdata_ready = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 56:10:@48375.4 AXIProtocol.scala 82:21:@48405.4]
  assign io_in_wresp_valid = io_out_wresp_valid; // @[AXIProtocol.scala 56:10:@48272.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 56:10:@48271.4]
  assign io_out_cmd_valid = io_in_cmd_valid & _T_210; // @[AXIProtocol.scala 56:10:@48381.4 AXIProtocol.scala 84:20:@48409.4]
  assign io_out_cmd_bits_addr = io_in_cmd_bits_addr; // @[AXIProtocol.scala 56:10:@48380.4]
  assign io_out_cmd_bits_size = io_in_cmd_bits_size; // @[AXIProtocol.scala 56:10:@48379.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 56:10:@48377.4]
  assign io_out_cmd_bits_tag = io_in_cmd_bits_tag; // @[AXIProtocol.scala 56:10:@48376.4]
  assign io_out_wdata_valid = io_in_wdata_valid & writeIssued; // @[AXIProtocol.scala 56:10:@48374.4 AXIProtocol.scala 86:22:@48411.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 56:10:@48358.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 56:10:@48359.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 56:10:@48360.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 56:10:@48361.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 56:10:@48362.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 56:10:@48363.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 56:10:@48364.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 56:10:@48365.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 56:10:@48366.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 56:10:@48367.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 56:10:@48368.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 56:10:@48369.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 56:10:@48370.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 56:10:@48371.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 56:10:@48372.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 56:10:@48373.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 56:10:@48294.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 56:10:@48295.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 56:10:@48296.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 56:10:@48297.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 56:10:@48298.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 56:10:@48299.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 56:10:@48300.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 56:10:@48301.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 56:10:@48302.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 56:10:@48303.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 56:10:@48304.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 56:10:@48305.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 56:10:@48306.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 56:10:@48307.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 56:10:@48308.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 56:10:@48309.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 56:10:@48310.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 56:10:@48311.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 56:10:@48312.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 56:10:@48313.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 56:10:@48314.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 56:10:@48315.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 56:10:@48316.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 56:10:@48317.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 56:10:@48318.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 56:10:@48319.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 56:10:@48320.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 56:10:@48321.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 56:10:@48322.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 56:10:@48323.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 56:10:@48324.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 56:10:@48325.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 56:10:@48326.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 56:10:@48327.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 56:10:@48328.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 56:10:@48329.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 56:10:@48330.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 56:10:@48331.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 56:10:@48332.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 56:10:@48333.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 56:10:@48334.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 56:10:@48335.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 56:10:@48336.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 56:10:@48337.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 56:10:@48338.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 56:10:@48339.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 56:10:@48340.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 56:10:@48341.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 56:10:@48342.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 56:10:@48343.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 56:10:@48344.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 56:10:@48345.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 56:10:@48346.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 56:10:@48347.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 56:10:@48348.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 56:10:@48349.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 56:10:@48350.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 56:10:@48351.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 56:10:@48352.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 56:10:@48353.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 56:10:@48354.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 56:10:@48355.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 56:10:@48356.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 56:10:@48357.4]
  assign io_out_wdata_bits_wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 56:10:@48293.4 AXIProtocol.scala 87:27:@48412.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 56:10:@48292.4]
  assign io_out_wresp_ready = io_in_wresp_ready; // @[AXIProtocol.scala 56:10:@48273.4]
  assign wdataCounter_clock = clock; // @[:@48384.4]
  assign wdataCounter_reset = reset; // @[:@48385.4]
  assign wdataCounter_io_reset = dramWriteIssue & _T_201; // @[AXIProtocol.scala 76:25:@48400.4]
  assign wdataCounter_io_enable = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 77:26:@48401.4]
  assign wdataCounter_io_stride = 32'h1; // @[AXIProtocol.scala 78:26:@48402.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeIssued = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      writeIssued <= 1'h0;
    end else begin
      if (wlast) begin
        writeIssued <= 1'h0;
      end else begin
        if (_T_203) begin
          writeIssued <= 1'h1;
        end
      end
    end
  end
endmodule
module DRAMArbiter( // @[:@48414.2]
  input         clock, // @[:@48415.4]
  input         reset, // @[:@48416.4]
  input         io_enable, // @[:@48417.4]
  output        io_app_stores_0_cmd_ready, // @[:@48417.4]
  input         io_app_stores_0_cmd_valid, // @[:@48417.4]
  input  [63:0] io_app_stores_0_cmd_bits_addr, // @[:@48417.4]
  input  [31:0] io_app_stores_0_cmd_bits_size, // @[:@48417.4]
  output        io_app_stores_0_data_ready, // @[:@48417.4]
  input         io_app_stores_0_data_valid, // @[:@48417.4]
  input  [31:0] io_app_stores_0_data_bits_wdata_0, // @[:@48417.4]
  input         io_app_stores_0_data_bits_wstrb, // @[:@48417.4]
  input         io_app_stores_0_wresp_ready, // @[:@48417.4]
  output        io_app_stores_0_wresp_valid, // @[:@48417.4]
  output        io_app_stores_0_wresp_bits, // @[:@48417.4]
  input         io_dram_cmd_ready, // @[:@48417.4]
  output        io_dram_cmd_valid, // @[:@48417.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@48417.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@48417.4]
  output        io_dram_cmd_bits_isWr, // @[:@48417.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@48417.4]
  input         io_dram_wdata_ready, // @[:@48417.4]
  output        io_dram_wdata_valid, // @[:@48417.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@48417.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@48417.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@48417.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@48417.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@48417.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@48417.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@48417.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@48417.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@48417.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@48417.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@48417.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@48417.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@48417.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@48417.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@48417.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@48417.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@48417.4]
  output        io_dram_wdata_bits_wlast, // @[:@48417.4]
  output        io_dram_rresp_ready, // @[:@48417.4]
  output        io_dram_wresp_ready, // @[:@48417.4]
  input         io_dram_wresp_valid, // @[:@48417.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@48417.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@49303.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@49317.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@49545.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@49660.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@49660.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@49303.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@49317.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@49545.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@49660.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_app_stores_0_cmd_ready = StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 68:18:@49316.4]
  assign io_app_stores_0_data_ready = StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 68:18:@49312.4]
  assign io_app_stores_0_wresp_valid = StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 68:18:@49307.4]
  assign io_app_stores_0_wresp_bits = StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 68:18:@49306.4]
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@49885.4 DRAMArbiter.scala 100:23:@49888.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@49884.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@49883.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@49881.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@49880.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@49878.4 DRAMArbiter.scala 101:25:@49890.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@49862.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@49863.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@49864.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@49865.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@49866.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@49867.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@49868.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@49869.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@49870.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@49871.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@49872.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@49873.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@49874.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@49875.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@49876.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@49877.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@49798.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@49799.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@49800.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@49801.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@49802.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@49803.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@49804.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@49805.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@49806.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@49807.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@49808.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@49809.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@49810.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@49811.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@49812.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@49813.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@49814.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@49815.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@49816.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@49817.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@49818.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@49819.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@49820.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@49821.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@49822.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@49823.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@49824.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@49825.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@49826.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@49827.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@49828.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@49829.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@49830.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@49831.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@49832.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@49833.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@49834.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@49835.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@49836.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@49837.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@49838.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@49839.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@49840.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@49841.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@49842.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@49843.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@49844.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@49845.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@49846.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@49847.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@49848.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@49849.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@49850.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@49851.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@49852.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@49853.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@49854.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@49855.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@49856.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@49857.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@49858.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@49859.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@49860.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@49861.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@49797.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@49796.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@49777.4]
  assign StreamControllerStore_clock = clock; // @[:@49304.4]
  assign StreamControllerStore_reset = reset; // @[:@49305.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@49432.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@49425.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@49322.4]
  assign StreamControllerStore_io_store_cmd_valid = io_app_stores_0_cmd_valid; // @[DRAMArbiter.scala 68:18:@49315.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = io_app_stores_0_cmd_bits_addr; // @[DRAMArbiter.scala 68:18:@49314.4]
  assign StreamControllerStore_io_store_cmd_bits_size = io_app_stores_0_cmd_bits_size; // @[DRAMArbiter.scala 68:18:@49313.4]
  assign StreamControllerStore_io_store_data_valid = io_app_stores_0_data_valid; // @[DRAMArbiter.scala 68:18:@49311.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = io_app_stores_0_data_bits_wdata_0; // @[DRAMArbiter.scala 68:18:@49310.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = io_app_stores_0_data_bits_wstrb; // @[DRAMArbiter.scala 68:18:@49309.4]
  assign StreamControllerStore_io_store_wresp_ready = io_app_stores_0_wresp_ready; // @[DRAMArbiter.scala 68:18:@49308.4]
  assign StreamArbiter_clock = clock; // @[:@49318.4]
  assign StreamArbiter_reset = reset; // @[:@49319.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@49543.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@49542.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@49541.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@49539.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@49538.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@49536.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@49520.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@49521.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@49522.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@49523.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@49524.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@49525.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@49526.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@49527.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@49528.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@49529.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@49530.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@49531.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@49532.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@49533.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@49534.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@49535.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@49456.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@49457.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@49458.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@49459.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@49460.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@49461.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@49462.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@49463.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@49464.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@49465.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@49466.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@49467.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@49468.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@49469.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@49470.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@49471.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@49472.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@49473.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@49474.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@49475.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@49476.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@49477.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@49478.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@49479.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@49480.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@49481.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@49482.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@49483.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@49484.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@49485.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@49486.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@49487.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@49488.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@49489.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@49490.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@49491.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@49492.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@49493.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@49494.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@49495.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@49496.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@49497.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@49498.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@49499.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@49500.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@49501.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@49502.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@49503.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@49504.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@49505.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@49506.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@49507.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@49508.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@49509.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@49510.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@49511.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@49512.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@49513.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@49514.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@49515.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@49516.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@49517.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@49518.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@49519.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@49454.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@49435.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@49659.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@49652.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@49549.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@49548.4]
  assign AXICmdSplit_clock = clock; // @[:@49546.4]
  assign AXICmdSplit_reset = reset; // @[:@49547.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@49658.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@49657.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@49656.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@49654.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@49653.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@49651.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@49635.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@49636.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@49637.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@49638.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@49639.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@49640.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@49641.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@49642.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@49643.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@49644.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@49645.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@49646.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@49647.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@49648.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@49649.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@49650.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@49571.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@49572.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@49573.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@49574.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@49575.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@49576.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@49577.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@49578.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@49579.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@49580.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@49581.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@49582.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@49583.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@49584.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@49585.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@49586.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@49587.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@49588.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@49589.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@49590.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@49591.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@49592.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@49593.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@49594.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@49595.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@49596.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@49597.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@49598.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@49599.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@49600.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@49601.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@49602.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@49603.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@49604.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@49605.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@49606.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@49607.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@49608.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@49609.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@49610.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@49611.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@49612.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@49613.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@49614.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@49615.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@49616.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@49617.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@49618.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@49619.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@49620.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@49621.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@49622.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@49623.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@49624.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@49625.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@49626.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@49627.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@49628.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@49629.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@49630.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@49631.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@49632.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@49633.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@49634.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@49569.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@49550.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@49774.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@49767.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@49664.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@49663.4]
  assign AXICmdIssue_clock = clock; // @[:@49661.4]
  assign AXICmdIssue_reset = reset; // @[:@49662.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@49773.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@49772.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@49771.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@49769.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@49768.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@49766.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@49750.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@49751.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@49752.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@49753.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@49754.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@49755.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@49756.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@49757.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@49758.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@49759.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@49760.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@49761.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@49762.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@49763.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@49764.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@49765.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@49686.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@49687.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@49688.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@49689.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@49690.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@49691.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@49692.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@49693.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@49694.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@49695.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@49696.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@49697.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@49698.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@49699.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@49700.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@49701.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@49702.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@49703.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@49704.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@49705.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@49706.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@49707.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@49708.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@49709.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@49710.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@49711.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@49712.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@49713.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@49714.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@49715.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@49716.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@49717.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@49718.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@49719.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@49720.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@49721.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@49722.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@49723.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@49724.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@49725.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@49726.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@49727.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@49728.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@49729.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@49730.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@49731.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@49732.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@49733.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@49734.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@49735.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@49736.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@49737.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@49738.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@49739.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@49740.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@49741.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@49742.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@49743.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@49744.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@49745.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@49746.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@49747.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@49748.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@49749.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@49684.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@49665.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@49886.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@49879.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@49776.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@49775.4]
endmodule
module DRAMArbiter_1( // @[:@64115.2]
  input         clock, // @[:@64116.4]
  input         reset, // @[:@64117.4]
  input         io_enable, // @[:@64118.4]
  input         io_dram_cmd_ready, // @[:@64118.4]
  output        io_dram_cmd_valid, // @[:@64118.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@64118.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@64118.4]
  output        io_dram_cmd_bits_isWr, // @[:@64118.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@64118.4]
  input         io_dram_wdata_ready, // @[:@64118.4]
  output        io_dram_wdata_valid, // @[:@64118.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@64118.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@64118.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@64118.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@64118.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@64118.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@64118.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@64118.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@64118.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@64118.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@64118.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@64118.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@64118.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@64118.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@64118.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@64118.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@64118.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@64118.4]
  output        io_dram_wdata_bits_wlast, // @[:@64118.4]
  output        io_dram_rresp_ready, // @[:@64118.4]
  output        io_dram_wresp_ready, // @[:@64118.4]
  input         io_dram_wresp_valid, // @[:@64118.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@64118.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@65004.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@65018.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@65246.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@65361.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@65361.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@65004.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@65018.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@65246.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@65361.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@65586.4 DRAMArbiter.scala 100:23:@65589.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@65585.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@65584.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@65582.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@65581.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@65579.4 DRAMArbiter.scala 101:25:@65591.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@65563.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@65564.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@65565.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@65566.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@65567.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@65568.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@65569.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@65570.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@65571.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@65572.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@65573.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@65574.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@65575.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@65576.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@65577.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@65578.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@65499.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@65500.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@65501.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@65502.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@65503.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@65504.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@65505.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@65506.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@65507.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@65508.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@65509.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@65510.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@65511.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@65512.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@65513.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@65514.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@65515.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@65516.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@65517.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@65518.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@65519.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@65520.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@65521.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@65522.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@65523.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@65524.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@65525.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@65526.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@65527.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@65528.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@65529.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@65530.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@65531.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@65532.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@65533.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@65534.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@65535.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@65536.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@65537.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@65538.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@65539.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@65540.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@65541.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@65542.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@65543.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@65544.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@65545.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@65546.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@65547.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@65548.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@65549.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@65550.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@65551.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@65552.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@65553.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@65554.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@65555.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@65556.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@65557.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@65558.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@65559.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@65560.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@65561.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@65562.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@65498.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@65497.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@65478.4]
  assign StreamControllerStore_clock = clock; // @[:@65005.4]
  assign StreamControllerStore_reset = reset; // @[:@65006.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@65133.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@65126.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@65023.4]
  assign StreamControllerStore_io_store_cmd_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@65016.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = 64'h0; // @[DRAMArbiter.scala 68:18:@65015.4]
  assign StreamControllerStore_io_store_cmd_bits_size = 32'h0; // @[DRAMArbiter.scala 68:18:@65014.4]
  assign StreamControllerStore_io_store_data_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@65012.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = 32'h0; // @[DRAMArbiter.scala 68:18:@65011.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = 1'h0; // @[DRAMArbiter.scala 68:18:@65010.4]
  assign StreamControllerStore_io_store_wresp_ready = 1'h0; // @[DRAMArbiter.scala 68:18:@65009.4]
  assign StreamArbiter_clock = clock; // @[:@65019.4]
  assign StreamArbiter_reset = reset; // @[:@65020.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@65244.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@65243.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@65242.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@65240.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@65239.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@65237.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@65221.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@65222.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@65223.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@65224.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@65225.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@65226.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@65227.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@65228.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@65229.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@65230.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@65231.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@65232.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@65233.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@65234.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@65235.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@65236.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@65157.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@65158.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@65159.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@65160.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@65161.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@65162.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@65163.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@65164.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@65165.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@65166.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@65167.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@65168.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@65169.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@65170.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@65171.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@65172.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@65173.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@65174.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@65175.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@65176.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@65177.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@65178.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@65179.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@65180.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@65181.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@65182.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@65183.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@65184.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@65185.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@65186.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@65187.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@65188.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@65189.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@65190.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@65191.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@65192.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@65193.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@65194.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@65195.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@65196.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@65197.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@65198.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@65199.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@65200.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@65201.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@65202.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@65203.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@65204.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@65205.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@65206.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@65207.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@65208.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@65209.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@65210.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@65211.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@65212.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@65213.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@65214.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@65215.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@65216.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@65217.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@65218.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@65219.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@65220.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@65155.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@65136.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@65360.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@65353.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@65250.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@65249.4]
  assign AXICmdSplit_clock = clock; // @[:@65247.4]
  assign AXICmdSplit_reset = reset; // @[:@65248.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@65359.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@65358.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@65357.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@65355.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@65354.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@65352.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@65336.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@65337.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@65338.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@65339.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@65340.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@65341.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@65342.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@65343.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@65344.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@65345.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@65346.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@65347.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@65348.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@65349.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@65350.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@65351.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@65272.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@65273.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@65274.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@65275.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@65276.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@65277.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@65278.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@65279.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@65280.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@65281.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@65282.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@65283.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@65284.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@65285.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@65286.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@65287.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@65288.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@65289.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@65290.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@65291.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@65292.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@65293.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@65294.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@65295.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@65296.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@65297.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@65298.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@65299.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@65300.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@65301.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@65302.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@65303.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@65304.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@65305.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@65306.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@65307.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@65308.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@65309.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@65310.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@65311.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@65312.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@65313.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@65314.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@65315.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@65316.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@65317.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@65318.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@65319.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@65320.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@65321.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@65322.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@65323.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@65324.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@65325.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@65326.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@65327.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@65328.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@65329.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@65330.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@65331.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@65332.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@65333.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@65334.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@65335.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@65270.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@65251.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@65475.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@65468.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@65365.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@65364.4]
  assign AXICmdIssue_clock = clock; // @[:@65362.4]
  assign AXICmdIssue_reset = reset; // @[:@65363.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@65474.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@65473.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@65472.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@65470.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@65469.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@65467.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@65451.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@65452.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@65453.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@65454.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@65455.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@65456.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@65457.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@65458.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@65459.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@65460.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@65461.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@65462.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@65463.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@65464.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@65465.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@65466.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@65387.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@65388.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@65389.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@65390.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@65391.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@65392.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@65393.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@65394.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@65395.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@65396.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@65397.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@65398.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@65399.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@65400.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@65401.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@65402.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@65403.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@65404.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@65405.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@65406.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@65407.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@65408.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@65409.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@65410.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@65411.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@65412.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@65413.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@65414.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@65415.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@65416.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@65417.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@65418.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@65419.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@65420.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@65421.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@65422.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@65423.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@65424.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@65425.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@65426.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@65427.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@65428.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@65429.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@65430.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@65431.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@65432.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@65433.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@65434.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@65435.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@65436.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@65437.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@65438.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@65439.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@65440.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@65441.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@65442.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@65443.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@65444.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@65445.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@65446.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@65447.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@65448.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@65449.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@65450.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@65385.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@65366.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@65587.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@65580.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@65477.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@65476.4]
endmodule
module DRAMHeap( // @[:@96223.2]
  input         io_accel_0_req_valid, // @[:@96226.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@96226.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@96226.4]
  output        io_accel_0_resp_valid, // @[:@96226.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@96226.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@96226.4]
  output        io_host_0_req_valid, // @[:@96226.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@96226.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@96226.4]
  input         io_host_0_resp_valid, // @[:@96226.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@96226.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@96226.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@96233.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@96235.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@96234.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@96230.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@96229.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@96228.4]
endmodule
module RetimeWrapper_333( // @[:@96249.2]
  input         clock, // @[:@96250.4]
  input         reset, // @[:@96251.4]
  input         io_flow, // @[:@96252.4]
  input  [63:0] io_in, // @[:@96252.4]
  output [63:0] io_out // @[:@96252.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@96254.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@96254.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@96254.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@96254.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@96254.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@96254.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@96254.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@96267.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@96266.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@96265.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@96264.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@96263.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@96261.4]
endmodule
module FringeFF( // @[:@96269.2]
  input         clock, // @[:@96270.4]
  input         reset, // @[:@96271.4]
  input  [63:0] io_in, // @[:@96272.4]
  input         io_reset, // @[:@96272.4]
  output [63:0] io_out, // @[:@96272.4]
  input         io_enable // @[:@96272.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@96275.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@96275.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@96275.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@96275.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@96275.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@96280.4 package.scala 96:25:@96281.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@96286.6]
  RetimeWrapper_333 RetimeWrapper ( // @[package.scala 93:22:@96275.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@96280.4 package.scala 96:25:@96281.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@96286.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@96292.4]
  assign RetimeWrapper_clock = clock; // @[:@96276.4]
  assign RetimeWrapper_reset = reset; // @[:@96277.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@96279.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@96278.4]
endmodule
module MuxN( // @[:@124908.2]
  input  [63:0] io_ins_0, // @[:@124911.4]
  input  [63:0] io_ins_1, // @[:@124911.4]
  input  [63:0] io_ins_2, // @[:@124911.4]
  input  [63:0] io_ins_3, // @[:@124911.4]
  input  [63:0] io_ins_4, // @[:@124911.4]
  input  [63:0] io_ins_5, // @[:@124911.4]
  input  [63:0] io_ins_6, // @[:@124911.4]
  input  [63:0] io_ins_7, // @[:@124911.4]
  input  [63:0] io_ins_8, // @[:@124911.4]
  input  [63:0] io_ins_9, // @[:@124911.4]
  input  [63:0] io_ins_10, // @[:@124911.4]
  input  [63:0] io_ins_11, // @[:@124911.4]
  input  [63:0] io_ins_12, // @[:@124911.4]
  input  [63:0] io_ins_13, // @[:@124911.4]
  input  [63:0] io_ins_14, // @[:@124911.4]
  input  [63:0] io_ins_15, // @[:@124911.4]
  input  [63:0] io_ins_16, // @[:@124911.4]
  input  [63:0] io_ins_17, // @[:@124911.4]
  input  [63:0] io_ins_18, // @[:@124911.4]
  input  [63:0] io_ins_19, // @[:@124911.4]
  input  [63:0] io_ins_20, // @[:@124911.4]
  input  [63:0] io_ins_21, // @[:@124911.4]
  input  [63:0] io_ins_22, // @[:@124911.4]
  input  [63:0] io_ins_23, // @[:@124911.4]
  input  [63:0] io_ins_24, // @[:@124911.4]
  input  [63:0] io_ins_25, // @[:@124911.4]
  input  [63:0] io_ins_26, // @[:@124911.4]
  input  [63:0] io_ins_27, // @[:@124911.4]
  input  [63:0] io_ins_28, // @[:@124911.4]
  input  [63:0] io_ins_29, // @[:@124911.4]
  input  [63:0] io_ins_30, // @[:@124911.4]
  input  [63:0] io_ins_31, // @[:@124911.4]
  input  [63:0] io_ins_32, // @[:@124911.4]
  input  [63:0] io_ins_33, // @[:@124911.4]
  input  [63:0] io_ins_34, // @[:@124911.4]
  input  [63:0] io_ins_35, // @[:@124911.4]
  input  [63:0] io_ins_36, // @[:@124911.4]
  input  [63:0] io_ins_37, // @[:@124911.4]
  input  [63:0] io_ins_38, // @[:@124911.4]
  input  [63:0] io_ins_39, // @[:@124911.4]
  input  [63:0] io_ins_40, // @[:@124911.4]
  input  [63:0] io_ins_41, // @[:@124911.4]
  input  [63:0] io_ins_42, // @[:@124911.4]
  input  [63:0] io_ins_43, // @[:@124911.4]
  input  [63:0] io_ins_44, // @[:@124911.4]
  input  [63:0] io_ins_45, // @[:@124911.4]
  input  [63:0] io_ins_46, // @[:@124911.4]
  input  [63:0] io_ins_47, // @[:@124911.4]
  input  [63:0] io_ins_48, // @[:@124911.4]
  input  [63:0] io_ins_49, // @[:@124911.4]
  input  [63:0] io_ins_50, // @[:@124911.4]
  input  [63:0] io_ins_51, // @[:@124911.4]
  input  [63:0] io_ins_52, // @[:@124911.4]
  input  [63:0] io_ins_53, // @[:@124911.4]
  input  [63:0] io_ins_54, // @[:@124911.4]
  input  [63:0] io_ins_55, // @[:@124911.4]
  input  [63:0] io_ins_56, // @[:@124911.4]
  input  [63:0] io_ins_57, // @[:@124911.4]
  input  [63:0] io_ins_58, // @[:@124911.4]
  input  [63:0] io_ins_59, // @[:@124911.4]
  input  [63:0] io_ins_60, // @[:@124911.4]
  input  [63:0] io_ins_61, // @[:@124911.4]
  input  [63:0] io_ins_62, // @[:@124911.4]
  input  [63:0] io_ins_63, // @[:@124911.4]
  input  [63:0] io_ins_64, // @[:@124911.4]
  input  [63:0] io_ins_65, // @[:@124911.4]
  input  [63:0] io_ins_66, // @[:@124911.4]
  input  [63:0] io_ins_67, // @[:@124911.4]
  input  [63:0] io_ins_68, // @[:@124911.4]
  input  [63:0] io_ins_69, // @[:@124911.4]
  input  [63:0] io_ins_70, // @[:@124911.4]
  input  [63:0] io_ins_71, // @[:@124911.4]
  input  [63:0] io_ins_72, // @[:@124911.4]
  input  [63:0] io_ins_73, // @[:@124911.4]
  input  [63:0] io_ins_74, // @[:@124911.4]
  input  [63:0] io_ins_75, // @[:@124911.4]
  input  [63:0] io_ins_76, // @[:@124911.4]
  input  [63:0] io_ins_77, // @[:@124911.4]
  input  [63:0] io_ins_78, // @[:@124911.4]
  input  [63:0] io_ins_79, // @[:@124911.4]
  input  [63:0] io_ins_80, // @[:@124911.4]
  input  [63:0] io_ins_81, // @[:@124911.4]
  input  [63:0] io_ins_82, // @[:@124911.4]
  input  [63:0] io_ins_83, // @[:@124911.4]
  input  [63:0] io_ins_84, // @[:@124911.4]
  input  [63:0] io_ins_85, // @[:@124911.4]
  input  [63:0] io_ins_86, // @[:@124911.4]
  input  [63:0] io_ins_87, // @[:@124911.4]
  input  [63:0] io_ins_88, // @[:@124911.4]
  input  [63:0] io_ins_89, // @[:@124911.4]
  input  [63:0] io_ins_90, // @[:@124911.4]
  input  [63:0] io_ins_91, // @[:@124911.4]
  input  [63:0] io_ins_92, // @[:@124911.4]
  input  [63:0] io_ins_93, // @[:@124911.4]
  input  [63:0] io_ins_94, // @[:@124911.4]
  input  [63:0] io_ins_95, // @[:@124911.4]
  input  [63:0] io_ins_96, // @[:@124911.4]
  input  [63:0] io_ins_97, // @[:@124911.4]
  input  [63:0] io_ins_98, // @[:@124911.4]
  input  [63:0] io_ins_99, // @[:@124911.4]
  input  [63:0] io_ins_100, // @[:@124911.4]
  input  [63:0] io_ins_101, // @[:@124911.4]
  input  [63:0] io_ins_102, // @[:@124911.4]
  input  [63:0] io_ins_103, // @[:@124911.4]
  input  [63:0] io_ins_104, // @[:@124911.4]
  input  [63:0] io_ins_105, // @[:@124911.4]
  input  [63:0] io_ins_106, // @[:@124911.4]
  input  [63:0] io_ins_107, // @[:@124911.4]
  input  [63:0] io_ins_108, // @[:@124911.4]
  input  [63:0] io_ins_109, // @[:@124911.4]
  input  [63:0] io_ins_110, // @[:@124911.4]
  input  [63:0] io_ins_111, // @[:@124911.4]
  input  [63:0] io_ins_112, // @[:@124911.4]
  input  [63:0] io_ins_113, // @[:@124911.4]
  input  [63:0] io_ins_114, // @[:@124911.4]
  input  [63:0] io_ins_115, // @[:@124911.4]
  input  [63:0] io_ins_116, // @[:@124911.4]
  input  [63:0] io_ins_117, // @[:@124911.4]
  input  [63:0] io_ins_118, // @[:@124911.4]
  input  [63:0] io_ins_119, // @[:@124911.4]
  input  [63:0] io_ins_120, // @[:@124911.4]
  input  [63:0] io_ins_121, // @[:@124911.4]
  input  [63:0] io_ins_122, // @[:@124911.4]
  input  [63:0] io_ins_123, // @[:@124911.4]
  input  [63:0] io_ins_124, // @[:@124911.4]
  input  [63:0] io_ins_125, // @[:@124911.4]
  input  [63:0] io_ins_126, // @[:@124911.4]
  input  [63:0] io_ins_127, // @[:@124911.4]
  input  [63:0] io_ins_128, // @[:@124911.4]
  input  [63:0] io_ins_129, // @[:@124911.4]
  input  [63:0] io_ins_130, // @[:@124911.4]
  input  [63:0] io_ins_131, // @[:@124911.4]
  input  [63:0] io_ins_132, // @[:@124911.4]
  input  [63:0] io_ins_133, // @[:@124911.4]
  input  [63:0] io_ins_134, // @[:@124911.4]
  input  [63:0] io_ins_135, // @[:@124911.4]
  input  [63:0] io_ins_136, // @[:@124911.4]
  input  [63:0] io_ins_137, // @[:@124911.4]
  input  [63:0] io_ins_138, // @[:@124911.4]
  input  [63:0] io_ins_139, // @[:@124911.4]
  input  [63:0] io_ins_140, // @[:@124911.4]
  input  [63:0] io_ins_141, // @[:@124911.4]
  input  [63:0] io_ins_142, // @[:@124911.4]
  input  [63:0] io_ins_143, // @[:@124911.4]
  input  [63:0] io_ins_144, // @[:@124911.4]
  input  [63:0] io_ins_145, // @[:@124911.4]
  input  [63:0] io_ins_146, // @[:@124911.4]
  input  [63:0] io_ins_147, // @[:@124911.4]
  input  [63:0] io_ins_148, // @[:@124911.4]
  input  [63:0] io_ins_149, // @[:@124911.4]
  input  [63:0] io_ins_150, // @[:@124911.4]
  input  [63:0] io_ins_151, // @[:@124911.4]
  input  [63:0] io_ins_152, // @[:@124911.4]
  input  [63:0] io_ins_153, // @[:@124911.4]
  input  [63:0] io_ins_154, // @[:@124911.4]
  input  [63:0] io_ins_155, // @[:@124911.4]
  input  [63:0] io_ins_156, // @[:@124911.4]
  input  [63:0] io_ins_157, // @[:@124911.4]
  input  [63:0] io_ins_158, // @[:@124911.4]
  input  [63:0] io_ins_159, // @[:@124911.4]
  input  [63:0] io_ins_160, // @[:@124911.4]
  input  [63:0] io_ins_161, // @[:@124911.4]
  input  [63:0] io_ins_162, // @[:@124911.4]
  input  [63:0] io_ins_163, // @[:@124911.4]
  input  [63:0] io_ins_164, // @[:@124911.4]
  input  [63:0] io_ins_165, // @[:@124911.4]
  input  [63:0] io_ins_166, // @[:@124911.4]
  input  [63:0] io_ins_167, // @[:@124911.4]
  input  [63:0] io_ins_168, // @[:@124911.4]
  input  [63:0] io_ins_169, // @[:@124911.4]
  input  [63:0] io_ins_170, // @[:@124911.4]
  input  [63:0] io_ins_171, // @[:@124911.4]
  input  [63:0] io_ins_172, // @[:@124911.4]
  input  [63:0] io_ins_173, // @[:@124911.4]
  input  [63:0] io_ins_174, // @[:@124911.4]
  input  [63:0] io_ins_175, // @[:@124911.4]
  input  [63:0] io_ins_176, // @[:@124911.4]
  input  [63:0] io_ins_177, // @[:@124911.4]
  input  [63:0] io_ins_178, // @[:@124911.4]
  input  [63:0] io_ins_179, // @[:@124911.4]
  input  [63:0] io_ins_180, // @[:@124911.4]
  input  [63:0] io_ins_181, // @[:@124911.4]
  input  [63:0] io_ins_182, // @[:@124911.4]
  input  [63:0] io_ins_183, // @[:@124911.4]
  input  [63:0] io_ins_184, // @[:@124911.4]
  input  [63:0] io_ins_185, // @[:@124911.4]
  input  [63:0] io_ins_186, // @[:@124911.4]
  input  [63:0] io_ins_187, // @[:@124911.4]
  input  [63:0] io_ins_188, // @[:@124911.4]
  input  [63:0] io_ins_189, // @[:@124911.4]
  input  [63:0] io_ins_190, // @[:@124911.4]
  input  [63:0] io_ins_191, // @[:@124911.4]
  input  [63:0] io_ins_192, // @[:@124911.4]
  input  [63:0] io_ins_193, // @[:@124911.4]
  input  [63:0] io_ins_194, // @[:@124911.4]
  input  [63:0] io_ins_195, // @[:@124911.4]
  input  [63:0] io_ins_196, // @[:@124911.4]
  input  [63:0] io_ins_197, // @[:@124911.4]
  input  [63:0] io_ins_198, // @[:@124911.4]
  input  [63:0] io_ins_199, // @[:@124911.4]
  input  [63:0] io_ins_200, // @[:@124911.4]
  input  [63:0] io_ins_201, // @[:@124911.4]
  input  [63:0] io_ins_202, // @[:@124911.4]
  input  [63:0] io_ins_203, // @[:@124911.4]
  input  [63:0] io_ins_204, // @[:@124911.4]
  input  [63:0] io_ins_205, // @[:@124911.4]
  input  [63:0] io_ins_206, // @[:@124911.4]
  input  [63:0] io_ins_207, // @[:@124911.4]
  input  [63:0] io_ins_208, // @[:@124911.4]
  input  [63:0] io_ins_209, // @[:@124911.4]
  input  [63:0] io_ins_210, // @[:@124911.4]
  input  [63:0] io_ins_211, // @[:@124911.4]
  input  [63:0] io_ins_212, // @[:@124911.4]
  input  [63:0] io_ins_213, // @[:@124911.4]
  input  [63:0] io_ins_214, // @[:@124911.4]
  input  [63:0] io_ins_215, // @[:@124911.4]
  input  [63:0] io_ins_216, // @[:@124911.4]
  input  [63:0] io_ins_217, // @[:@124911.4]
  input  [63:0] io_ins_218, // @[:@124911.4]
  input  [63:0] io_ins_219, // @[:@124911.4]
  input  [63:0] io_ins_220, // @[:@124911.4]
  input  [63:0] io_ins_221, // @[:@124911.4]
  input  [63:0] io_ins_222, // @[:@124911.4]
  input  [63:0] io_ins_223, // @[:@124911.4]
  input  [63:0] io_ins_224, // @[:@124911.4]
  input  [63:0] io_ins_225, // @[:@124911.4]
  input  [63:0] io_ins_226, // @[:@124911.4]
  input  [63:0] io_ins_227, // @[:@124911.4]
  input  [63:0] io_ins_228, // @[:@124911.4]
  input  [63:0] io_ins_229, // @[:@124911.4]
  input  [63:0] io_ins_230, // @[:@124911.4]
  input  [63:0] io_ins_231, // @[:@124911.4]
  input  [63:0] io_ins_232, // @[:@124911.4]
  input  [63:0] io_ins_233, // @[:@124911.4]
  input  [63:0] io_ins_234, // @[:@124911.4]
  input  [63:0] io_ins_235, // @[:@124911.4]
  input  [63:0] io_ins_236, // @[:@124911.4]
  input  [63:0] io_ins_237, // @[:@124911.4]
  input  [63:0] io_ins_238, // @[:@124911.4]
  input  [63:0] io_ins_239, // @[:@124911.4]
  input  [63:0] io_ins_240, // @[:@124911.4]
  input  [63:0] io_ins_241, // @[:@124911.4]
  input  [63:0] io_ins_242, // @[:@124911.4]
  input  [63:0] io_ins_243, // @[:@124911.4]
  input  [63:0] io_ins_244, // @[:@124911.4]
  input  [63:0] io_ins_245, // @[:@124911.4]
  input  [63:0] io_ins_246, // @[:@124911.4]
  input  [63:0] io_ins_247, // @[:@124911.4]
  input  [63:0] io_ins_248, // @[:@124911.4]
  input  [63:0] io_ins_249, // @[:@124911.4]
  input  [63:0] io_ins_250, // @[:@124911.4]
  input  [63:0] io_ins_251, // @[:@124911.4]
  input  [63:0] io_ins_252, // @[:@124911.4]
  input  [63:0] io_ins_253, // @[:@124911.4]
  input  [63:0] io_ins_254, // @[:@124911.4]
  input  [63:0] io_ins_255, // @[:@124911.4]
  input  [63:0] io_ins_256, // @[:@124911.4]
  input  [63:0] io_ins_257, // @[:@124911.4]
  input  [63:0] io_ins_258, // @[:@124911.4]
  input  [63:0] io_ins_259, // @[:@124911.4]
  input  [63:0] io_ins_260, // @[:@124911.4]
  input  [63:0] io_ins_261, // @[:@124911.4]
  input  [63:0] io_ins_262, // @[:@124911.4]
  input  [63:0] io_ins_263, // @[:@124911.4]
  input  [63:0] io_ins_264, // @[:@124911.4]
  input  [63:0] io_ins_265, // @[:@124911.4]
  input  [63:0] io_ins_266, // @[:@124911.4]
  input  [63:0] io_ins_267, // @[:@124911.4]
  input  [63:0] io_ins_268, // @[:@124911.4]
  input  [63:0] io_ins_269, // @[:@124911.4]
  input  [63:0] io_ins_270, // @[:@124911.4]
  input  [63:0] io_ins_271, // @[:@124911.4]
  input  [63:0] io_ins_272, // @[:@124911.4]
  input  [63:0] io_ins_273, // @[:@124911.4]
  input  [63:0] io_ins_274, // @[:@124911.4]
  input  [63:0] io_ins_275, // @[:@124911.4]
  input  [63:0] io_ins_276, // @[:@124911.4]
  input  [63:0] io_ins_277, // @[:@124911.4]
  input  [63:0] io_ins_278, // @[:@124911.4]
  input  [63:0] io_ins_279, // @[:@124911.4]
  input  [63:0] io_ins_280, // @[:@124911.4]
  input  [63:0] io_ins_281, // @[:@124911.4]
  input  [63:0] io_ins_282, // @[:@124911.4]
  input  [63:0] io_ins_283, // @[:@124911.4]
  input  [63:0] io_ins_284, // @[:@124911.4]
  input  [63:0] io_ins_285, // @[:@124911.4]
  input  [63:0] io_ins_286, // @[:@124911.4]
  input  [63:0] io_ins_287, // @[:@124911.4]
  input  [63:0] io_ins_288, // @[:@124911.4]
  input  [63:0] io_ins_289, // @[:@124911.4]
  input  [63:0] io_ins_290, // @[:@124911.4]
  input  [63:0] io_ins_291, // @[:@124911.4]
  input  [63:0] io_ins_292, // @[:@124911.4]
  input  [63:0] io_ins_293, // @[:@124911.4]
  input  [63:0] io_ins_294, // @[:@124911.4]
  input  [63:0] io_ins_295, // @[:@124911.4]
  input  [63:0] io_ins_296, // @[:@124911.4]
  input  [63:0] io_ins_297, // @[:@124911.4]
  input  [63:0] io_ins_298, // @[:@124911.4]
  input  [63:0] io_ins_299, // @[:@124911.4]
  input  [63:0] io_ins_300, // @[:@124911.4]
  input  [63:0] io_ins_301, // @[:@124911.4]
  input  [63:0] io_ins_302, // @[:@124911.4]
  input  [63:0] io_ins_303, // @[:@124911.4]
  input  [63:0] io_ins_304, // @[:@124911.4]
  input  [63:0] io_ins_305, // @[:@124911.4]
  input  [63:0] io_ins_306, // @[:@124911.4]
  input  [63:0] io_ins_307, // @[:@124911.4]
  input  [63:0] io_ins_308, // @[:@124911.4]
  input  [63:0] io_ins_309, // @[:@124911.4]
  input  [63:0] io_ins_310, // @[:@124911.4]
  input  [63:0] io_ins_311, // @[:@124911.4]
  input  [63:0] io_ins_312, // @[:@124911.4]
  input  [63:0] io_ins_313, // @[:@124911.4]
  input  [63:0] io_ins_314, // @[:@124911.4]
  input  [63:0] io_ins_315, // @[:@124911.4]
  input  [63:0] io_ins_316, // @[:@124911.4]
  input  [63:0] io_ins_317, // @[:@124911.4]
  input  [63:0] io_ins_318, // @[:@124911.4]
  input  [63:0] io_ins_319, // @[:@124911.4]
  input  [63:0] io_ins_320, // @[:@124911.4]
  input  [63:0] io_ins_321, // @[:@124911.4]
  input  [63:0] io_ins_322, // @[:@124911.4]
  input  [63:0] io_ins_323, // @[:@124911.4]
  input  [63:0] io_ins_324, // @[:@124911.4]
  input  [63:0] io_ins_325, // @[:@124911.4]
  input  [63:0] io_ins_326, // @[:@124911.4]
  input  [63:0] io_ins_327, // @[:@124911.4]
  input  [63:0] io_ins_328, // @[:@124911.4]
  input  [63:0] io_ins_329, // @[:@124911.4]
  input  [63:0] io_ins_330, // @[:@124911.4]
  input  [63:0] io_ins_331, // @[:@124911.4]
  input  [63:0] io_ins_332, // @[:@124911.4]
  input  [63:0] io_ins_333, // @[:@124911.4]
  input  [63:0] io_ins_334, // @[:@124911.4]
  input  [63:0] io_ins_335, // @[:@124911.4]
  input  [63:0] io_ins_336, // @[:@124911.4]
  input  [63:0] io_ins_337, // @[:@124911.4]
  input  [63:0] io_ins_338, // @[:@124911.4]
  input  [63:0] io_ins_339, // @[:@124911.4]
  input  [63:0] io_ins_340, // @[:@124911.4]
  input  [63:0] io_ins_341, // @[:@124911.4]
  input  [63:0] io_ins_342, // @[:@124911.4]
  input  [63:0] io_ins_343, // @[:@124911.4]
  input  [63:0] io_ins_344, // @[:@124911.4]
  input  [63:0] io_ins_345, // @[:@124911.4]
  input  [63:0] io_ins_346, // @[:@124911.4]
  input  [63:0] io_ins_347, // @[:@124911.4]
  input  [63:0] io_ins_348, // @[:@124911.4]
  input  [63:0] io_ins_349, // @[:@124911.4]
  input  [63:0] io_ins_350, // @[:@124911.4]
  input  [63:0] io_ins_351, // @[:@124911.4]
  input  [63:0] io_ins_352, // @[:@124911.4]
  input  [63:0] io_ins_353, // @[:@124911.4]
  input  [63:0] io_ins_354, // @[:@124911.4]
  input  [63:0] io_ins_355, // @[:@124911.4]
  input  [63:0] io_ins_356, // @[:@124911.4]
  input  [63:0] io_ins_357, // @[:@124911.4]
  input  [63:0] io_ins_358, // @[:@124911.4]
  input  [63:0] io_ins_359, // @[:@124911.4]
  input  [63:0] io_ins_360, // @[:@124911.4]
  input  [63:0] io_ins_361, // @[:@124911.4]
  input  [63:0] io_ins_362, // @[:@124911.4]
  input  [63:0] io_ins_363, // @[:@124911.4]
  input  [63:0] io_ins_364, // @[:@124911.4]
  input  [63:0] io_ins_365, // @[:@124911.4]
  input  [63:0] io_ins_366, // @[:@124911.4]
  input  [63:0] io_ins_367, // @[:@124911.4]
  input  [63:0] io_ins_368, // @[:@124911.4]
  input  [63:0] io_ins_369, // @[:@124911.4]
  input  [63:0] io_ins_370, // @[:@124911.4]
  input  [63:0] io_ins_371, // @[:@124911.4]
  input  [63:0] io_ins_372, // @[:@124911.4]
  input  [63:0] io_ins_373, // @[:@124911.4]
  input  [63:0] io_ins_374, // @[:@124911.4]
  input  [63:0] io_ins_375, // @[:@124911.4]
  input  [63:0] io_ins_376, // @[:@124911.4]
  input  [63:0] io_ins_377, // @[:@124911.4]
  input  [63:0] io_ins_378, // @[:@124911.4]
  input  [63:0] io_ins_379, // @[:@124911.4]
  input  [63:0] io_ins_380, // @[:@124911.4]
  input  [63:0] io_ins_381, // @[:@124911.4]
  input  [63:0] io_ins_382, // @[:@124911.4]
  input  [63:0] io_ins_383, // @[:@124911.4]
  input  [63:0] io_ins_384, // @[:@124911.4]
  input  [63:0] io_ins_385, // @[:@124911.4]
  input  [63:0] io_ins_386, // @[:@124911.4]
  input  [63:0] io_ins_387, // @[:@124911.4]
  input  [63:0] io_ins_388, // @[:@124911.4]
  input  [63:0] io_ins_389, // @[:@124911.4]
  input  [63:0] io_ins_390, // @[:@124911.4]
  input  [63:0] io_ins_391, // @[:@124911.4]
  input  [63:0] io_ins_392, // @[:@124911.4]
  input  [63:0] io_ins_393, // @[:@124911.4]
  input  [63:0] io_ins_394, // @[:@124911.4]
  input  [63:0] io_ins_395, // @[:@124911.4]
  input  [63:0] io_ins_396, // @[:@124911.4]
  input  [63:0] io_ins_397, // @[:@124911.4]
  input  [63:0] io_ins_398, // @[:@124911.4]
  input  [63:0] io_ins_399, // @[:@124911.4]
  input  [63:0] io_ins_400, // @[:@124911.4]
  input  [63:0] io_ins_401, // @[:@124911.4]
  input  [63:0] io_ins_402, // @[:@124911.4]
  input  [63:0] io_ins_403, // @[:@124911.4]
  input  [63:0] io_ins_404, // @[:@124911.4]
  input  [63:0] io_ins_405, // @[:@124911.4]
  input  [63:0] io_ins_406, // @[:@124911.4]
  input  [63:0] io_ins_407, // @[:@124911.4]
  input  [63:0] io_ins_408, // @[:@124911.4]
  input  [63:0] io_ins_409, // @[:@124911.4]
  input  [63:0] io_ins_410, // @[:@124911.4]
  input  [63:0] io_ins_411, // @[:@124911.4]
  input  [63:0] io_ins_412, // @[:@124911.4]
  input  [63:0] io_ins_413, // @[:@124911.4]
  input  [63:0] io_ins_414, // @[:@124911.4]
  input  [63:0] io_ins_415, // @[:@124911.4]
  input  [63:0] io_ins_416, // @[:@124911.4]
  input  [63:0] io_ins_417, // @[:@124911.4]
  input  [63:0] io_ins_418, // @[:@124911.4]
  input  [63:0] io_ins_419, // @[:@124911.4]
  input  [63:0] io_ins_420, // @[:@124911.4]
  input  [63:0] io_ins_421, // @[:@124911.4]
  input  [63:0] io_ins_422, // @[:@124911.4]
  input  [63:0] io_ins_423, // @[:@124911.4]
  input  [63:0] io_ins_424, // @[:@124911.4]
  input  [63:0] io_ins_425, // @[:@124911.4]
  input  [63:0] io_ins_426, // @[:@124911.4]
  input  [63:0] io_ins_427, // @[:@124911.4]
  input  [63:0] io_ins_428, // @[:@124911.4]
  input  [63:0] io_ins_429, // @[:@124911.4]
  input  [63:0] io_ins_430, // @[:@124911.4]
  input  [63:0] io_ins_431, // @[:@124911.4]
  input  [63:0] io_ins_432, // @[:@124911.4]
  input  [63:0] io_ins_433, // @[:@124911.4]
  input  [63:0] io_ins_434, // @[:@124911.4]
  input  [63:0] io_ins_435, // @[:@124911.4]
  input  [63:0] io_ins_436, // @[:@124911.4]
  input  [63:0] io_ins_437, // @[:@124911.4]
  input  [63:0] io_ins_438, // @[:@124911.4]
  input  [63:0] io_ins_439, // @[:@124911.4]
  input  [63:0] io_ins_440, // @[:@124911.4]
  input  [63:0] io_ins_441, // @[:@124911.4]
  input  [63:0] io_ins_442, // @[:@124911.4]
  input  [63:0] io_ins_443, // @[:@124911.4]
  input  [63:0] io_ins_444, // @[:@124911.4]
  input  [63:0] io_ins_445, // @[:@124911.4]
  input  [63:0] io_ins_446, // @[:@124911.4]
  input  [63:0] io_ins_447, // @[:@124911.4]
  input  [63:0] io_ins_448, // @[:@124911.4]
  input  [63:0] io_ins_449, // @[:@124911.4]
  input  [63:0] io_ins_450, // @[:@124911.4]
  input  [63:0] io_ins_451, // @[:@124911.4]
  input  [63:0] io_ins_452, // @[:@124911.4]
  input  [63:0] io_ins_453, // @[:@124911.4]
  input  [63:0] io_ins_454, // @[:@124911.4]
  input  [63:0] io_ins_455, // @[:@124911.4]
  input  [63:0] io_ins_456, // @[:@124911.4]
  input  [63:0] io_ins_457, // @[:@124911.4]
  input  [63:0] io_ins_458, // @[:@124911.4]
  input  [63:0] io_ins_459, // @[:@124911.4]
  input  [63:0] io_ins_460, // @[:@124911.4]
  input  [63:0] io_ins_461, // @[:@124911.4]
  input  [63:0] io_ins_462, // @[:@124911.4]
  input  [63:0] io_ins_463, // @[:@124911.4]
  input  [63:0] io_ins_464, // @[:@124911.4]
  input  [63:0] io_ins_465, // @[:@124911.4]
  input  [63:0] io_ins_466, // @[:@124911.4]
  input  [63:0] io_ins_467, // @[:@124911.4]
  input  [63:0] io_ins_468, // @[:@124911.4]
  input  [63:0] io_ins_469, // @[:@124911.4]
  input  [63:0] io_ins_470, // @[:@124911.4]
  input  [63:0] io_ins_471, // @[:@124911.4]
  input  [63:0] io_ins_472, // @[:@124911.4]
  input  [63:0] io_ins_473, // @[:@124911.4]
  input  [63:0] io_ins_474, // @[:@124911.4]
  input  [63:0] io_ins_475, // @[:@124911.4]
  input  [63:0] io_ins_476, // @[:@124911.4]
  input  [63:0] io_ins_477, // @[:@124911.4]
  input  [63:0] io_ins_478, // @[:@124911.4]
  input  [63:0] io_ins_479, // @[:@124911.4]
  input  [63:0] io_ins_480, // @[:@124911.4]
  input  [63:0] io_ins_481, // @[:@124911.4]
  input  [63:0] io_ins_482, // @[:@124911.4]
  input  [63:0] io_ins_483, // @[:@124911.4]
  input  [63:0] io_ins_484, // @[:@124911.4]
  input  [63:0] io_ins_485, // @[:@124911.4]
  input  [63:0] io_ins_486, // @[:@124911.4]
  input  [63:0] io_ins_487, // @[:@124911.4]
  input  [63:0] io_ins_488, // @[:@124911.4]
  input  [63:0] io_ins_489, // @[:@124911.4]
  input  [63:0] io_ins_490, // @[:@124911.4]
  input  [63:0] io_ins_491, // @[:@124911.4]
  input  [63:0] io_ins_492, // @[:@124911.4]
  input  [63:0] io_ins_493, // @[:@124911.4]
  input  [63:0] io_ins_494, // @[:@124911.4]
  input  [63:0] io_ins_495, // @[:@124911.4]
  input  [63:0] io_ins_496, // @[:@124911.4]
  input  [63:0] io_ins_497, // @[:@124911.4]
  input  [63:0] io_ins_498, // @[:@124911.4]
  input  [63:0] io_ins_499, // @[:@124911.4]
  input  [63:0] io_ins_500, // @[:@124911.4]
  input  [63:0] io_ins_501, // @[:@124911.4]
  input  [63:0] io_ins_502, // @[:@124911.4]
  input  [8:0]  io_sel, // @[:@124911.4]
  output [63:0] io_out // @[:@124911.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@124913.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_1 = 9'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_2 = 9'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_3 = 9'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_4 = 9'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_5 = 9'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_6 = 9'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_7 = 9'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_8 = 9'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_9 = 9'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_10 = 9'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_11 = 9'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_12 = 9'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_13 = 9'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_14 = 9'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_15 = 9'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_16 = 9'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_17 = 9'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_18 = 9'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_19 = 9'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_20 = 9'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_21 = 9'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_22 = 9'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_23 = 9'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_24 = 9'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_25 = 9'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_26 = 9'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_27 = 9'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_28 = 9'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_29 = 9'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_30 = 9'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_31 = 9'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_32 = 9'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_33 = 9'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_34 = 9'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_35 = 9'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_36 = 9'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_37 = 9'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_38 = 9'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_39 = 9'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_40 = 9'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_41 = 9'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_42 = 9'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_43 = 9'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_44 = 9'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_45 = 9'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_46 = 9'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_47 = 9'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_48 = 9'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_49 = 9'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_50 = 9'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_51 = 9'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_52 = 9'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_53 = 9'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_54 = 9'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_55 = 9'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_56 = 9'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_57 = 9'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_58 = 9'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_59 = 9'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_60 = 9'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_61 = 9'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_62 = 9'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_63 = 9'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_64 = 9'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_65 = 9'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_66 = 9'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_67 = 9'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_68 = 9'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_69 = 9'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_70 = 9'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_71 = 9'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_72 = 9'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_73 = 9'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_74 = 9'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_75 = 9'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_76 = 9'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_77 = 9'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_78 = 9'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_79 = 9'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_80 = 9'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_81 = 9'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_82 = 9'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_83 = 9'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_84 = 9'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_85 = 9'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_86 = 9'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_87 = 9'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_88 = 9'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_89 = 9'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_90 = 9'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_91 = 9'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_92 = 9'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_93 = 9'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_94 = 9'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_95 = 9'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_96 = 9'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_97 = 9'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_98 = 9'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_99 = 9'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_100 = 9'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_101 = 9'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_102 = 9'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_103 = 9'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_104 = 9'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_105 = 9'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_106 = 9'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_107 = 9'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_108 = 9'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_109 = 9'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_110 = 9'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_111 = 9'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_112 = 9'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_113 = 9'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_114 = 9'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_115 = 9'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_116 = 9'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_117 = 9'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_118 = 9'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_119 = 9'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_120 = 9'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_121 = 9'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_122 = 9'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_123 = 9'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_124 = 9'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_125 = 9'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_126 = 9'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_127 = 9'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_128 = 9'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_129 = 9'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_130 = 9'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_131 = 9'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_132 = 9'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_133 = 9'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_134 = 9'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_135 = 9'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_136 = 9'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_137 = 9'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_138 = 9'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_139 = 9'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_140 = 9'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_141 = 9'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_142 = 9'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_143 = 9'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_144 = 9'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_145 = 9'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_146 = 9'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_147 = 9'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_148 = 9'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_149 = 9'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_150 = 9'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_151 = 9'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_152 = 9'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_153 = 9'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_154 = 9'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_155 = 9'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_156 = 9'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_157 = 9'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_158 = 9'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_159 = 9'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_160 = 9'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_161 = 9'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_162 = 9'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_163 = 9'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_164 = 9'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_165 = 9'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_166 = 9'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_167 = 9'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_168 = 9'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_169 = 9'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_170 = 9'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_171 = 9'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_172 = 9'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_173 = 9'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_174 = 9'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_175 = 9'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_176 = 9'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_177 = 9'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_178 = 9'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_179 = 9'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_180 = 9'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_181 = 9'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_182 = 9'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_183 = 9'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_184 = 9'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_185 = 9'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_186 = 9'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_187 = 9'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_188 = 9'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_189 = 9'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_190 = 9'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_191 = 9'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_192 = 9'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_193 = 9'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_194 = 9'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_195 = 9'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_196 = 9'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_197 = 9'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_198 = 9'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_199 = 9'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_200 = 9'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_201 = 9'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_202 = 9'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_203 = 9'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_204 = 9'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_205 = 9'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_206 = 9'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_207 = 9'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_208 = 9'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_209 = 9'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_210 = 9'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_211 = 9'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_212 = 9'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_213 = 9'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_214 = 9'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_215 = 9'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_216 = 9'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_217 = 9'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_218 = 9'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_219 = 9'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_220 = 9'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_221 = 9'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_222 = 9'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_223 = 9'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_224 = 9'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_225 = 9'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_226 = 9'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_227 = 9'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_228 = 9'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_229 = 9'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_230 = 9'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_231 = 9'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_232 = 9'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_233 = 9'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_234 = 9'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_235 = 9'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_236 = 9'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_237 = 9'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_238 = 9'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_239 = 9'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_240 = 9'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_241 = 9'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_242 = 9'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_243 = 9'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_244 = 9'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_245 = 9'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_246 = 9'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_247 = 9'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_248 = 9'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_249 = 9'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_250 = 9'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_251 = 9'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_252 = 9'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_253 = 9'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_254 = 9'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_255 = 9'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_256 = 9'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_257 = 9'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_258 = 9'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_259 = 9'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_260 = 9'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_261 = 9'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_262 = 9'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_263 = 9'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_264 = 9'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_265 = 9'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_266 = 9'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_267 = 9'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_268 = 9'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_269 = 9'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_270 = 9'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_271 = 9'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_272 = 9'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_273 = 9'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_274 = 9'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_275 = 9'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_276 = 9'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_277 = 9'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_278 = 9'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_279 = 9'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_280 = 9'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_281 = 9'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_282 = 9'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_283 = 9'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_284 = 9'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_285 = 9'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_286 = 9'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_287 = 9'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_288 = 9'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_289 = 9'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_290 = 9'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_291 = 9'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_292 = 9'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_293 = 9'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_294 = 9'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_295 = 9'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_296 = 9'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_297 = 9'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_298 = 9'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_299 = 9'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_300 = 9'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_301 = 9'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_302 = 9'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_303 = 9'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_304 = 9'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_305 = 9'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_306 = 9'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_307 = 9'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_308 = 9'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_309 = 9'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_310 = 9'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_311 = 9'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_312 = 9'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_313 = 9'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_314 = 9'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_315 = 9'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_316 = 9'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_317 = 9'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_318 = 9'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_319 = 9'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_320 = 9'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_321 = 9'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_322 = 9'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_323 = 9'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_324 = 9'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_325 = 9'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_326 = 9'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_327 = 9'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_328 = 9'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_329 = 9'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_330 = 9'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_331 = 9'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_332 = 9'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_333 = 9'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_334 = 9'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_335 = 9'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_336 = 9'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_337 = 9'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_338 = 9'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_339 = 9'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_340 = 9'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_341 = 9'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_342 = 9'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_343 = 9'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_344 = 9'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_345 = 9'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_346 = 9'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_347 = 9'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_348 = 9'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_349 = 9'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_350 = 9'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_351 = 9'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_352 = 9'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_353 = 9'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_354 = 9'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_355 = 9'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_356 = 9'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_357 = 9'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_358 = 9'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_359 = 9'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_360 = 9'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_361 = 9'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_362 = 9'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_363 = 9'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_364 = 9'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_365 = 9'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_366 = 9'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_367 = 9'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_368 = 9'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_369 = 9'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_370 = 9'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_371 = 9'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_372 = 9'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_373 = 9'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_374 = 9'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_375 = 9'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_376 = 9'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_377 = 9'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_378 = 9'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_379 = 9'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_380 = 9'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_381 = 9'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_382 = 9'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_383 = 9'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_384 = 9'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_385 = 9'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_386 = 9'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_387 = 9'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_388 = 9'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_389 = 9'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_390 = 9'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_391 = 9'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_392 = 9'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_393 = 9'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_394 = 9'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_395 = 9'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_396 = 9'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_397 = 9'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_398 = 9'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_399 = 9'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_400 = 9'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_401 = 9'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_402 = 9'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_403 = 9'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_404 = 9'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_405 = 9'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_406 = 9'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_407 = 9'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_408 = 9'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_409 = 9'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_410 = 9'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_411 = 9'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_412 = 9'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_413 = 9'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_414 = 9'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_415 = 9'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_416 = 9'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_417 = 9'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_418 = 9'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_419 = 9'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_420 = 9'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_421 = 9'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_422 = 9'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_423 = 9'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_424 = 9'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_425 = 9'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_426 = 9'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_427 = 9'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_428 = 9'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_429 = 9'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_430 = 9'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_431 = 9'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_432 = 9'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_433 = 9'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_434 = 9'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_435 = 9'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_436 = 9'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_437 = 9'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_438 = 9'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_439 = 9'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_440 = 9'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_441 = 9'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_442 = 9'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_443 = 9'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_444 = 9'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_445 = 9'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_446 = 9'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_447 = 9'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_448 = 9'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_449 = 9'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_450 = 9'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_451 = 9'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_452 = 9'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_453 = 9'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_454 = 9'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_455 = 9'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_456 = 9'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_457 = 9'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_458 = 9'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_459 = 9'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_460 = 9'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_461 = 9'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_462 = 9'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_463 = 9'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_464 = 9'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_465 = 9'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_466 = 9'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_467 = 9'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_468 = 9'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_469 = 9'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_470 = 9'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_471 = 9'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_472 = 9'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_473 = 9'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_474 = 9'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_475 = 9'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_476 = 9'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_477 = 9'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_478 = 9'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_479 = 9'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_480 = 9'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_481 = 9'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_482 = 9'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_483 = 9'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_484 = 9'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_485 = 9'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_486 = 9'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_487 = 9'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_488 = 9'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_489 = 9'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_490 = 9'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_491 = 9'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_492 = 9'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_493 = 9'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_494 = 9'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_495 = 9'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_496 = 9'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_497 = 9'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_498 = 9'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_499 = 9'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_500 = 9'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@124913.4]
  assign _GEN_501 = 9'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@124913.4]
  assign io_out = 9'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@124913.4]
endmodule
module RegFile( // @[:@124915.2]
  input         clock, // @[:@124916.4]
  input         reset, // @[:@124917.4]
  input  [31:0] io_raddr, // @[:@124918.4]
  input         io_wen, // @[:@124918.4]
  input  [31:0] io_waddr, // @[:@124918.4]
  input  [63:0] io_wdata, // @[:@124918.4]
  output [63:0] io_rdata, // @[:@124918.4]
  input         io_reset, // @[:@124918.4]
  output [63:0] io_argIns_0, // @[:@124918.4]
  output [63:0] io_argIns_1, // @[:@124918.4]
  output [63:0] io_argIns_2, // @[:@124918.4]
  output [63:0] io_argIns_3, // @[:@124918.4]
  input         io_argOuts_0_valid, // @[:@124918.4]
  input  [63:0] io_argOuts_0_bits, // @[:@124918.4]
  input         io_argOuts_1_valid, // @[:@124918.4]
  input  [63:0] io_argOuts_1_bits // @[:@124918.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@126928.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@126928.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@126928.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@126928.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@126928.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@126928.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@126940.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@126940.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@126940.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@126940.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@126940.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@126940.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@126959.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@126959.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@126959.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@126959.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@126959.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@126959.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@126971.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@126971.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@126971.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@126971.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@126971.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@126971.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@126983.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@126983.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@126983.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@126983.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@126983.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@126983.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@126997.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@126997.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@126997.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@126997.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@126997.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@126997.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@127011.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@127011.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@127011.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@127011.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@127011.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@127011.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@127025.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@127025.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@127025.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@127025.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@127025.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@127025.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@127039.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@127039.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@127039.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@127039.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@127039.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@127039.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@127053.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@127053.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@127053.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@127053.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@127053.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@127053.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@127067.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@127067.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@127067.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@127067.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@127067.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@127067.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@127081.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@127081.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@127081.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@127081.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@127081.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@127081.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@127095.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@127095.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@127095.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@127095.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@127095.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@127095.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@127109.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@127109.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@127109.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@127109.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@127109.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@127109.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@127123.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@127123.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@127123.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@127123.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@127123.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@127123.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@127137.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@127137.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@127137.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@127137.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@127137.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@127137.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@127151.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@127151.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@127151.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@127151.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@127151.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@127151.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@127165.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@127165.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@127165.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@127165.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@127165.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@127165.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@127179.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@127179.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@127179.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@127179.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@127179.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@127179.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@127193.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@127193.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@127193.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@127193.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@127193.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@127193.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@127207.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@127207.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@127207.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@127207.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@127207.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@127207.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@127221.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@127221.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@127221.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@127221.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@127221.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@127221.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@127235.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@127235.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@127235.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@127235.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@127235.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@127235.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@127249.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@127249.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@127249.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@127249.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@127249.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@127249.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@127263.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@127263.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@127263.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@127263.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@127263.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@127263.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@127277.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@127277.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@127277.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@127277.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@127277.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@127277.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@127291.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@127291.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@127291.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@127291.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@127291.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@127291.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@127305.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@127305.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@127305.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@127305.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@127305.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@127305.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@127319.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@127319.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@127319.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@127319.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@127319.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@127319.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@127333.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@127333.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@127333.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@127333.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@127333.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@127333.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@127347.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@127347.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@127347.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@127347.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@127347.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@127347.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@127361.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@127361.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@127361.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@127361.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@127361.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@127361.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@127375.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@127375.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@127375.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@127375.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@127375.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@127375.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@127389.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@127389.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@127389.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@127389.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@127389.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@127389.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@127403.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@127403.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@127403.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@127403.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@127403.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@127403.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@127417.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@127417.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@127417.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@127417.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@127417.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@127417.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@127431.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@127431.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@127431.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@127431.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@127431.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@127431.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@127445.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@127445.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@127445.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@127445.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@127445.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@127445.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@127459.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@127459.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@127459.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@127459.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@127459.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@127459.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@127473.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@127473.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@127473.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@127473.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@127473.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@127473.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@127487.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@127487.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@127487.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@127487.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@127487.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@127487.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@127501.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@127501.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@127501.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@127501.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@127501.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@127501.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@127515.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@127515.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@127515.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@127515.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@127515.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@127515.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@127529.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@127529.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@127529.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@127529.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@127529.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@127529.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@127543.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@127543.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@127543.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@127543.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@127543.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@127543.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@127557.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@127557.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@127557.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@127557.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@127557.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@127557.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@127571.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@127571.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@127571.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@127571.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@127571.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@127571.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@127585.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@127585.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@127585.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@127585.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@127585.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@127585.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@127599.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@127599.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@127599.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@127599.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@127599.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@127599.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@127613.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@127613.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@127613.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@127613.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@127613.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@127613.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@127627.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@127627.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@127627.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@127627.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@127627.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@127627.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@127641.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@127641.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@127641.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@127641.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@127641.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@127641.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@127655.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@127655.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@127655.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@127655.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@127655.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@127655.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@127669.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@127669.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@127669.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@127669.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@127669.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@127669.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@127683.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@127683.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@127683.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@127683.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@127683.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@127683.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@127697.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@127697.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@127697.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@127697.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@127697.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@127697.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@127711.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@127711.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@127711.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@127711.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@127711.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@127711.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@127725.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@127725.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@127725.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@127725.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@127725.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@127725.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@127739.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@127739.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@127739.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@127739.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@127739.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@127739.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@127753.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@127753.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@127753.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@127753.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@127753.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@127753.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@127767.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@127767.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@127767.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@127767.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@127767.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@127767.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@127781.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@127781.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@127781.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@127781.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@127781.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@127781.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@127795.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@127795.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@127795.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@127795.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@127795.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@127795.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@127809.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@127809.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@127809.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@127809.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@127809.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@127809.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@127823.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@127823.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@127823.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@127823.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@127823.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@127823.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@127837.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@127837.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@127837.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@127837.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@127837.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@127837.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@127851.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@127851.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@127851.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@127851.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@127851.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@127851.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@127865.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@127865.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@127865.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@127865.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@127865.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@127865.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@127879.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@127879.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@127879.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@127879.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@127879.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@127879.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@127893.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@127893.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@127893.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@127893.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@127893.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@127893.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@127907.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@127907.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@127907.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@127907.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@127907.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@127907.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@127921.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@127921.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@127921.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@127921.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@127921.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@127921.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@127935.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@127935.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@127935.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@127935.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@127935.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@127935.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@127949.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@127949.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@127949.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@127949.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@127949.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@127949.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@127963.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@127963.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@127963.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@127963.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@127963.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@127963.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@127977.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@127977.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@127977.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@127977.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@127977.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@127977.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@127991.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@127991.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@127991.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@127991.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@127991.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@127991.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@128005.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@128005.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@128005.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@128005.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@128005.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@128005.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@128019.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@128019.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@128019.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@128019.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@128019.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@128019.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@128033.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@128033.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@128033.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@128033.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@128033.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@128033.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@128047.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@128047.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@128047.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@128047.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@128047.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@128047.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@128061.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@128061.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@128061.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@128061.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@128061.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@128061.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@128075.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@128075.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@128075.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@128075.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@128075.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@128075.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@128089.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@128089.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@128089.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@128089.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@128089.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@128089.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@128103.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@128103.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@128103.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@128103.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@128103.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@128103.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@128117.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@128117.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@128117.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@128117.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@128117.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@128117.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@128131.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@128131.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@128131.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@128131.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@128131.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@128131.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@128145.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@128145.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@128145.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@128145.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@128145.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@128145.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@128159.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@128159.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@128159.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@128159.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@128159.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@128159.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@128173.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@128173.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@128173.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@128173.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@128173.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@128173.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@128187.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@128187.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@128187.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@128187.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@128187.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@128187.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@128201.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@128201.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@128201.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@128201.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@128201.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@128201.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@128215.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@128215.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@128215.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@128215.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@128215.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@128215.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@128229.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@128229.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@128229.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@128229.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@128229.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@128229.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@128243.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@128243.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@128243.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@128243.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@128243.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@128243.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@128257.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@128257.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@128257.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@128257.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@128257.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@128257.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@128271.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@128271.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@128271.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@128271.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@128271.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@128271.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@128285.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@128285.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@128285.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@128285.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@128285.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@128285.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@128299.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@128299.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@128299.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@128299.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@128299.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@128299.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@128313.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@128313.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@128313.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@128313.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@128313.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@128313.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@128327.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@128327.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@128327.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@128327.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@128327.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@128327.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@128341.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@128341.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@128341.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@128341.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@128341.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@128341.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@128355.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@128355.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@128355.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@128355.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@128355.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@128355.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@128369.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@128369.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@128369.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@128369.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@128369.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@128369.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@128383.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@128383.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@128383.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@128383.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@128383.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@128383.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@128397.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@128397.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@128397.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@128397.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@128397.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@128397.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@128411.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@128411.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@128411.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@128411.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@128411.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@128411.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@128425.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@128425.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@128425.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@128425.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@128425.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@128425.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@128439.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@128439.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@128439.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@128439.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@128439.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@128439.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@128453.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@128453.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@128453.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@128453.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@128453.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@128453.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@128467.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@128467.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@128467.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@128467.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@128467.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@128467.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@128481.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@128481.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@128481.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@128481.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@128481.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@128481.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@128495.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@128495.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@128495.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@128495.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@128495.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@128495.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@128509.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@128509.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@128509.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@128509.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@128509.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@128509.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@128523.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@128523.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@128523.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@128523.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@128523.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@128523.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@128537.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@128537.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@128537.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@128537.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@128537.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@128537.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@128551.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@128551.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@128551.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@128551.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@128551.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@128551.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@128565.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@128565.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@128565.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@128565.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@128565.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@128565.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@128579.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@128579.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@128579.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@128579.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@128579.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@128579.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@128593.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@128593.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@128593.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@128593.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@128593.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@128593.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@128607.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@128607.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@128607.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@128607.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@128607.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@128607.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@128621.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@128621.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@128621.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@128621.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@128621.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@128621.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@128635.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@128635.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@128635.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@128635.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@128635.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@128635.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@128649.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@128649.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@128649.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@128649.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@128649.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@128649.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@128663.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@128663.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@128663.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@128663.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@128663.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@128663.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@128677.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@128677.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@128677.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@128677.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@128677.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@128677.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@128691.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@128691.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@128691.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@128691.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@128691.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@128691.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@128705.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@128705.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@128705.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@128705.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@128705.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@128705.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@128719.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@128719.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@128719.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@128719.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@128719.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@128719.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@128733.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@128733.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@128733.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@128733.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@128733.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@128733.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@128747.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@128747.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@128747.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@128747.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@128747.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@128747.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@128761.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@128761.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@128761.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@128761.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@128761.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@128761.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@128775.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@128775.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@128775.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@128775.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@128775.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@128775.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@128789.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@128789.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@128789.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@128789.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@128789.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@128789.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@128803.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@128803.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@128803.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@128803.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@128803.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@128803.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@128817.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@128817.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@128817.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@128817.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@128817.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@128817.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@128831.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@128831.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@128831.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@128831.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@128831.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@128831.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@128845.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@128845.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@128845.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@128845.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@128845.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@128845.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@128859.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@128859.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@128859.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@128859.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@128859.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@128859.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@128873.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@128873.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@128873.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@128873.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@128873.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@128873.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@128887.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@128887.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@128887.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@128887.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@128887.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@128887.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@128901.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@128901.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@128901.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@128901.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@128901.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@128901.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@128915.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@128915.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@128915.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@128915.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@128915.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@128915.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@128929.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@128929.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@128929.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@128929.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@128929.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@128929.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@128943.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@128943.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@128943.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@128943.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@128943.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@128943.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@128957.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@128957.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@128957.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@128957.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@128957.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@128957.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@128971.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@128971.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@128971.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@128971.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@128971.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@128971.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@128985.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@128985.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@128985.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@128985.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@128985.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@128985.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@128999.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@128999.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@128999.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@128999.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@128999.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@128999.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@129013.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@129013.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@129013.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@129013.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@129013.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@129013.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@129027.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@129027.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@129027.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@129027.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@129027.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@129027.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@129041.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@129041.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@129041.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@129041.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@129041.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@129041.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@129055.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@129055.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@129055.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@129055.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@129055.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@129055.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@129069.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@129069.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@129069.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@129069.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@129069.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@129069.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@129083.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@129083.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@129083.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@129083.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@129083.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@129083.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@129097.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@129097.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@129097.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@129097.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@129097.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@129097.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@129111.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@129111.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@129111.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@129111.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@129111.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@129111.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@129125.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@129125.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@129125.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@129125.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@129125.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@129125.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@129139.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@129139.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@129139.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@129139.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@129139.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@129139.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@129153.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@129153.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@129153.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@129153.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@129153.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@129153.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@129167.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@129167.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@129167.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@129167.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@129167.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@129167.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@129181.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@129181.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@129181.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@129181.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@129181.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@129181.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@129195.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@129195.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@129195.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@129195.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@129195.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@129195.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@129209.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@129209.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@129209.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@129209.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@129209.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@129209.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@129223.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@129223.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@129223.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@129223.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@129223.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@129223.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@129237.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@129237.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@129237.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@129237.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@129237.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@129237.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@129251.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@129251.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@129251.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@129251.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@129251.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@129251.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@129265.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@129265.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@129265.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@129265.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@129265.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@129265.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@129279.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@129279.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@129279.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@129279.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@129279.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@129279.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@129293.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@129293.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@129293.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@129293.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@129293.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@129293.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@129307.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@129307.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@129307.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@129307.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@129307.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@129307.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@129321.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@129321.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@129321.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@129321.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@129321.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@129321.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@129335.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@129335.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@129335.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@129335.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@129335.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@129335.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@129349.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@129349.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@129349.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@129349.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@129349.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@129349.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@129363.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@129363.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@129363.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@129363.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@129363.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@129363.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@129377.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@129377.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@129377.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@129377.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@129377.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@129377.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@129391.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@129391.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@129391.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@129391.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@129391.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@129391.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@129405.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@129405.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@129405.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@129405.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@129405.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@129405.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@129419.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@129419.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@129419.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@129419.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@129419.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@129419.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@129433.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@129433.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@129433.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@129433.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@129433.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@129433.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@129447.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@129447.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@129447.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@129447.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@129447.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@129447.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@129461.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@129461.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@129461.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@129461.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@129461.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@129461.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@129475.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@129475.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@129475.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@129475.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@129475.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@129475.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@129489.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@129489.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@129489.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@129489.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@129489.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@129489.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@129503.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@129503.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@129503.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@129503.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@129503.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@129503.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@129517.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@129517.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@129517.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@129517.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@129517.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@129517.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@129531.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@129531.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@129531.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@129531.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@129531.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@129531.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@129545.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@129545.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@129545.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@129545.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@129545.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@129545.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@129559.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@129559.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@129559.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@129559.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@129559.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@129559.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@129573.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@129573.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@129573.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@129573.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@129573.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@129573.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@129587.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@129587.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@129587.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@129587.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@129587.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@129587.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@129601.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@129601.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@129601.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@129601.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@129601.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@129601.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@129615.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@129615.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@129615.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@129615.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@129615.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@129615.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@129629.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@129629.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@129629.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@129629.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@129629.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@129629.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@129643.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@129643.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@129643.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@129643.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@129643.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@129643.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@129657.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@129657.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@129657.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@129657.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@129657.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@129657.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@129671.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@129671.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@129671.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@129671.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@129671.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@129671.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@129685.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@129685.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@129685.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@129685.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@129685.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@129685.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@129699.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@129699.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@129699.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@129699.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@129699.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@129699.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@129713.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@129713.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@129713.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@129713.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@129713.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@129713.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@129727.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@129727.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@129727.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@129727.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@129727.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@129727.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@129741.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@129741.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@129741.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@129741.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@129741.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@129741.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@129755.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@129755.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@129755.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@129755.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@129755.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@129755.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@129769.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@129769.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@129769.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@129769.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@129769.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@129769.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@129783.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@129783.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@129783.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@129783.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@129783.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@129783.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@129797.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@129797.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@129797.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@129797.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@129797.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@129797.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@129811.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@129811.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@129811.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@129811.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@129811.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@129811.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@129825.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@129825.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@129825.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@129825.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@129825.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@129825.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@129839.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@129839.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@129839.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@129839.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@129839.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@129839.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@129853.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@129853.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@129853.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@129853.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@129853.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@129853.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@129867.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@129867.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@129867.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@129867.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@129867.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@129867.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@129881.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@129881.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@129881.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@129881.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@129881.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@129881.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@129895.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@129895.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@129895.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@129895.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@129895.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@129895.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@129909.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@129909.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@129909.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@129909.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@129909.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@129909.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@129923.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@129923.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@129923.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@129923.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@129923.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@129923.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@129937.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@129937.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@129937.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@129937.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@129937.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@129937.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@129951.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@129951.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@129951.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@129951.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@129951.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@129951.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@129965.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@129965.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@129965.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@129965.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@129965.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@129965.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@129979.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@129979.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@129979.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@129979.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@129979.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@129979.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@129993.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@129993.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@129993.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@129993.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@129993.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@129993.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@130007.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@130007.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@130007.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@130007.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@130007.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@130007.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@130021.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@130021.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@130021.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@130021.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@130021.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@130021.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@130035.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@130035.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@130035.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@130035.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@130035.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@130035.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@130049.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@130049.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@130049.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@130049.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@130049.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@130049.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@130063.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@130063.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@130063.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@130063.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@130063.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@130063.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@130077.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@130077.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@130077.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@130077.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@130077.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@130077.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@130091.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@130091.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@130091.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@130091.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@130091.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@130091.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@130105.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@130105.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@130105.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@130105.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@130105.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@130105.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@130119.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@130119.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@130119.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@130119.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@130119.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@130119.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@130133.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@130133.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@130133.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@130133.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@130133.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@130133.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@130147.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@130147.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@130147.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@130147.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@130147.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@130147.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@130161.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@130161.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@130161.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@130161.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@130161.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@130161.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@130175.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@130175.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@130175.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@130175.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@130175.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@130175.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@130189.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@130189.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@130189.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@130189.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@130189.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@130189.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@130203.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@130203.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@130203.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@130203.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@130203.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@130203.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@130217.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@130217.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@130217.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@130217.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@130217.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@130217.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@130231.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@130231.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@130231.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@130231.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@130231.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@130231.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@130245.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@130245.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@130245.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@130245.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@130245.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@130245.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@130259.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@130259.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@130259.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@130259.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@130259.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@130259.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@130273.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@130273.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@130273.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@130273.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@130273.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@130273.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@130287.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@130287.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@130287.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@130287.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@130287.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@130287.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@130301.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@130301.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@130301.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@130301.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@130301.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@130301.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@130315.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@130315.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@130315.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@130315.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@130315.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@130315.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@130329.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@130329.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@130329.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@130329.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@130329.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@130329.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@130343.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@130343.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@130343.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@130343.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@130343.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@130343.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@130357.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@130357.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@130357.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@130357.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@130357.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@130357.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@130371.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@130371.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@130371.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@130371.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@130371.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@130371.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@130385.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@130385.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@130385.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@130385.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@130385.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@130385.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@130399.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@130399.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@130399.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@130399.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@130399.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@130399.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@130413.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@130413.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@130413.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@130413.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@130413.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@130413.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@130427.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@130427.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@130427.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@130427.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@130427.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@130427.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@130441.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@130441.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@130441.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@130441.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@130441.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@130441.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@130455.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@130455.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@130455.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@130455.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@130455.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@130455.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@130469.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@130469.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@130469.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@130469.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@130469.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@130469.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@130483.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@130483.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@130483.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@130483.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@130483.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@130483.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@130497.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@130497.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@130497.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@130497.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@130497.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@130497.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@130511.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@130511.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@130511.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@130511.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@130511.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@130511.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@130525.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@130525.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@130525.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@130525.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@130525.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@130525.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@130539.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@130539.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@130539.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@130539.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@130539.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@130539.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@130553.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@130553.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@130553.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@130553.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@130553.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@130553.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@130567.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@130567.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@130567.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@130567.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@130567.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@130567.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@130581.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@130581.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@130581.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@130581.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@130581.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@130581.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@130595.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@130595.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@130595.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@130595.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@130595.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@130595.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@130609.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@130609.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@130609.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@130609.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@130609.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@130609.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@130623.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@130623.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@130623.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@130623.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@130623.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@130623.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@130637.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@130637.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@130637.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@130637.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@130637.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@130637.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@130651.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@130651.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@130651.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@130651.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@130651.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@130651.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@130665.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@130665.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@130665.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@130665.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@130665.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@130665.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@130679.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@130679.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@130679.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@130679.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@130679.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@130679.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@130693.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@130693.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@130693.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@130693.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@130693.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@130693.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@130707.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@130707.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@130707.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@130707.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@130707.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@130707.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@130721.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@130721.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@130721.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@130721.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@130721.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@130721.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@130735.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@130735.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@130735.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@130735.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@130735.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@130735.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@130749.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@130749.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@130749.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@130749.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@130749.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@130749.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@130763.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@130763.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@130763.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@130763.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@130763.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@130763.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@130777.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@130777.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@130777.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@130777.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@130777.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@130777.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@130791.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@130791.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@130791.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@130791.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@130791.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@130791.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@130805.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@130805.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@130805.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@130805.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@130805.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@130805.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@130819.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@130819.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@130819.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@130819.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@130819.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@130819.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@130833.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@130833.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@130833.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@130833.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@130833.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@130833.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@130847.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@130847.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@130847.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@130847.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@130847.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@130847.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@130861.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@130861.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@130861.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@130861.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@130861.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@130861.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@130875.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@130875.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@130875.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@130875.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@130875.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@130875.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@130889.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@130889.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@130889.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@130889.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@130889.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@130889.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@130903.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@130903.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@130903.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@130903.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@130903.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@130903.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@130917.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@130917.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@130917.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@130917.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@130917.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@130917.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@130931.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@130931.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@130931.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@130931.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@130931.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@130931.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@130945.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@130945.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@130945.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@130945.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@130945.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@130945.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@130959.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@130959.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@130959.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@130959.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@130959.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@130959.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@130973.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@130973.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@130973.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@130973.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@130973.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@130973.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@130987.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@130987.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@130987.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@130987.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@130987.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@130987.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@131001.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@131001.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@131001.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@131001.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@131001.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@131001.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@131015.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@131015.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@131015.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@131015.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@131015.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@131015.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@131029.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@131029.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@131029.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@131029.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@131029.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@131029.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@131043.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@131043.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@131043.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@131043.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@131043.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@131043.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@131057.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@131057.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@131057.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@131057.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@131057.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@131057.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@131071.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@131071.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@131071.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@131071.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@131071.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@131071.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@131085.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@131085.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@131085.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@131085.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@131085.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@131085.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@131099.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@131099.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@131099.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@131099.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@131099.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@131099.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@131113.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@131113.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@131113.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@131113.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@131113.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@131113.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@131127.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@131127.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@131127.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@131127.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@131127.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@131127.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@131141.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@131141.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@131141.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@131141.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@131141.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@131141.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@131155.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@131155.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@131155.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@131155.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@131155.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@131155.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@131169.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@131169.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@131169.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@131169.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@131169.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@131169.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@131183.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@131183.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@131183.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@131183.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@131183.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@131183.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@131197.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@131197.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@131197.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@131197.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@131197.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@131197.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@131211.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@131211.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@131211.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@131211.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@131211.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@131211.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@131225.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@131225.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@131225.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@131225.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@131225.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@131225.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@131239.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@131239.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@131239.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@131239.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@131239.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@131239.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@131253.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@131253.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@131253.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@131253.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@131253.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@131253.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@131267.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@131267.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@131267.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@131267.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@131267.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@131267.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@131281.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@131281.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@131281.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@131281.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@131281.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@131281.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@131295.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@131295.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@131295.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@131295.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@131295.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@131295.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@131309.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@131309.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@131309.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@131309.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@131309.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@131309.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@131323.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@131323.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@131323.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@131323.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@131323.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@131323.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@131337.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@131337.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@131337.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@131337.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@131337.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@131337.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@131351.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@131351.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@131351.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@131351.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@131351.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@131351.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@131365.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@131365.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@131365.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@131365.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@131365.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@131365.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@131379.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@131379.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@131379.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@131379.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@131379.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@131379.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@131393.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@131393.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@131393.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@131393.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@131393.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@131393.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@131407.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@131407.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@131407.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@131407.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@131407.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@131407.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@131421.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@131421.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@131421.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@131421.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@131421.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@131421.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@131435.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@131435.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@131435.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@131435.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@131435.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@131435.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@131449.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@131449.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@131449.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@131449.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@131449.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@131449.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@131463.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@131463.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@131463.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@131463.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@131463.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@131463.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@131477.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@131477.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@131477.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@131477.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@131477.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@131477.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@131491.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@131491.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@131491.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@131491.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@131491.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@131491.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@131505.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@131505.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@131505.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@131505.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@131505.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@131505.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@131519.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@131519.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@131519.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@131519.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@131519.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@131519.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@131533.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@131533.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@131533.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@131533.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@131533.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@131533.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@131547.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@131547.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@131547.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@131547.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@131547.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@131547.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@131561.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@131561.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@131561.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@131561.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@131561.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@131561.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@131575.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@131575.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@131575.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@131575.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@131575.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@131575.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@131589.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@131589.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@131589.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@131589.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@131589.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@131589.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@131603.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@131603.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@131603.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@131603.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@131603.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@131603.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@131617.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@131617.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@131617.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@131617.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@131617.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@131617.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@131631.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@131631.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@131631.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@131631.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@131631.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@131631.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@131645.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@131645.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@131645.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@131645.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@131645.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@131645.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@131659.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@131659.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@131659.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@131659.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@131659.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@131659.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@131673.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@131673.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@131673.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@131673.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@131673.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@131673.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@131687.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@131687.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@131687.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@131687.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@131687.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@131687.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@131701.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@131701.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@131701.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@131701.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@131701.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@131701.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@131715.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@131715.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@131715.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@131715.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@131715.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@131715.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@131729.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@131729.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@131729.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@131729.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@131729.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@131729.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@131743.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@131743.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@131743.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@131743.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@131743.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@131743.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@131757.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@131757.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@131757.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@131757.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@131757.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@131757.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@131771.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@131771.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@131771.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@131771.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@131771.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@131771.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@131785.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@131785.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@131785.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@131785.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@131785.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@131785.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@131799.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@131799.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@131799.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@131799.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@131799.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@131799.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@131813.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@131813.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@131813.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@131813.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@131813.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@131813.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@131827.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@131827.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@131827.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@131827.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@131827.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@131827.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@131841.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@131841.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@131841.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@131841.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@131841.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@131841.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@131855.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@131855.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@131855.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@131855.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@131855.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@131855.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@131869.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@131869.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@131869.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@131869.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@131869.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@131869.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@131883.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@131883.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@131883.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@131883.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@131883.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@131883.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@131897.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@131897.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@131897.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@131897.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@131897.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@131897.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@131911.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@131911.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@131911.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@131911.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@131911.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@131911.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@131925.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@131925.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@131925.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@131925.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@131925.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@131925.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@131939.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@131939.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@131939.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@131939.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@131939.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@131939.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@131953.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@131953.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@131953.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@131953.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@131953.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@131953.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@131967.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@131967.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@131967.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@131967.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@131967.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@131967.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@131981.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@131981.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@131981.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@131981.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@131981.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@131981.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@131995.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@131995.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@131995.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@131995.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@131995.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@131995.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@132009.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@132009.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@132009.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@132009.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@132009.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@132009.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@132023.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@132023.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@132023.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@132023.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@132023.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@132023.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@132037.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@132037.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@132037.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@132037.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@132037.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@132037.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@132051.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@132051.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@132051.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@132051.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@132051.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@132051.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@132065.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@132065.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@132065.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@132065.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@132065.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@132065.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@132079.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@132079.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@132079.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@132079.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@132079.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@132079.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@132093.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@132093.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@132093.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@132093.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@132093.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@132093.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@132107.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@132107.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@132107.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@132107.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@132107.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@132107.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@132121.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@132121.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@132121.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@132121.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@132121.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@132121.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@132135.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@132135.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@132135.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@132135.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@132135.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@132135.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@132149.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@132149.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@132149.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@132149.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@132149.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@132149.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@132163.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@132163.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@132163.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@132163.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@132163.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@132163.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@132177.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@132177.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@132177.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@132177.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@132177.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@132177.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@132191.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@132191.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@132191.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@132191.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@132191.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@132191.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@132205.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@132205.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@132205.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@132205.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@132205.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@132205.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@132219.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@132219.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@132219.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@132219.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@132219.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@132219.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@132233.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@132233.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@132233.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@132233.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@132233.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@132233.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@132247.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@132247.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@132247.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@132247.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@132247.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@132247.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@132261.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@132261.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@132261.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@132261.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@132261.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@132261.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@132275.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@132275.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@132275.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@132275.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@132275.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@132275.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@132289.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@132289.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@132289.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@132289.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@132289.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@132289.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@132303.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@132303.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@132303.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@132303.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@132303.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@132303.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@132317.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@132317.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@132317.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@132317.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@132317.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@132317.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@132331.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@132331.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@132331.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@132331.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@132331.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@132331.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@132345.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@132345.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@132345.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@132345.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@132345.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@132345.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@132359.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@132359.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@132359.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@132359.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@132359.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@132359.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@132373.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@132373.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@132373.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@132373.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@132373.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@132373.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@132387.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@132387.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@132387.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@132387.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@132387.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@132387.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@132401.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@132401.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@132401.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@132401.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@132401.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@132401.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@132415.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@132415.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@132415.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@132415.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@132415.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@132415.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@132429.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@132429.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@132429.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@132429.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@132429.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@132429.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@132443.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@132443.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@132443.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@132443.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@132443.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@132443.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@132457.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@132457.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@132457.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@132457.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@132457.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@132457.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@132471.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@132471.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@132471.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@132471.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@132471.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@132471.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@132485.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@132485.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@132485.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@132485.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@132485.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@132485.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@132499.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@132499.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@132499.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@132499.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@132499.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@132499.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@132513.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@132513.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@132513.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@132513.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@132513.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@132513.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@132527.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@132527.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@132527.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@132527.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@132527.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@132527.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@132541.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@132541.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@132541.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@132541.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@132541.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@132541.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@132555.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@132555.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@132555.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@132555.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@132555.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@132555.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@132569.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@132569.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@132569.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@132569.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@132569.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@132569.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@132583.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@132583.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@132583.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@132583.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@132583.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@132583.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@132597.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@132597.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@132597.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@132597.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@132597.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@132597.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@132611.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@132611.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@132611.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@132611.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@132611.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@132611.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@132625.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@132625.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@132625.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@132625.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@132625.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@132625.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@132639.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@132639.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@132639.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@132639.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@132639.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@132639.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@132653.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@132653.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@132653.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@132653.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@132653.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@132653.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@132667.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@132667.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@132667.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@132667.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@132667.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@132667.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@132681.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@132681.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@132681.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@132681.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@132681.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@132681.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@132695.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@132695.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@132695.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@132695.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@132695.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@132695.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@132709.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@132709.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@132709.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@132709.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@132709.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@132709.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@132723.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@132723.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@132723.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@132723.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@132723.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@132723.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@132737.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@132737.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@132737.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@132737.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@132737.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@132737.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@132751.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@132751.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@132751.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@132751.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@132751.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@132751.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@132765.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@132765.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@132765.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@132765.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@132765.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@132765.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@132779.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@132779.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@132779.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@132779.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@132779.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@132779.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@132793.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@132793.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@132793.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@132793.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@132793.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@132793.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@132807.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@132807.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@132807.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@132807.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@132807.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@132807.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@132821.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@132821.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@132821.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@132821.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@132821.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@132821.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@132835.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@132835.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@132835.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@132835.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@132835.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@132835.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@132849.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@132849.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@132849.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@132849.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@132849.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@132849.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@132863.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@132863.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@132863.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@132863.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@132863.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@132863.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@132877.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@132877.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@132877.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@132877.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@132877.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@132877.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@132891.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@132891.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@132891.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@132891.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@132891.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@132891.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@132905.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@132905.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@132905.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@132905.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@132905.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@132905.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@132919.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@132919.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@132919.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@132919.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@132919.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@132919.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@132933.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@132933.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@132933.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@132933.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@132933.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@132933.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@132947.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@132947.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@132947.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@132947.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@132947.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@132947.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@132961.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@132961.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@132961.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@132961.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@132961.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@132961.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@132975.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@132975.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@132975.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@132975.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@132975.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@132975.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@132989.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@132989.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@132989.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@132989.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@132989.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@132989.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@133003.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@133003.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@133003.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@133003.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@133003.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@133003.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@133017.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@133017.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@133017.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@133017.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@133017.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@133017.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@133031.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@133031.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@133031.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@133031.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@133031.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@133031.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@133045.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@133045.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@133045.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@133045.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@133045.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@133045.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@133059.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@133059.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@133059.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@133059.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@133059.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@133059.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@133073.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@133073.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@133073.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@133073.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@133073.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@133073.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@133087.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@133087.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@133087.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@133087.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@133087.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@133087.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@133101.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@133101.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@133101.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@133101.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@133101.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@133101.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@133115.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@133115.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@133115.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@133115.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@133115.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@133115.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@133129.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@133129.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@133129.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@133129.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@133129.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@133129.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@133143.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@133143.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@133143.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@133143.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@133143.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@133143.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@133157.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@133157.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@133157.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@133157.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@133157.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@133157.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@133171.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@133171.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@133171.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@133171.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@133171.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@133171.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@133185.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@133185.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@133185.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@133185.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@133185.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@133185.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@133199.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@133199.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@133199.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@133199.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@133199.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@133199.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@133213.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@133213.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@133213.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@133213.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@133213.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@133213.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@133227.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@133227.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@133227.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@133227.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@133227.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@133227.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@133241.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@133241.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@133241.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@133241.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@133241.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@133241.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@133255.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@133255.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@133255.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@133255.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@133255.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@133255.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@133269.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@133269.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@133269.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@133269.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@133269.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@133269.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@133283.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@133283.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@133283.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@133283.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@133283.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@133283.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@133297.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@133297.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@133297.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@133297.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@133297.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@133297.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@133311.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@133311.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@133311.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@133311.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@133311.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@133311.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@133325.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@133325.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@133325.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@133325.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@133325.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@133325.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@133339.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@133339.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@133339.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@133339.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@133339.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@133339.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@133353.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@133353.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@133353.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@133353.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@133353.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@133353.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@133367.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@133367.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@133367.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@133367.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@133367.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@133367.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@133381.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@133381.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@133381.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@133381.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@133381.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@133381.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@133395.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@133395.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@133395.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@133395.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@133395.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@133395.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@133409.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@133409.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@133409.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@133409.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@133409.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@133409.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@133423.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@133423.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@133423.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@133423.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@133423.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@133423.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@133437.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@133437.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@133437.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@133437.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@133437.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@133437.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@133451.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@133451.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@133451.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@133451.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@133451.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@133451.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@133465.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@133465.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@133465.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@133465.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@133465.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@133465.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@133479.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@133479.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@133479.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@133479.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@133479.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@133479.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@133493.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@133493.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@133493.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@133493.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@133493.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@133493.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@133507.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@133507.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@133507.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@133507.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@133507.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@133507.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@133521.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@133521.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@133521.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@133521.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@133521.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@133521.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@133535.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@133535.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@133535.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@133535.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@133535.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@133535.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@133549.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@133549.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@133549.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@133549.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@133549.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@133549.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@133563.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@133563.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@133563.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@133563.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@133563.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@133563.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@133577.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@133577.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@133577.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@133577.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@133577.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@133577.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@133591.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@133591.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@133591.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@133591.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@133591.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@133591.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@133605.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@133605.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@133605.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@133605.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@133605.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@133605.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@133619.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@133619.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@133619.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@133619.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@133619.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@133619.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@133633.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@133633.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@133633.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@133633.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@133633.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@133633.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@133647.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@133647.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@133647.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@133647.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@133647.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@133647.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@133661.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@133661.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@133661.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@133661.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@133661.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@133661.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@133675.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@133675.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@133675.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@133675.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@133675.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@133675.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@133689.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@133689.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@133689.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@133689.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@133689.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@133689.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@133703.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@133703.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@133703.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@133703.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@133703.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@133703.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@133717.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@133717.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@133717.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@133717.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@133717.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@133717.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@133731.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@133731.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@133731.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@133731.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@133731.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@133731.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@133745.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@133745.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@133745.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@133745.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@133745.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@133745.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@133759.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@133759.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@133759.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@133759.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@133759.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@133759.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@133773.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@133773.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@133773.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@133773.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@133773.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@133773.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@133787.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@133787.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@133787.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@133787.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@133787.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@133787.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@133801.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@133801.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@133801.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@133801.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@133801.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@133801.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@133815.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@133815.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@133815.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@133815.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@133815.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@133815.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@133829.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@133829.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@133829.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@133829.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@133829.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@133829.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@133843.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@133843.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@133843.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@133843.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@133843.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@133843.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@133857.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@133857.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@133857.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@133857.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@133857.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@133857.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@133871.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@133871.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@133871.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@133871.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@133871.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@133871.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@133885.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@133885.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@133885.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@133885.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@133885.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@133885.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@133899.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@133899.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@133899.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@133899.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@133899.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@133899.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@133913.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@133913.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@133913.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@133913.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@133913.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@133913.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@133927.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@133927.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@133927.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@133927.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@133927.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@133927.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@133941.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@133941.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@133941.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@133941.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@133941.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@133941.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@133955.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@133955.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@133955.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@133955.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@133955.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@133955.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@133969.4]
  wire [8:0] rport_io_sel; // @[RegFile.scala 95:21:@133969.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@133969.4]
  wire  _T_3078; // @[RegFile.scala 80:42:@126931.4]
  wire  _T_3084; // @[RegFile.scala 68:46:@126943.4]
  wire  _T_3085; // @[RegFile.scala 68:34:@126944.4]
  wire  _T_3098; // @[RegFile.scala 80:42:@126962.4]
  wire  _T_3104; // @[RegFile.scala 80:42:@126974.4]
  wire  _T_3110; // @[RegFile.scala 74:80:@126986.4]
  wire  _T_3111; // @[RegFile.scala 74:68:@126987.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@126928.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@126940.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@126959.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@126971.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@126983.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@126997.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@127011.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@127025.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@127039.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@127053.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@127067.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@127081.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@127095.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@127109.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@127123.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@127137.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@127151.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@127165.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@127179.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@127193.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@127207.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@127221.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@127235.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@127249.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@127263.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@127277.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@127291.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@127305.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@127319.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@127333.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@127347.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@127361.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@127375.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@127389.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@127403.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@127417.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@127431.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@127445.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@127459.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@127473.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@127487.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@127501.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@127515.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@127529.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@127543.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@127557.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@127571.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@127585.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@127599.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@127613.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@127627.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@127641.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@127655.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@127669.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@127683.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@127697.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@127711.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@127725.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@127739.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@127753.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@127767.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@127781.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@127795.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@127809.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@127823.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@127837.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@127851.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@127865.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@127879.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@127893.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@127907.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@127921.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@127935.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@127949.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@127963.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@127977.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@127991.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@128005.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@128019.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@128033.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@128047.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@128061.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@128075.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@128089.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@128103.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@128117.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@128131.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@128145.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@128159.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@128173.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@128187.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@128201.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@128215.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@128229.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@128243.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@128257.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@128271.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@128285.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@128299.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@128313.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@128327.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@128341.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@128355.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@128369.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@128383.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@128397.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@128411.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@128425.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@128439.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@128453.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@128467.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@128481.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@128495.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@128509.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@128523.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@128537.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@128551.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@128565.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@128579.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@128593.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@128607.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@128621.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@128635.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@128649.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@128663.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@128677.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@128691.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@128705.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@128719.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@128733.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@128747.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@128761.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@128775.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@128789.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@128803.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@128817.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@128831.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@128845.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@128859.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@128873.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@128887.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@128901.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@128915.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@128929.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@128943.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@128957.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@128971.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@128985.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@128999.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@129013.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@129027.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@129041.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@129055.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@129069.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@129083.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@129097.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@129111.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@129125.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@129139.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@129153.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@129167.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@129181.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@129195.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@129209.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@129223.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@129237.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@129251.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@129265.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@129279.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@129293.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@129307.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@129321.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@129335.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@129349.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@129363.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@129377.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@129391.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@129405.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@129419.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@129433.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@129447.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@129461.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@129475.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@129489.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@129503.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@129517.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@129531.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@129545.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@129559.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@129573.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@129587.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@129601.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@129615.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@129629.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@129643.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@129657.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@129671.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@129685.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@129699.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@129713.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@129727.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@129741.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@129755.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@129769.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@129783.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@129797.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@129811.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@129825.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@129839.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@129853.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@129867.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@129881.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@129895.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@129909.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@129923.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@129937.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@129951.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@129965.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@129979.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@129993.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@130007.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@130021.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@130035.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@130049.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@130063.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@130077.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@130091.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@130105.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@130119.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@130133.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@130147.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@130161.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@130175.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@130189.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@130203.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@130217.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@130231.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@130245.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@130259.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@130273.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@130287.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@130301.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@130315.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@130329.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@130343.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@130357.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@130371.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@130385.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@130399.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@130413.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@130427.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@130441.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@130455.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@130469.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@130483.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@130497.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@130511.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@130525.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@130539.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@130553.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@130567.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@130581.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@130595.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@130609.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@130623.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@130637.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@130651.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@130665.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@130679.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@130693.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@130707.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@130721.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@130735.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@130749.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@130763.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@130777.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@130791.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@130805.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@130819.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@130833.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@130847.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@130861.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@130875.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@130889.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@130903.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@130917.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@130931.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@130945.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@130959.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@130973.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@130987.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@131001.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@131015.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@131029.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@131043.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@131057.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@131071.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@131085.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@131099.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@131113.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@131127.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@131141.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@131155.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@131169.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@131183.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@131197.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@131211.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@131225.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@131239.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@131253.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@131267.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@131281.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@131295.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@131309.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@131323.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@131337.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@131351.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@131365.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@131379.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@131393.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@131407.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@131421.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@131435.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@131449.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@131463.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@131477.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@131491.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@131505.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@131519.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@131533.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@131547.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@131561.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@131575.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@131589.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@131603.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@131617.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@131631.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@131645.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@131659.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@131673.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@131687.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@131701.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@131715.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@131729.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@131743.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@131757.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@131771.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@131785.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@131799.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@131813.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@131827.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@131841.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@131855.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@131869.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@131883.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@131897.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@131911.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@131925.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@131939.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@131953.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@131967.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@131981.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@131995.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@132009.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@132023.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@132037.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@132051.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@132065.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@132079.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@132093.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@132107.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@132121.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@132135.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@132149.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@132163.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@132177.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@132191.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@132205.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@132219.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@132233.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@132247.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@132261.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@132275.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@132289.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@132303.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@132317.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@132331.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@132345.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@132359.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@132373.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@132387.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@132401.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@132415.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@132429.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@132443.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@132457.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@132471.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@132485.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@132499.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@132513.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@132527.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@132541.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@132555.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@132569.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@132583.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@132597.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@132611.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@132625.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@132639.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@132653.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@132667.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@132681.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@132695.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@132709.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@132723.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@132737.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@132751.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@132765.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@132779.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@132793.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@132807.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@132821.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@132835.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@132849.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@132863.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@132877.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@132891.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@132905.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@132919.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@132933.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@132947.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@132961.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@132975.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@132989.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@133003.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@133017.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@133031.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@133045.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@133059.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@133073.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@133087.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@133101.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@133115.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@133129.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@133143.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@133157.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@133171.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@133185.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@133199.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@133213.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@133227.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@133241.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@133255.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@133269.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@133283.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@133297.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@133311.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@133325.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@133339.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@133353.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@133367.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@133381.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@133395.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@133409.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@133423.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@133437.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@133451.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@133465.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@133479.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@133493.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@133507.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@133521.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@133535.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@133549.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@133563.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@133577.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@133591.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@133605.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@133619.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@133633.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@133647.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@133661.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@133675.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@133689.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@133703.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@133717.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@133731.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@133745.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@133759.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@133773.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@133787.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@133801.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@133815.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@133829.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@133843.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@133857.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@133871.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@133885.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@133899.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@133913.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@133927.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@133941.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@133955.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  MuxN rport ( // @[RegFile.scala 95:21:@133969.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3078 = io_waddr == 32'h0; // @[RegFile.scala 80:42:@126931.4]
  assign _T_3084 = io_waddr == 32'h1; // @[RegFile.scala 68:46:@126943.4]
  assign _T_3085 = io_wen & _T_3084; // @[RegFile.scala 68:34:@126944.4]
  assign _T_3098 = io_waddr == 32'h2; // @[RegFile.scala 80:42:@126962.4]
  assign _T_3104 = io_waddr == 32'h3; // @[RegFile.scala 80:42:@126974.4]
  assign _T_3110 = io_waddr == 32'h4; // @[RegFile.scala 74:80:@126986.4]
  assign _T_3111 = io_wen & _T_3110; // @[RegFile.scala 74:68:@126987.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@134980.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@134986.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@134987.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@134988.4]
  assign io_argIns_3 = regs_3_io_out; // @[RegFile.scala 111:13:@134989.4]
  assign regs_0_clock = clock; // @[:@126929.4]
  assign regs_0_reset = reset; // @[:@126930.4 RegFile.scala 82:16:@126936.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@126934.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@126938.4]
  assign regs_0_io_enable = io_wen & _T_3078; // @[RegFile.scala 80:20:@126933.4]
  assign regs_1_clock = clock; // @[:@126941.4]
  assign regs_1_reset = reset; // @[:@126942.4 RegFile.scala 70:16:@126954.4]
  assign regs_1_io_in = _T_3085 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@126952.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@126957.4]
  assign regs_1_io_enable = _T_3085 ? _T_3085 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@126948.4]
  assign regs_2_clock = clock; // @[:@126960.4]
  assign regs_2_reset = reset; // @[:@126961.4 RegFile.scala 82:16:@126967.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@126965.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@126969.4]
  assign regs_2_io_enable = io_wen & _T_3098; // @[RegFile.scala 80:20:@126964.4]
  assign regs_3_clock = clock; // @[:@126972.4]
  assign regs_3_reset = reset; // @[:@126973.4 RegFile.scala 82:16:@126979.4]
  assign regs_3_io_in = io_wdata; // @[RegFile.scala 81:16:@126977.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 83:19:@126981.4]
  assign regs_3_io_enable = io_wen & _T_3104; // @[RegFile.scala 80:20:@126976.4]
  assign regs_4_clock = clock; // @[:@126984.4]
  assign regs_4_reset = io_reset; // @[:@126985.4 RegFile.scala 76:16:@126992.4]
  assign regs_4_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@126991.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@126995.4]
  assign regs_4_io_enable = io_argOuts_1_valid | _T_3111; // @[RegFile.scala 74:20:@126989.4]
  assign regs_5_clock = clock; // @[:@126998.4]
  assign regs_5_reset = io_reset; // @[:@126999.4 RegFile.scala 76:16:@127006.4]
  assign regs_5_io_in = 64'h0; // @[RegFile.scala 75:16:@127005.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@127009.4]
  assign regs_5_io_enable = 1'h1; // @[RegFile.scala 74:20:@127003.4]
  assign regs_6_clock = clock; // @[:@127012.4]
  assign regs_6_reset = io_reset; // @[:@127013.4 RegFile.scala 76:16:@127020.4]
  assign regs_6_io_in = 64'h0; // @[RegFile.scala 75:16:@127019.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@127023.4]
  assign regs_6_io_enable = 1'h1; // @[RegFile.scala 74:20:@127017.4]
  assign regs_7_clock = clock; // @[:@127026.4]
  assign regs_7_reset = io_reset; // @[:@127027.4 RegFile.scala 76:16:@127034.4]
  assign regs_7_io_in = 64'h0; // @[RegFile.scala 75:16:@127033.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@127037.4]
  assign regs_7_io_enable = 1'h1; // @[RegFile.scala 74:20:@127031.4]
  assign regs_8_clock = clock; // @[:@127040.4]
  assign regs_8_reset = io_reset; // @[:@127041.4 RegFile.scala 76:16:@127048.4]
  assign regs_8_io_in = 64'h0; // @[RegFile.scala 75:16:@127047.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@127051.4]
  assign regs_8_io_enable = 1'h1; // @[RegFile.scala 74:20:@127045.4]
  assign regs_9_clock = clock; // @[:@127054.4]
  assign regs_9_reset = io_reset; // @[:@127055.4 RegFile.scala 76:16:@127062.4]
  assign regs_9_io_in = 64'h0; // @[RegFile.scala 75:16:@127061.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@127065.4]
  assign regs_9_io_enable = 1'h1; // @[RegFile.scala 74:20:@127059.4]
  assign regs_10_clock = clock; // @[:@127068.4]
  assign regs_10_reset = io_reset; // @[:@127069.4 RegFile.scala 76:16:@127076.4]
  assign regs_10_io_in = 64'h0; // @[RegFile.scala 75:16:@127075.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@127079.4]
  assign regs_10_io_enable = 1'h1; // @[RegFile.scala 74:20:@127073.4]
  assign regs_11_clock = clock; // @[:@127082.4]
  assign regs_11_reset = io_reset; // @[:@127083.4 RegFile.scala 76:16:@127090.4]
  assign regs_11_io_in = 64'h0; // @[RegFile.scala 75:16:@127089.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@127093.4]
  assign regs_11_io_enable = 1'h1; // @[RegFile.scala 74:20:@127087.4]
  assign regs_12_clock = clock; // @[:@127096.4]
  assign regs_12_reset = io_reset; // @[:@127097.4 RegFile.scala 76:16:@127104.4]
  assign regs_12_io_in = 64'h0; // @[RegFile.scala 75:16:@127103.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@127107.4]
  assign regs_12_io_enable = 1'h1; // @[RegFile.scala 74:20:@127101.4]
  assign regs_13_clock = clock; // @[:@127110.4]
  assign regs_13_reset = io_reset; // @[:@127111.4 RegFile.scala 76:16:@127118.4]
  assign regs_13_io_in = 64'h0; // @[RegFile.scala 75:16:@127117.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@127121.4]
  assign regs_13_io_enable = 1'h1; // @[RegFile.scala 74:20:@127115.4]
  assign regs_14_clock = clock; // @[:@127124.4]
  assign regs_14_reset = io_reset; // @[:@127125.4 RegFile.scala 76:16:@127132.4]
  assign regs_14_io_in = 64'h0; // @[RegFile.scala 75:16:@127131.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@127135.4]
  assign regs_14_io_enable = 1'h1; // @[RegFile.scala 74:20:@127129.4]
  assign regs_15_clock = clock; // @[:@127138.4]
  assign regs_15_reset = io_reset; // @[:@127139.4 RegFile.scala 76:16:@127146.4]
  assign regs_15_io_in = 64'h0; // @[RegFile.scala 75:16:@127145.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@127149.4]
  assign regs_15_io_enable = 1'h1; // @[RegFile.scala 74:20:@127143.4]
  assign regs_16_clock = clock; // @[:@127152.4]
  assign regs_16_reset = io_reset; // @[:@127153.4 RegFile.scala 76:16:@127160.4]
  assign regs_16_io_in = 64'h0; // @[RegFile.scala 75:16:@127159.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@127163.4]
  assign regs_16_io_enable = 1'h1; // @[RegFile.scala 74:20:@127157.4]
  assign regs_17_clock = clock; // @[:@127166.4]
  assign regs_17_reset = io_reset; // @[:@127167.4 RegFile.scala 76:16:@127174.4]
  assign regs_17_io_in = 64'h0; // @[RegFile.scala 75:16:@127173.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@127177.4]
  assign regs_17_io_enable = 1'h1; // @[RegFile.scala 74:20:@127171.4]
  assign regs_18_clock = clock; // @[:@127180.4]
  assign regs_18_reset = io_reset; // @[:@127181.4 RegFile.scala 76:16:@127188.4]
  assign regs_18_io_in = 64'h0; // @[RegFile.scala 75:16:@127187.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@127191.4]
  assign regs_18_io_enable = 1'h1; // @[RegFile.scala 74:20:@127185.4]
  assign regs_19_clock = clock; // @[:@127194.4]
  assign regs_19_reset = io_reset; // @[:@127195.4 RegFile.scala 76:16:@127202.4]
  assign regs_19_io_in = 64'h0; // @[RegFile.scala 75:16:@127201.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@127205.4]
  assign regs_19_io_enable = 1'h1; // @[RegFile.scala 74:20:@127199.4]
  assign regs_20_clock = clock; // @[:@127208.4]
  assign regs_20_reset = io_reset; // @[:@127209.4 RegFile.scala 76:16:@127216.4]
  assign regs_20_io_in = 64'h0; // @[RegFile.scala 75:16:@127215.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@127219.4]
  assign regs_20_io_enable = 1'h1; // @[RegFile.scala 74:20:@127213.4]
  assign regs_21_clock = clock; // @[:@127222.4]
  assign regs_21_reset = io_reset; // @[:@127223.4 RegFile.scala 76:16:@127230.4]
  assign regs_21_io_in = 64'h0; // @[RegFile.scala 75:16:@127229.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@127233.4]
  assign regs_21_io_enable = 1'h1; // @[RegFile.scala 74:20:@127227.4]
  assign regs_22_clock = clock; // @[:@127236.4]
  assign regs_22_reset = io_reset; // @[:@127237.4 RegFile.scala 76:16:@127244.4]
  assign regs_22_io_in = 64'h0; // @[RegFile.scala 75:16:@127243.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@127247.4]
  assign regs_22_io_enable = 1'h1; // @[RegFile.scala 74:20:@127241.4]
  assign regs_23_clock = clock; // @[:@127250.4]
  assign regs_23_reset = io_reset; // @[:@127251.4 RegFile.scala 76:16:@127258.4]
  assign regs_23_io_in = 64'h0; // @[RegFile.scala 75:16:@127257.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@127261.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 74:20:@127255.4]
  assign regs_24_clock = clock; // @[:@127264.4]
  assign regs_24_reset = io_reset; // @[:@127265.4 RegFile.scala 76:16:@127272.4]
  assign regs_24_io_in = 64'h0; // @[RegFile.scala 75:16:@127271.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@127275.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 74:20:@127269.4]
  assign regs_25_clock = clock; // @[:@127278.4]
  assign regs_25_reset = io_reset; // @[:@127279.4 RegFile.scala 76:16:@127286.4]
  assign regs_25_io_in = 64'h0; // @[RegFile.scala 75:16:@127285.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@127289.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 74:20:@127283.4]
  assign regs_26_clock = clock; // @[:@127292.4]
  assign regs_26_reset = io_reset; // @[:@127293.4 RegFile.scala 76:16:@127300.4]
  assign regs_26_io_in = 64'h0; // @[RegFile.scala 75:16:@127299.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@127303.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 74:20:@127297.4]
  assign regs_27_clock = clock; // @[:@127306.4]
  assign regs_27_reset = io_reset; // @[:@127307.4 RegFile.scala 76:16:@127314.4]
  assign regs_27_io_in = 64'h0; // @[RegFile.scala 75:16:@127313.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@127317.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 74:20:@127311.4]
  assign regs_28_clock = clock; // @[:@127320.4]
  assign regs_28_reset = io_reset; // @[:@127321.4 RegFile.scala 76:16:@127328.4]
  assign regs_28_io_in = 64'h0; // @[RegFile.scala 75:16:@127327.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@127331.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 74:20:@127325.4]
  assign regs_29_clock = clock; // @[:@127334.4]
  assign regs_29_reset = io_reset; // @[:@127335.4 RegFile.scala 76:16:@127342.4]
  assign regs_29_io_in = 64'h0; // @[RegFile.scala 75:16:@127341.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@127345.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 74:20:@127339.4]
  assign regs_30_clock = clock; // @[:@127348.4]
  assign regs_30_reset = io_reset; // @[:@127349.4 RegFile.scala 76:16:@127356.4]
  assign regs_30_io_in = 64'h0; // @[RegFile.scala 75:16:@127355.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@127359.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 74:20:@127353.4]
  assign regs_31_clock = clock; // @[:@127362.4]
  assign regs_31_reset = io_reset; // @[:@127363.4 RegFile.scala 76:16:@127370.4]
  assign regs_31_io_in = 64'h0; // @[RegFile.scala 75:16:@127369.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@127373.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 74:20:@127367.4]
  assign regs_32_clock = clock; // @[:@127376.4]
  assign regs_32_reset = io_reset; // @[:@127377.4 RegFile.scala 76:16:@127384.4]
  assign regs_32_io_in = 64'h0; // @[RegFile.scala 75:16:@127383.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@127387.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 74:20:@127381.4]
  assign regs_33_clock = clock; // @[:@127390.4]
  assign regs_33_reset = io_reset; // @[:@127391.4 RegFile.scala 76:16:@127398.4]
  assign regs_33_io_in = 64'h0; // @[RegFile.scala 75:16:@127397.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@127401.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 74:20:@127395.4]
  assign regs_34_clock = clock; // @[:@127404.4]
  assign regs_34_reset = io_reset; // @[:@127405.4 RegFile.scala 76:16:@127412.4]
  assign regs_34_io_in = 64'h0; // @[RegFile.scala 75:16:@127411.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@127415.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 74:20:@127409.4]
  assign regs_35_clock = clock; // @[:@127418.4]
  assign regs_35_reset = io_reset; // @[:@127419.4 RegFile.scala 76:16:@127426.4]
  assign regs_35_io_in = 64'h0; // @[RegFile.scala 75:16:@127425.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@127429.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@127423.4]
  assign regs_36_clock = clock; // @[:@127432.4]
  assign regs_36_reset = io_reset; // @[:@127433.4 RegFile.scala 76:16:@127440.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 75:16:@127439.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@127443.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@127437.4]
  assign regs_37_clock = clock; // @[:@127446.4]
  assign regs_37_reset = io_reset; // @[:@127447.4 RegFile.scala 76:16:@127454.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 75:16:@127453.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@127457.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@127451.4]
  assign regs_38_clock = clock; // @[:@127460.4]
  assign regs_38_reset = io_reset; // @[:@127461.4 RegFile.scala 76:16:@127468.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 75:16:@127467.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@127471.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@127465.4]
  assign regs_39_clock = clock; // @[:@127474.4]
  assign regs_39_reset = io_reset; // @[:@127475.4 RegFile.scala 76:16:@127482.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 75:16:@127481.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@127485.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@127479.4]
  assign regs_40_clock = clock; // @[:@127488.4]
  assign regs_40_reset = io_reset; // @[:@127489.4 RegFile.scala 76:16:@127496.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 75:16:@127495.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@127499.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@127493.4]
  assign regs_41_clock = clock; // @[:@127502.4]
  assign regs_41_reset = io_reset; // @[:@127503.4 RegFile.scala 76:16:@127510.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 75:16:@127509.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@127513.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@127507.4]
  assign regs_42_clock = clock; // @[:@127516.4]
  assign regs_42_reset = io_reset; // @[:@127517.4 RegFile.scala 76:16:@127524.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 75:16:@127523.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@127527.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@127521.4]
  assign regs_43_clock = clock; // @[:@127530.4]
  assign regs_43_reset = io_reset; // @[:@127531.4 RegFile.scala 76:16:@127538.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 75:16:@127537.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@127541.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@127535.4]
  assign regs_44_clock = clock; // @[:@127544.4]
  assign regs_44_reset = io_reset; // @[:@127545.4 RegFile.scala 76:16:@127552.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 75:16:@127551.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@127555.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@127549.4]
  assign regs_45_clock = clock; // @[:@127558.4]
  assign regs_45_reset = io_reset; // @[:@127559.4 RegFile.scala 76:16:@127566.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 75:16:@127565.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@127569.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@127563.4]
  assign regs_46_clock = clock; // @[:@127572.4]
  assign regs_46_reset = io_reset; // @[:@127573.4 RegFile.scala 76:16:@127580.4]
  assign regs_46_io_in = 64'h0; // @[RegFile.scala 75:16:@127579.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@127583.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@127577.4]
  assign regs_47_clock = clock; // @[:@127586.4]
  assign regs_47_reset = io_reset; // @[:@127587.4 RegFile.scala 76:16:@127594.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 75:16:@127593.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@127597.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@127591.4]
  assign regs_48_clock = clock; // @[:@127600.4]
  assign regs_48_reset = io_reset; // @[:@127601.4 RegFile.scala 76:16:@127608.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 75:16:@127607.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@127611.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@127605.4]
  assign regs_49_clock = clock; // @[:@127614.4]
  assign regs_49_reset = io_reset; // @[:@127615.4 RegFile.scala 76:16:@127622.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@127621.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@127625.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@127619.4]
  assign regs_50_clock = clock; // @[:@127628.4]
  assign regs_50_reset = io_reset; // @[:@127629.4 RegFile.scala 76:16:@127636.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@127635.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@127639.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@127633.4]
  assign regs_51_clock = clock; // @[:@127642.4]
  assign regs_51_reset = io_reset; // @[:@127643.4 RegFile.scala 76:16:@127650.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@127649.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@127653.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@127647.4]
  assign regs_52_clock = clock; // @[:@127656.4]
  assign regs_52_reset = io_reset; // @[:@127657.4 RegFile.scala 76:16:@127664.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@127663.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@127667.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@127661.4]
  assign regs_53_clock = clock; // @[:@127670.4]
  assign regs_53_reset = io_reset; // @[:@127671.4 RegFile.scala 76:16:@127678.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@127677.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@127681.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@127675.4]
  assign regs_54_clock = clock; // @[:@127684.4]
  assign regs_54_reset = io_reset; // @[:@127685.4 RegFile.scala 76:16:@127692.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@127691.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@127695.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@127689.4]
  assign regs_55_clock = clock; // @[:@127698.4]
  assign regs_55_reset = io_reset; // @[:@127699.4 RegFile.scala 76:16:@127706.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@127705.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@127709.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@127703.4]
  assign regs_56_clock = clock; // @[:@127712.4]
  assign regs_56_reset = io_reset; // @[:@127713.4 RegFile.scala 76:16:@127720.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@127719.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@127723.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@127717.4]
  assign regs_57_clock = clock; // @[:@127726.4]
  assign regs_57_reset = io_reset; // @[:@127727.4 RegFile.scala 76:16:@127734.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@127733.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@127737.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@127731.4]
  assign regs_58_clock = clock; // @[:@127740.4]
  assign regs_58_reset = io_reset; // @[:@127741.4 RegFile.scala 76:16:@127748.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@127747.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@127751.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@127745.4]
  assign regs_59_clock = clock; // @[:@127754.4]
  assign regs_59_reset = io_reset; // @[:@127755.4 RegFile.scala 76:16:@127762.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 75:16:@127761.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@127765.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@127759.4]
  assign regs_60_clock = clock; // @[:@127768.4]
  assign regs_60_reset = io_reset; // @[:@127769.4 RegFile.scala 76:16:@127776.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@127775.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@127779.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@127773.4]
  assign regs_61_clock = clock; // @[:@127782.4]
  assign regs_61_reset = io_reset; // @[:@127783.4 RegFile.scala 76:16:@127790.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@127789.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@127793.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@127787.4]
  assign regs_62_clock = clock; // @[:@127796.4]
  assign regs_62_reset = io_reset; // @[:@127797.4 RegFile.scala 76:16:@127804.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@127803.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@127807.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@127801.4]
  assign regs_63_clock = clock; // @[:@127810.4]
  assign regs_63_reset = io_reset; // @[:@127811.4 RegFile.scala 76:16:@127818.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@127817.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@127821.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@127815.4]
  assign regs_64_clock = clock; // @[:@127824.4]
  assign regs_64_reset = io_reset; // @[:@127825.4 RegFile.scala 76:16:@127832.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@127831.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@127835.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@127829.4]
  assign regs_65_clock = clock; // @[:@127838.4]
  assign regs_65_reset = io_reset; // @[:@127839.4 RegFile.scala 76:16:@127846.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@127845.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@127849.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@127843.4]
  assign regs_66_clock = clock; // @[:@127852.4]
  assign regs_66_reset = io_reset; // @[:@127853.4 RegFile.scala 76:16:@127860.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@127859.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@127863.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@127857.4]
  assign regs_67_clock = clock; // @[:@127866.4]
  assign regs_67_reset = io_reset; // @[:@127867.4 RegFile.scala 76:16:@127874.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@127873.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@127877.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@127871.4]
  assign regs_68_clock = clock; // @[:@127880.4]
  assign regs_68_reset = io_reset; // @[:@127881.4 RegFile.scala 76:16:@127888.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@127887.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@127891.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@127885.4]
  assign regs_69_clock = clock; // @[:@127894.4]
  assign regs_69_reset = io_reset; // @[:@127895.4 RegFile.scala 76:16:@127902.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@127901.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@127905.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@127899.4]
  assign regs_70_clock = clock; // @[:@127908.4]
  assign regs_70_reset = io_reset; // @[:@127909.4 RegFile.scala 76:16:@127916.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@127915.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@127919.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@127913.4]
  assign regs_71_clock = clock; // @[:@127922.4]
  assign regs_71_reset = io_reset; // @[:@127923.4 RegFile.scala 76:16:@127930.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@127929.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@127933.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@127927.4]
  assign regs_72_clock = clock; // @[:@127936.4]
  assign regs_72_reset = io_reset; // @[:@127937.4 RegFile.scala 76:16:@127944.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@127943.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@127947.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@127941.4]
  assign regs_73_clock = clock; // @[:@127950.4]
  assign regs_73_reset = io_reset; // @[:@127951.4 RegFile.scala 76:16:@127958.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@127957.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@127961.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@127955.4]
  assign regs_74_clock = clock; // @[:@127964.4]
  assign regs_74_reset = io_reset; // @[:@127965.4 RegFile.scala 76:16:@127972.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@127971.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@127975.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@127969.4]
  assign regs_75_clock = clock; // @[:@127978.4]
  assign regs_75_reset = io_reset; // @[:@127979.4 RegFile.scala 76:16:@127986.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@127985.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@127989.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@127983.4]
  assign regs_76_clock = clock; // @[:@127992.4]
  assign regs_76_reset = io_reset; // @[:@127993.4 RegFile.scala 76:16:@128000.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@127999.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@128003.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@127997.4]
  assign regs_77_clock = clock; // @[:@128006.4]
  assign regs_77_reset = io_reset; // @[:@128007.4 RegFile.scala 76:16:@128014.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@128013.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@128017.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@128011.4]
  assign regs_78_clock = clock; // @[:@128020.4]
  assign regs_78_reset = io_reset; // @[:@128021.4 RegFile.scala 76:16:@128028.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@128027.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@128031.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@128025.4]
  assign regs_79_clock = clock; // @[:@128034.4]
  assign regs_79_reset = io_reset; // @[:@128035.4 RegFile.scala 76:16:@128042.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@128041.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@128045.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@128039.4]
  assign regs_80_clock = clock; // @[:@128048.4]
  assign regs_80_reset = io_reset; // @[:@128049.4 RegFile.scala 76:16:@128056.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@128055.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@128059.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@128053.4]
  assign regs_81_clock = clock; // @[:@128062.4]
  assign regs_81_reset = io_reset; // @[:@128063.4 RegFile.scala 76:16:@128070.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@128069.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@128073.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@128067.4]
  assign regs_82_clock = clock; // @[:@128076.4]
  assign regs_82_reset = io_reset; // @[:@128077.4 RegFile.scala 76:16:@128084.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@128083.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@128087.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@128081.4]
  assign regs_83_clock = clock; // @[:@128090.4]
  assign regs_83_reset = io_reset; // @[:@128091.4 RegFile.scala 76:16:@128098.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@128097.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@128101.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@128095.4]
  assign regs_84_clock = clock; // @[:@128104.4]
  assign regs_84_reset = io_reset; // @[:@128105.4 RegFile.scala 76:16:@128112.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@128111.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@128115.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@128109.4]
  assign regs_85_clock = clock; // @[:@128118.4]
  assign regs_85_reset = io_reset; // @[:@128119.4 RegFile.scala 76:16:@128126.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@128125.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@128129.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@128123.4]
  assign regs_86_clock = clock; // @[:@128132.4]
  assign regs_86_reset = io_reset; // @[:@128133.4 RegFile.scala 76:16:@128140.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@128139.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@128143.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@128137.4]
  assign regs_87_clock = clock; // @[:@128146.4]
  assign regs_87_reset = io_reset; // @[:@128147.4 RegFile.scala 76:16:@128154.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@128153.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@128157.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@128151.4]
  assign regs_88_clock = clock; // @[:@128160.4]
  assign regs_88_reset = io_reset; // @[:@128161.4 RegFile.scala 76:16:@128168.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@128167.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@128171.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@128165.4]
  assign regs_89_clock = clock; // @[:@128174.4]
  assign regs_89_reset = io_reset; // @[:@128175.4 RegFile.scala 76:16:@128182.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@128181.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@128185.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@128179.4]
  assign regs_90_clock = clock; // @[:@128188.4]
  assign regs_90_reset = io_reset; // @[:@128189.4 RegFile.scala 76:16:@128196.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@128195.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@128199.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@128193.4]
  assign regs_91_clock = clock; // @[:@128202.4]
  assign regs_91_reset = io_reset; // @[:@128203.4 RegFile.scala 76:16:@128210.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@128209.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@128213.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@128207.4]
  assign regs_92_clock = clock; // @[:@128216.4]
  assign regs_92_reset = io_reset; // @[:@128217.4 RegFile.scala 76:16:@128224.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@128223.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@128227.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@128221.4]
  assign regs_93_clock = clock; // @[:@128230.4]
  assign regs_93_reset = io_reset; // @[:@128231.4 RegFile.scala 76:16:@128238.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@128237.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@128241.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@128235.4]
  assign regs_94_clock = clock; // @[:@128244.4]
  assign regs_94_reset = io_reset; // @[:@128245.4 RegFile.scala 76:16:@128252.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@128251.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@128255.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@128249.4]
  assign regs_95_clock = clock; // @[:@128258.4]
  assign regs_95_reset = io_reset; // @[:@128259.4 RegFile.scala 76:16:@128266.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@128265.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@128269.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@128263.4]
  assign regs_96_clock = clock; // @[:@128272.4]
  assign regs_96_reset = io_reset; // @[:@128273.4 RegFile.scala 76:16:@128280.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@128279.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@128283.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@128277.4]
  assign regs_97_clock = clock; // @[:@128286.4]
  assign regs_97_reset = io_reset; // @[:@128287.4 RegFile.scala 76:16:@128294.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@128293.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@128297.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@128291.4]
  assign regs_98_clock = clock; // @[:@128300.4]
  assign regs_98_reset = io_reset; // @[:@128301.4 RegFile.scala 76:16:@128308.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@128307.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@128311.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@128305.4]
  assign regs_99_clock = clock; // @[:@128314.4]
  assign regs_99_reset = io_reset; // @[:@128315.4 RegFile.scala 76:16:@128322.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@128321.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@128325.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@128319.4]
  assign regs_100_clock = clock; // @[:@128328.4]
  assign regs_100_reset = io_reset; // @[:@128329.4 RegFile.scala 76:16:@128336.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@128335.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@128339.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@128333.4]
  assign regs_101_clock = clock; // @[:@128342.4]
  assign regs_101_reset = io_reset; // @[:@128343.4 RegFile.scala 76:16:@128350.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@128349.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@128353.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@128347.4]
  assign regs_102_clock = clock; // @[:@128356.4]
  assign regs_102_reset = io_reset; // @[:@128357.4 RegFile.scala 76:16:@128364.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@128363.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@128367.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@128361.4]
  assign regs_103_clock = clock; // @[:@128370.4]
  assign regs_103_reset = io_reset; // @[:@128371.4 RegFile.scala 76:16:@128378.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@128377.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@128381.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@128375.4]
  assign regs_104_clock = clock; // @[:@128384.4]
  assign regs_104_reset = io_reset; // @[:@128385.4 RegFile.scala 76:16:@128392.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@128391.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@128395.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@128389.4]
  assign regs_105_clock = clock; // @[:@128398.4]
  assign regs_105_reset = io_reset; // @[:@128399.4 RegFile.scala 76:16:@128406.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@128405.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@128409.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@128403.4]
  assign regs_106_clock = clock; // @[:@128412.4]
  assign regs_106_reset = io_reset; // @[:@128413.4 RegFile.scala 76:16:@128420.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@128419.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@128423.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@128417.4]
  assign regs_107_clock = clock; // @[:@128426.4]
  assign regs_107_reset = io_reset; // @[:@128427.4 RegFile.scala 76:16:@128434.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@128433.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@128437.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@128431.4]
  assign regs_108_clock = clock; // @[:@128440.4]
  assign regs_108_reset = io_reset; // @[:@128441.4 RegFile.scala 76:16:@128448.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@128447.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@128451.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@128445.4]
  assign regs_109_clock = clock; // @[:@128454.4]
  assign regs_109_reset = io_reset; // @[:@128455.4 RegFile.scala 76:16:@128462.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@128461.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@128465.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@128459.4]
  assign regs_110_clock = clock; // @[:@128468.4]
  assign regs_110_reset = io_reset; // @[:@128469.4 RegFile.scala 76:16:@128476.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@128475.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@128479.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@128473.4]
  assign regs_111_clock = clock; // @[:@128482.4]
  assign regs_111_reset = io_reset; // @[:@128483.4 RegFile.scala 76:16:@128490.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@128489.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@128493.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@128487.4]
  assign regs_112_clock = clock; // @[:@128496.4]
  assign regs_112_reset = io_reset; // @[:@128497.4 RegFile.scala 76:16:@128504.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@128503.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@128507.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@128501.4]
  assign regs_113_clock = clock; // @[:@128510.4]
  assign regs_113_reset = io_reset; // @[:@128511.4 RegFile.scala 76:16:@128518.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@128517.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@128521.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@128515.4]
  assign regs_114_clock = clock; // @[:@128524.4]
  assign regs_114_reset = io_reset; // @[:@128525.4 RegFile.scala 76:16:@128532.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@128531.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@128535.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@128529.4]
  assign regs_115_clock = clock; // @[:@128538.4]
  assign regs_115_reset = io_reset; // @[:@128539.4 RegFile.scala 76:16:@128546.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@128545.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@128549.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@128543.4]
  assign regs_116_clock = clock; // @[:@128552.4]
  assign regs_116_reset = io_reset; // @[:@128553.4 RegFile.scala 76:16:@128560.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@128559.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@128563.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@128557.4]
  assign regs_117_clock = clock; // @[:@128566.4]
  assign regs_117_reset = io_reset; // @[:@128567.4 RegFile.scala 76:16:@128574.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@128573.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@128577.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@128571.4]
  assign regs_118_clock = clock; // @[:@128580.4]
  assign regs_118_reset = io_reset; // @[:@128581.4 RegFile.scala 76:16:@128588.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@128587.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@128591.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@128585.4]
  assign regs_119_clock = clock; // @[:@128594.4]
  assign regs_119_reset = io_reset; // @[:@128595.4 RegFile.scala 76:16:@128602.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@128601.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@128605.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@128599.4]
  assign regs_120_clock = clock; // @[:@128608.4]
  assign regs_120_reset = io_reset; // @[:@128609.4 RegFile.scala 76:16:@128616.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@128615.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@128619.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@128613.4]
  assign regs_121_clock = clock; // @[:@128622.4]
  assign regs_121_reset = io_reset; // @[:@128623.4 RegFile.scala 76:16:@128630.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@128629.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@128633.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@128627.4]
  assign regs_122_clock = clock; // @[:@128636.4]
  assign regs_122_reset = io_reset; // @[:@128637.4 RegFile.scala 76:16:@128644.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@128643.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@128647.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@128641.4]
  assign regs_123_clock = clock; // @[:@128650.4]
  assign regs_123_reset = io_reset; // @[:@128651.4 RegFile.scala 76:16:@128658.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@128657.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@128661.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@128655.4]
  assign regs_124_clock = clock; // @[:@128664.4]
  assign regs_124_reset = io_reset; // @[:@128665.4 RegFile.scala 76:16:@128672.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@128671.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@128675.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@128669.4]
  assign regs_125_clock = clock; // @[:@128678.4]
  assign regs_125_reset = io_reset; // @[:@128679.4 RegFile.scala 76:16:@128686.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@128685.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@128689.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@128683.4]
  assign regs_126_clock = clock; // @[:@128692.4]
  assign regs_126_reset = io_reset; // @[:@128693.4 RegFile.scala 76:16:@128700.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@128699.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@128703.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@128697.4]
  assign regs_127_clock = clock; // @[:@128706.4]
  assign regs_127_reset = io_reset; // @[:@128707.4 RegFile.scala 76:16:@128714.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@128713.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@128717.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@128711.4]
  assign regs_128_clock = clock; // @[:@128720.4]
  assign regs_128_reset = io_reset; // @[:@128721.4 RegFile.scala 76:16:@128728.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@128727.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@128731.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@128725.4]
  assign regs_129_clock = clock; // @[:@128734.4]
  assign regs_129_reset = io_reset; // @[:@128735.4 RegFile.scala 76:16:@128742.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@128741.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@128745.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@128739.4]
  assign regs_130_clock = clock; // @[:@128748.4]
  assign regs_130_reset = io_reset; // @[:@128749.4 RegFile.scala 76:16:@128756.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@128755.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@128759.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@128753.4]
  assign regs_131_clock = clock; // @[:@128762.4]
  assign regs_131_reset = io_reset; // @[:@128763.4 RegFile.scala 76:16:@128770.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@128769.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@128773.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@128767.4]
  assign regs_132_clock = clock; // @[:@128776.4]
  assign regs_132_reset = io_reset; // @[:@128777.4 RegFile.scala 76:16:@128784.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@128783.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@128787.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@128781.4]
  assign regs_133_clock = clock; // @[:@128790.4]
  assign regs_133_reset = io_reset; // @[:@128791.4 RegFile.scala 76:16:@128798.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@128797.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@128801.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@128795.4]
  assign regs_134_clock = clock; // @[:@128804.4]
  assign regs_134_reset = io_reset; // @[:@128805.4 RegFile.scala 76:16:@128812.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@128811.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@128815.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@128809.4]
  assign regs_135_clock = clock; // @[:@128818.4]
  assign regs_135_reset = io_reset; // @[:@128819.4 RegFile.scala 76:16:@128826.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@128825.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@128829.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@128823.4]
  assign regs_136_clock = clock; // @[:@128832.4]
  assign regs_136_reset = io_reset; // @[:@128833.4 RegFile.scala 76:16:@128840.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@128839.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@128843.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@128837.4]
  assign regs_137_clock = clock; // @[:@128846.4]
  assign regs_137_reset = io_reset; // @[:@128847.4 RegFile.scala 76:16:@128854.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@128853.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@128857.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@128851.4]
  assign regs_138_clock = clock; // @[:@128860.4]
  assign regs_138_reset = io_reset; // @[:@128861.4 RegFile.scala 76:16:@128868.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@128867.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@128871.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@128865.4]
  assign regs_139_clock = clock; // @[:@128874.4]
  assign regs_139_reset = io_reset; // @[:@128875.4 RegFile.scala 76:16:@128882.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@128881.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@128885.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@128879.4]
  assign regs_140_clock = clock; // @[:@128888.4]
  assign regs_140_reset = io_reset; // @[:@128889.4 RegFile.scala 76:16:@128896.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@128895.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@128899.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@128893.4]
  assign regs_141_clock = clock; // @[:@128902.4]
  assign regs_141_reset = io_reset; // @[:@128903.4 RegFile.scala 76:16:@128910.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@128909.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@128913.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@128907.4]
  assign regs_142_clock = clock; // @[:@128916.4]
  assign regs_142_reset = io_reset; // @[:@128917.4 RegFile.scala 76:16:@128924.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@128923.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@128927.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@128921.4]
  assign regs_143_clock = clock; // @[:@128930.4]
  assign regs_143_reset = io_reset; // @[:@128931.4 RegFile.scala 76:16:@128938.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@128937.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@128941.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@128935.4]
  assign regs_144_clock = clock; // @[:@128944.4]
  assign regs_144_reset = io_reset; // @[:@128945.4 RegFile.scala 76:16:@128952.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@128951.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@128955.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@128949.4]
  assign regs_145_clock = clock; // @[:@128958.4]
  assign regs_145_reset = io_reset; // @[:@128959.4 RegFile.scala 76:16:@128966.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@128965.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@128969.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@128963.4]
  assign regs_146_clock = clock; // @[:@128972.4]
  assign regs_146_reset = io_reset; // @[:@128973.4 RegFile.scala 76:16:@128980.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@128979.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@128983.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@128977.4]
  assign regs_147_clock = clock; // @[:@128986.4]
  assign regs_147_reset = io_reset; // @[:@128987.4 RegFile.scala 76:16:@128994.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@128993.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@128997.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@128991.4]
  assign regs_148_clock = clock; // @[:@129000.4]
  assign regs_148_reset = io_reset; // @[:@129001.4 RegFile.scala 76:16:@129008.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@129007.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@129011.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@129005.4]
  assign regs_149_clock = clock; // @[:@129014.4]
  assign regs_149_reset = io_reset; // @[:@129015.4 RegFile.scala 76:16:@129022.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@129021.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@129025.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@129019.4]
  assign regs_150_clock = clock; // @[:@129028.4]
  assign regs_150_reset = io_reset; // @[:@129029.4 RegFile.scala 76:16:@129036.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@129035.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@129039.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@129033.4]
  assign regs_151_clock = clock; // @[:@129042.4]
  assign regs_151_reset = io_reset; // @[:@129043.4 RegFile.scala 76:16:@129050.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@129049.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@129053.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@129047.4]
  assign regs_152_clock = clock; // @[:@129056.4]
  assign regs_152_reset = io_reset; // @[:@129057.4 RegFile.scala 76:16:@129064.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@129063.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@129067.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@129061.4]
  assign regs_153_clock = clock; // @[:@129070.4]
  assign regs_153_reset = io_reset; // @[:@129071.4 RegFile.scala 76:16:@129078.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@129077.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@129081.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@129075.4]
  assign regs_154_clock = clock; // @[:@129084.4]
  assign regs_154_reset = io_reset; // @[:@129085.4 RegFile.scala 76:16:@129092.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@129091.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@129095.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@129089.4]
  assign regs_155_clock = clock; // @[:@129098.4]
  assign regs_155_reset = io_reset; // @[:@129099.4 RegFile.scala 76:16:@129106.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@129105.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@129109.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@129103.4]
  assign regs_156_clock = clock; // @[:@129112.4]
  assign regs_156_reset = io_reset; // @[:@129113.4 RegFile.scala 76:16:@129120.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@129119.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@129123.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@129117.4]
  assign regs_157_clock = clock; // @[:@129126.4]
  assign regs_157_reset = io_reset; // @[:@129127.4 RegFile.scala 76:16:@129134.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@129133.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@129137.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@129131.4]
  assign regs_158_clock = clock; // @[:@129140.4]
  assign regs_158_reset = io_reset; // @[:@129141.4 RegFile.scala 76:16:@129148.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@129147.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@129151.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@129145.4]
  assign regs_159_clock = clock; // @[:@129154.4]
  assign regs_159_reset = io_reset; // @[:@129155.4 RegFile.scala 76:16:@129162.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@129161.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@129165.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@129159.4]
  assign regs_160_clock = clock; // @[:@129168.4]
  assign regs_160_reset = io_reset; // @[:@129169.4 RegFile.scala 76:16:@129176.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@129175.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@129179.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@129173.4]
  assign regs_161_clock = clock; // @[:@129182.4]
  assign regs_161_reset = io_reset; // @[:@129183.4 RegFile.scala 76:16:@129190.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@129189.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@129193.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@129187.4]
  assign regs_162_clock = clock; // @[:@129196.4]
  assign regs_162_reset = io_reset; // @[:@129197.4 RegFile.scala 76:16:@129204.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@129203.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@129207.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@129201.4]
  assign regs_163_clock = clock; // @[:@129210.4]
  assign regs_163_reset = io_reset; // @[:@129211.4 RegFile.scala 76:16:@129218.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@129217.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@129221.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@129215.4]
  assign regs_164_clock = clock; // @[:@129224.4]
  assign regs_164_reset = io_reset; // @[:@129225.4 RegFile.scala 76:16:@129232.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@129231.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@129235.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@129229.4]
  assign regs_165_clock = clock; // @[:@129238.4]
  assign regs_165_reset = io_reset; // @[:@129239.4 RegFile.scala 76:16:@129246.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@129245.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@129249.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@129243.4]
  assign regs_166_clock = clock; // @[:@129252.4]
  assign regs_166_reset = io_reset; // @[:@129253.4 RegFile.scala 76:16:@129260.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@129259.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@129263.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@129257.4]
  assign regs_167_clock = clock; // @[:@129266.4]
  assign regs_167_reset = io_reset; // @[:@129267.4 RegFile.scala 76:16:@129274.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@129273.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@129277.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@129271.4]
  assign regs_168_clock = clock; // @[:@129280.4]
  assign regs_168_reset = io_reset; // @[:@129281.4 RegFile.scala 76:16:@129288.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@129287.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@129291.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@129285.4]
  assign regs_169_clock = clock; // @[:@129294.4]
  assign regs_169_reset = io_reset; // @[:@129295.4 RegFile.scala 76:16:@129302.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@129301.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@129305.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@129299.4]
  assign regs_170_clock = clock; // @[:@129308.4]
  assign regs_170_reset = io_reset; // @[:@129309.4 RegFile.scala 76:16:@129316.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@129315.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@129319.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@129313.4]
  assign regs_171_clock = clock; // @[:@129322.4]
  assign regs_171_reset = io_reset; // @[:@129323.4 RegFile.scala 76:16:@129330.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@129329.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@129333.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@129327.4]
  assign regs_172_clock = clock; // @[:@129336.4]
  assign regs_172_reset = io_reset; // @[:@129337.4 RegFile.scala 76:16:@129344.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@129343.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@129347.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@129341.4]
  assign regs_173_clock = clock; // @[:@129350.4]
  assign regs_173_reset = io_reset; // @[:@129351.4 RegFile.scala 76:16:@129358.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@129357.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@129361.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@129355.4]
  assign regs_174_clock = clock; // @[:@129364.4]
  assign regs_174_reset = io_reset; // @[:@129365.4 RegFile.scala 76:16:@129372.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@129371.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@129375.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@129369.4]
  assign regs_175_clock = clock; // @[:@129378.4]
  assign regs_175_reset = io_reset; // @[:@129379.4 RegFile.scala 76:16:@129386.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@129385.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@129389.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@129383.4]
  assign regs_176_clock = clock; // @[:@129392.4]
  assign regs_176_reset = io_reset; // @[:@129393.4 RegFile.scala 76:16:@129400.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@129399.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@129403.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@129397.4]
  assign regs_177_clock = clock; // @[:@129406.4]
  assign regs_177_reset = io_reset; // @[:@129407.4 RegFile.scala 76:16:@129414.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@129413.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@129417.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@129411.4]
  assign regs_178_clock = clock; // @[:@129420.4]
  assign regs_178_reset = io_reset; // @[:@129421.4 RegFile.scala 76:16:@129428.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@129427.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@129431.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@129425.4]
  assign regs_179_clock = clock; // @[:@129434.4]
  assign regs_179_reset = io_reset; // @[:@129435.4 RegFile.scala 76:16:@129442.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@129441.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@129445.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@129439.4]
  assign regs_180_clock = clock; // @[:@129448.4]
  assign regs_180_reset = io_reset; // @[:@129449.4 RegFile.scala 76:16:@129456.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@129455.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@129459.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@129453.4]
  assign regs_181_clock = clock; // @[:@129462.4]
  assign regs_181_reset = io_reset; // @[:@129463.4 RegFile.scala 76:16:@129470.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@129469.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@129473.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@129467.4]
  assign regs_182_clock = clock; // @[:@129476.4]
  assign regs_182_reset = io_reset; // @[:@129477.4 RegFile.scala 76:16:@129484.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@129483.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@129487.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@129481.4]
  assign regs_183_clock = clock; // @[:@129490.4]
  assign regs_183_reset = io_reset; // @[:@129491.4 RegFile.scala 76:16:@129498.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@129497.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@129501.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@129495.4]
  assign regs_184_clock = clock; // @[:@129504.4]
  assign regs_184_reset = io_reset; // @[:@129505.4 RegFile.scala 76:16:@129512.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@129511.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@129515.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@129509.4]
  assign regs_185_clock = clock; // @[:@129518.4]
  assign regs_185_reset = io_reset; // @[:@129519.4 RegFile.scala 76:16:@129526.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@129525.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@129529.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@129523.4]
  assign regs_186_clock = clock; // @[:@129532.4]
  assign regs_186_reset = io_reset; // @[:@129533.4 RegFile.scala 76:16:@129540.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@129539.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@129543.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@129537.4]
  assign regs_187_clock = clock; // @[:@129546.4]
  assign regs_187_reset = io_reset; // @[:@129547.4 RegFile.scala 76:16:@129554.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@129553.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@129557.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@129551.4]
  assign regs_188_clock = clock; // @[:@129560.4]
  assign regs_188_reset = io_reset; // @[:@129561.4 RegFile.scala 76:16:@129568.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@129567.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@129571.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@129565.4]
  assign regs_189_clock = clock; // @[:@129574.4]
  assign regs_189_reset = io_reset; // @[:@129575.4 RegFile.scala 76:16:@129582.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@129581.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@129585.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@129579.4]
  assign regs_190_clock = clock; // @[:@129588.4]
  assign regs_190_reset = io_reset; // @[:@129589.4 RegFile.scala 76:16:@129596.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@129595.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@129599.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@129593.4]
  assign regs_191_clock = clock; // @[:@129602.4]
  assign regs_191_reset = io_reset; // @[:@129603.4 RegFile.scala 76:16:@129610.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@129609.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@129613.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@129607.4]
  assign regs_192_clock = clock; // @[:@129616.4]
  assign regs_192_reset = io_reset; // @[:@129617.4 RegFile.scala 76:16:@129624.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@129623.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@129627.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@129621.4]
  assign regs_193_clock = clock; // @[:@129630.4]
  assign regs_193_reset = io_reset; // @[:@129631.4 RegFile.scala 76:16:@129638.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@129637.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@129641.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@129635.4]
  assign regs_194_clock = clock; // @[:@129644.4]
  assign regs_194_reset = io_reset; // @[:@129645.4 RegFile.scala 76:16:@129652.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@129651.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@129655.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@129649.4]
  assign regs_195_clock = clock; // @[:@129658.4]
  assign regs_195_reset = io_reset; // @[:@129659.4 RegFile.scala 76:16:@129666.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@129665.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@129669.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@129663.4]
  assign regs_196_clock = clock; // @[:@129672.4]
  assign regs_196_reset = io_reset; // @[:@129673.4 RegFile.scala 76:16:@129680.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@129679.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@129683.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@129677.4]
  assign regs_197_clock = clock; // @[:@129686.4]
  assign regs_197_reset = io_reset; // @[:@129687.4 RegFile.scala 76:16:@129694.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@129693.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@129697.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@129691.4]
  assign regs_198_clock = clock; // @[:@129700.4]
  assign regs_198_reset = io_reset; // @[:@129701.4 RegFile.scala 76:16:@129708.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@129707.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@129711.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@129705.4]
  assign regs_199_clock = clock; // @[:@129714.4]
  assign regs_199_reset = io_reset; // @[:@129715.4 RegFile.scala 76:16:@129722.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@129721.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@129725.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@129719.4]
  assign regs_200_clock = clock; // @[:@129728.4]
  assign regs_200_reset = io_reset; // @[:@129729.4 RegFile.scala 76:16:@129736.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@129735.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@129739.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@129733.4]
  assign regs_201_clock = clock; // @[:@129742.4]
  assign regs_201_reset = io_reset; // @[:@129743.4 RegFile.scala 76:16:@129750.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@129749.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@129753.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@129747.4]
  assign regs_202_clock = clock; // @[:@129756.4]
  assign regs_202_reset = io_reset; // @[:@129757.4 RegFile.scala 76:16:@129764.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@129763.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@129767.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@129761.4]
  assign regs_203_clock = clock; // @[:@129770.4]
  assign regs_203_reset = io_reset; // @[:@129771.4 RegFile.scala 76:16:@129778.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@129777.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@129781.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@129775.4]
  assign regs_204_clock = clock; // @[:@129784.4]
  assign regs_204_reset = io_reset; // @[:@129785.4 RegFile.scala 76:16:@129792.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@129791.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@129795.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@129789.4]
  assign regs_205_clock = clock; // @[:@129798.4]
  assign regs_205_reset = io_reset; // @[:@129799.4 RegFile.scala 76:16:@129806.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@129805.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@129809.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@129803.4]
  assign regs_206_clock = clock; // @[:@129812.4]
  assign regs_206_reset = io_reset; // @[:@129813.4 RegFile.scala 76:16:@129820.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@129819.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@129823.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@129817.4]
  assign regs_207_clock = clock; // @[:@129826.4]
  assign regs_207_reset = io_reset; // @[:@129827.4 RegFile.scala 76:16:@129834.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@129833.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@129837.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@129831.4]
  assign regs_208_clock = clock; // @[:@129840.4]
  assign regs_208_reset = io_reset; // @[:@129841.4 RegFile.scala 76:16:@129848.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@129847.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@129851.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@129845.4]
  assign regs_209_clock = clock; // @[:@129854.4]
  assign regs_209_reset = io_reset; // @[:@129855.4 RegFile.scala 76:16:@129862.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@129861.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@129865.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@129859.4]
  assign regs_210_clock = clock; // @[:@129868.4]
  assign regs_210_reset = io_reset; // @[:@129869.4 RegFile.scala 76:16:@129876.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@129875.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@129879.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@129873.4]
  assign regs_211_clock = clock; // @[:@129882.4]
  assign regs_211_reset = io_reset; // @[:@129883.4 RegFile.scala 76:16:@129890.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@129889.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@129893.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@129887.4]
  assign regs_212_clock = clock; // @[:@129896.4]
  assign regs_212_reset = io_reset; // @[:@129897.4 RegFile.scala 76:16:@129904.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@129903.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@129907.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@129901.4]
  assign regs_213_clock = clock; // @[:@129910.4]
  assign regs_213_reset = io_reset; // @[:@129911.4 RegFile.scala 76:16:@129918.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@129917.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@129921.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@129915.4]
  assign regs_214_clock = clock; // @[:@129924.4]
  assign regs_214_reset = io_reset; // @[:@129925.4 RegFile.scala 76:16:@129932.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@129931.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@129935.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@129929.4]
  assign regs_215_clock = clock; // @[:@129938.4]
  assign regs_215_reset = io_reset; // @[:@129939.4 RegFile.scala 76:16:@129946.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@129945.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@129949.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@129943.4]
  assign regs_216_clock = clock; // @[:@129952.4]
  assign regs_216_reset = io_reset; // @[:@129953.4 RegFile.scala 76:16:@129960.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@129959.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@129963.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@129957.4]
  assign regs_217_clock = clock; // @[:@129966.4]
  assign regs_217_reset = io_reset; // @[:@129967.4 RegFile.scala 76:16:@129974.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@129973.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@129977.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@129971.4]
  assign regs_218_clock = clock; // @[:@129980.4]
  assign regs_218_reset = io_reset; // @[:@129981.4 RegFile.scala 76:16:@129988.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@129987.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@129991.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@129985.4]
  assign regs_219_clock = clock; // @[:@129994.4]
  assign regs_219_reset = io_reset; // @[:@129995.4 RegFile.scala 76:16:@130002.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@130001.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@130005.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@129999.4]
  assign regs_220_clock = clock; // @[:@130008.4]
  assign regs_220_reset = io_reset; // @[:@130009.4 RegFile.scala 76:16:@130016.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@130015.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@130019.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@130013.4]
  assign regs_221_clock = clock; // @[:@130022.4]
  assign regs_221_reset = io_reset; // @[:@130023.4 RegFile.scala 76:16:@130030.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@130029.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@130033.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@130027.4]
  assign regs_222_clock = clock; // @[:@130036.4]
  assign regs_222_reset = io_reset; // @[:@130037.4 RegFile.scala 76:16:@130044.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@130043.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@130047.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@130041.4]
  assign regs_223_clock = clock; // @[:@130050.4]
  assign regs_223_reset = io_reset; // @[:@130051.4 RegFile.scala 76:16:@130058.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@130057.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@130061.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@130055.4]
  assign regs_224_clock = clock; // @[:@130064.4]
  assign regs_224_reset = io_reset; // @[:@130065.4 RegFile.scala 76:16:@130072.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@130071.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@130075.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@130069.4]
  assign regs_225_clock = clock; // @[:@130078.4]
  assign regs_225_reset = io_reset; // @[:@130079.4 RegFile.scala 76:16:@130086.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@130085.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@130089.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@130083.4]
  assign regs_226_clock = clock; // @[:@130092.4]
  assign regs_226_reset = io_reset; // @[:@130093.4 RegFile.scala 76:16:@130100.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@130099.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@130103.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@130097.4]
  assign regs_227_clock = clock; // @[:@130106.4]
  assign regs_227_reset = io_reset; // @[:@130107.4 RegFile.scala 76:16:@130114.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@130113.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@130117.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@130111.4]
  assign regs_228_clock = clock; // @[:@130120.4]
  assign regs_228_reset = io_reset; // @[:@130121.4 RegFile.scala 76:16:@130128.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@130127.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@130131.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@130125.4]
  assign regs_229_clock = clock; // @[:@130134.4]
  assign regs_229_reset = io_reset; // @[:@130135.4 RegFile.scala 76:16:@130142.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@130141.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@130145.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@130139.4]
  assign regs_230_clock = clock; // @[:@130148.4]
  assign regs_230_reset = io_reset; // @[:@130149.4 RegFile.scala 76:16:@130156.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@130155.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@130159.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@130153.4]
  assign regs_231_clock = clock; // @[:@130162.4]
  assign regs_231_reset = io_reset; // @[:@130163.4 RegFile.scala 76:16:@130170.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@130169.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@130173.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@130167.4]
  assign regs_232_clock = clock; // @[:@130176.4]
  assign regs_232_reset = io_reset; // @[:@130177.4 RegFile.scala 76:16:@130184.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@130183.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@130187.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@130181.4]
  assign regs_233_clock = clock; // @[:@130190.4]
  assign regs_233_reset = io_reset; // @[:@130191.4 RegFile.scala 76:16:@130198.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@130197.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@130201.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@130195.4]
  assign regs_234_clock = clock; // @[:@130204.4]
  assign regs_234_reset = io_reset; // @[:@130205.4 RegFile.scala 76:16:@130212.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@130211.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@130215.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@130209.4]
  assign regs_235_clock = clock; // @[:@130218.4]
  assign regs_235_reset = io_reset; // @[:@130219.4 RegFile.scala 76:16:@130226.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@130225.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@130229.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@130223.4]
  assign regs_236_clock = clock; // @[:@130232.4]
  assign regs_236_reset = io_reset; // @[:@130233.4 RegFile.scala 76:16:@130240.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@130239.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@130243.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@130237.4]
  assign regs_237_clock = clock; // @[:@130246.4]
  assign regs_237_reset = io_reset; // @[:@130247.4 RegFile.scala 76:16:@130254.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@130253.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@130257.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@130251.4]
  assign regs_238_clock = clock; // @[:@130260.4]
  assign regs_238_reset = io_reset; // @[:@130261.4 RegFile.scala 76:16:@130268.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@130267.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@130271.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@130265.4]
  assign regs_239_clock = clock; // @[:@130274.4]
  assign regs_239_reset = io_reset; // @[:@130275.4 RegFile.scala 76:16:@130282.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@130281.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@130285.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@130279.4]
  assign regs_240_clock = clock; // @[:@130288.4]
  assign regs_240_reset = io_reset; // @[:@130289.4 RegFile.scala 76:16:@130296.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@130295.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@130299.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@130293.4]
  assign regs_241_clock = clock; // @[:@130302.4]
  assign regs_241_reset = io_reset; // @[:@130303.4 RegFile.scala 76:16:@130310.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@130309.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@130313.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@130307.4]
  assign regs_242_clock = clock; // @[:@130316.4]
  assign regs_242_reset = io_reset; // @[:@130317.4 RegFile.scala 76:16:@130324.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@130323.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@130327.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@130321.4]
  assign regs_243_clock = clock; // @[:@130330.4]
  assign regs_243_reset = io_reset; // @[:@130331.4 RegFile.scala 76:16:@130338.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@130337.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@130341.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@130335.4]
  assign regs_244_clock = clock; // @[:@130344.4]
  assign regs_244_reset = io_reset; // @[:@130345.4 RegFile.scala 76:16:@130352.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@130351.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@130355.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@130349.4]
  assign regs_245_clock = clock; // @[:@130358.4]
  assign regs_245_reset = io_reset; // @[:@130359.4 RegFile.scala 76:16:@130366.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@130365.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@130369.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@130363.4]
  assign regs_246_clock = clock; // @[:@130372.4]
  assign regs_246_reset = io_reset; // @[:@130373.4 RegFile.scala 76:16:@130380.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@130379.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@130383.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@130377.4]
  assign regs_247_clock = clock; // @[:@130386.4]
  assign regs_247_reset = io_reset; // @[:@130387.4 RegFile.scala 76:16:@130394.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@130393.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@130397.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@130391.4]
  assign regs_248_clock = clock; // @[:@130400.4]
  assign regs_248_reset = io_reset; // @[:@130401.4 RegFile.scala 76:16:@130408.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@130407.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@130411.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@130405.4]
  assign regs_249_clock = clock; // @[:@130414.4]
  assign regs_249_reset = io_reset; // @[:@130415.4 RegFile.scala 76:16:@130422.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@130421.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@130425.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@130419.4]
  assign regs_250_clock = clock; // @[:@130428.4]
  assign regs_250_reset = io_reset; // @[:@130429.4 RegFile.scala 76:16:@130436.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@130435.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@130439.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@130433.4]
  assign regs_251_clock = clock; // @[:@130442.4]
  assign regs_251_reset = io_reset; // @[:@130443.4 RegFile.scala 76:16:@130450.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@130449.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@130453.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@130447.4]
  assign regs_252_clock = clock; // @[:@130456.4]
  assign regs_252_reset = io_reset; // @[:@130457.4 RegFile.scala 76:16:@130464.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@130463.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@130467.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@130461.4]
  assign regs_253_clock = clock; // @[:@130470.4]
  assign regs_253_reset = io_reset; // @[:@130471.4 RegFile.scala 76:16:@130478.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@130477.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@130481.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@130475.4]
  assign regs_254_clock = clock; // @[:@130484.4]
  assign regs_254_reset = io_reset; // @[:@130485.4 RegFile.scala 76:16:@130492.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@130491.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@130495.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@130489.4]
  assign regs_255_clock = clock; // @[:@130498.4]
  assign regs_255_reset = io_reset; // @[:@130499.4 RegFile.scala 76:16:@130506.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@130505.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@130509.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@130503.4]
  assign regs_256_clock = clock; // @[:@130512.4]
  assign regs_256_reset = io_reset; // @[:@130513.4 RegFile.scala 76:16:@130520.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@130519.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@130523.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@130517.4]
  assign regs_257_clock = clock; // @[:@130526.4]
  assign regs_257_reset = io_reset; // @[:@130527.4 RegFile.scala 76:16:@130534.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@130533.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@130537.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@130531.4]
  assign regs_258_clock = clock; // @[:@130540.4]
  assign regs_258_reset = io_reset; // @[:@130541.4 RegFile.scala 76:16:@130548.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@130547.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@130551.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@130545.4]
  assign regs_259_clock = clock; // @[:@130554.4]
  assign regs_259_reset = io_reset; // @[:@130555.4 RegFile.scala 76:16:@130562.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@130561.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@130565.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@130559.4]
  assign regs_260_clock = clock; // @[:@130568.4]
  assign regs_260_reset = io_reset; // @[:@130569.4 RegFile.scala 76:16:@130576.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@130575.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@130579.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@130573.4]
  assign regs_261_clock = clock; // @[:@130582.4]
  assign regs_261_reset = io_reset; // @[:@130583.4 RegFile.scala 76:16:@130590.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@130589.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@130593.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@130587.4]
  assign regs_262_clock = clock; // @[:@130596.4]
  assign regs_262_reset = io_reset; // @[:@130597.4 RegFile.scala 76:16:@130604.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@130603.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@130607.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@130601.4]
  assign regs_263_clock = clock; // @[:@130610.4]
  assign regs_263_reset = io_reset; // @[:@130611.4 RegFile.scala 76:16:@130618.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@130617.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@130621.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@130615.4]
  assign regs_264_clock = clock; // @[:@130624.4]
  assign regs_264_reset = io_reset; // @[:@130625.4 RegFile.scala 76:16:@130632.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@130631.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@130635.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@130629.4]
  assign regs_265_clock = clock; // @[:@130638.4]
  assign regs_265_reset = io_reset; // @[:@130639.4 RegFile.scala 76:16:@130646.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@130645.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@130649.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@130643.4]
  assign regs_266_clock = clock; // @[:@130652.4]
  assign regs_266_reset = io_reset; // @[:@130653.4 RegFile.scala 76:16:@130660.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@130659.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@130663.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@130657.4]
  assign regs_267_clock = clock; // @[:@130666.4]
  assign regs_267_reset = io_reset; // @[:@130667.4 RegFile.scala 76:16:@130674.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@130673.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@130677.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@130671.4]
  assign regs_268_clock = clock; // @[:@130680.4]
  assign regs_268_reset = io_reset; // @[:@130681.4 RegFile.scala 76:16:@130688.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@130687.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@130691.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@130685.4]
  assign regs_269_clock = clock; // @[:@130694.4]
  assign regs_269_reset = io_reset; // @[:@130695.4 RegFile.scala 76:16:@130702.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@130701.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@130705.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@130699.4]
  assign regs_270_clock = clock; // @[:@130708.4]
  assign regs_270_reset = io_reset; // @[:@130709.4 RegFile.scala 76:16:@130716.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@130715.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@130719.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@130713.4]
  assign regs_271_clock = clock; // @[:@130722.4]
  assign regs_271_reset = io_reset; // @[:@130723.4 RegFile.scala 76:16:@130730.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@130729.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@130733.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@130727.4]
  assign regs_272_clock = clock; // @[:@130736.4]
  assign regs_272_reset = io_reset; // @[:@130737.4 RegFile.scala 76:16:@130744.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@130743.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@130747.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@130741.4]
  assign regs_273_clock = clock; // @[:@130750.4]
  assign regs_273_reset = io_reset; // @[:@130751.4 RegFile.scala 76:16:@130758.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@130757.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@130761.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@130755.4]
  assign regs_274_clock = clock; // @[:@130764.4]
  assign regs_274_reset = io_reset; // @[:@130765.4 RegFile.scala 76:16:@130772.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@130771.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@130775.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@130769.4]
  assign regs_275_clock = clock; // @[:@130778.4]
  assign regs_275_reset = io_reset; // @[:@130779.4 RegFile.scala 76:16:@130786.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@130785.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@130789.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@130783.4]
  assign regs_276_clock = clock; // @[:@130792.4]
  assign regs_276_reset = io_reset; // @[:@130793.4 RegFile.scala 76:16:@130800.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@130799.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@130803.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@130797.4]
  assign regs_277_clock = clock; // @[:@130806.4]
  assign regs_277_reset = io_reset; // @[:@130807.4 RegFile.scala 76:16:@130814.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@130813.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@130817.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@130811.4]
  assign regs_278_clock = clock; // @[:@130820.4]
  assign regs_278_reset = io_reset; // @[:@130821.4 RegFile.scala 76:16:@130828.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@130827.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@130831.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@130825.4]
  assign regs_279_clock = clock; // @[:@130834.4]
  assign regs_279_reset = io_reset; // @[:@130835.4 RegFile.scala 76:16:@130842.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@130841.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@130845.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@130839.4]
  assign regs_280_clock = clock; // @[:@130848.4]
  assign regs_280_reset = io_reset; // @[:@130849.4 RegFile.scala 76:16:@130856.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@130855.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@130859.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@130853.4]
  assign regs_281_clock = clock; // @[:@130862.4]
  assign regs_281_reset = io_reset; // @[:@130863.4 RegFile.scala 76:16:@130870.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@130869.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@130873.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@130867.4]
  assign regs_282_clock = clock; // @[:@130876.4]
  assign regs_282_reset = io_reset; // @[:@130877.4 RegFile.scala 76:16:@130884.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@130883.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@130887.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@130881.4]
  assign regs_283_clock = clock; // @[:@130890.4]
  assign regs_283_reset = io_reset; // @[:@130891.4 RegFile.scala 76:16:@130898.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@130897.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@130901.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@130895.4]
  assign regs_284_clock = clock; // @[:@130904.4]
  assign regs_284_reset = io_reset; // @[:@130905.4 RegFile.scala 76:16:@130912.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@130911.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@130915.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@130909.4]
  assign regs_285_clock = clock; // @[:@130918.4]
  assign regs_285_reset = io_reset; // @[:@130919.4 RegFile.scala 76:16:@130926.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@130925.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@130929.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@130923.4]
  assign regs_286_clock = clock; // @[:@130932.4]
  assign regs_286_reset = io_reset; // @[:@130933.4 RegFile.scala 76:16:@130940.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@130939.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@130943.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@130937.4]
  assign regs_287_clock = clock; // @[:@130946.4]
  assign regs_287_reset = io_reset; // @[:@130947.4 RegFile.scala 76:16:@130954.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@130953.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@130957.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@130951.4]
  assign regs_288_clock = clock; // @[:@130960.4]
  assign regs_288_reset = io_reset; // @[:@130961.4 RegFile.scala 76:16:@130968.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@130967.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@130971.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@130965.4]
  assign regs_289_clock = clock; // @[:@130974.4]
  assign regs_289_reset = io_reset; // @[:@130975.4 RegFile.scala 76:16:@130982.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@130981.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@130985.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@130979.4]
  assign regs_290_clock = clock; // @[:@130988.4]
  assign regs_290_reset = io_reset; // @[:@130989.4 RegFile.scala 76:16:@130996.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@130995.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@130999.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@130993.4]
  assign regs_291_clock = clock; // @[:@131002.4]
  assign regs_291_reset = io_reset; // @[:@131003.4 RegFile.scala 76:16:@131010.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@131009.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@131013.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@131007.4]
  assign regs_292_clock = clock; // @[:@131016.4]
  assign regs_292_reset = io_reset; // @[:@131017.4 RegFile.scala 76:16:@131024.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@131023.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@131027.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@131021.4]
  assign regs_293_clock = clock; // @[:@131030.4]
  assign regs_293_reset = io_reset; // @[:@131031.4 RegFile.scala 76:16:@131038.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@131037.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@131041.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@131035.4]
  assign regs_294_clock = clock; // @[:@131044.4]
  assign regs_294_reset = io_reset; // @[:@131045.4 RegFile.scala 76:16:@131052.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@131051.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@131055.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@131049.4]
  assign regs_295_clock = clock; // @[:@131058.4]
  assign regs_295_reset = io_reset; // @[:@131059.4 RegFile.scala 76:16:@131066.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@131065.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@131069.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@131063.4]
  assign regs_296_clock = clock; // @[:@131072.4]
  assign regs_296_reset = io_reset; // @[:@131073.4 RegFile.scala 76:16:@131080.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@131079.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@131083.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@131077.4]
  assign regs_297_clock = clock; // @[:@131086.4]
  assign regs_297_reset = io_reset; // @[:@131087.4 RegFile.scala 76:16:@131094.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@131093.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@131097.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@131091.4]
  assign regs_298_clock = clock; // @[:@131100.4]
  assign regs_298_reset = io_reset; // @[:@131101.4 RegFile.scala 76:16:@131108.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@131107.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@131111.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@131105.4]
  assign regs_299_clock = clock; // @[:@131114.4]
  assign regs_299_reset = io_reset; // @[:@131115.4 RegFile.scala 76:16:@131122.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@131121.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@131125.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@131119.4]
  assign regs_300_clock = clock; // @[:@131128.4]
  assign regs_300_reset = io_reset; // @[:@131129.4 RegFile.scala 76:16:@131136.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@131135.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@131139.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@131133.4]
  assign regs_301_clock = clock; // @[:@131142.4]
  assign regs_301_reset = io_reset; // @[:@131143.4 RegFile.scala 76:16:@131150.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@131149.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@131153.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@131147.4]
  assign regs_302_clock = clock; // @[:@131156.4]
  assign regs_302_reset = io_reset; // @[:@131157.4 RegFile.scala 76:16:@131164.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@131163.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@131167.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@131161.4]
  assign regs_303_clock = clock; // @[:@131170.4]
  assign regs_303_reset = io_reset; // @[:@131171.4 RegFile.scala 76:16:@131178.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@131177.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@131181.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@131175.4]
  assign regs_304_clock = clock; // @[:@131184.4]
  assign regs_304_reset = io_reset; // @[:@131185.4 RegFile.scala 76:16:@131192.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@131191.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@131195.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@131189.4]
  assign regs_305_clock = clock; // @[:@131198.4]
  assign regs_305_reset = io_reset; // @[:@131199.4 RegFile.scala 76:16:@131206.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@131205.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@131209.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@131203.4]
  assign regs_306_clock = clock; // @[:@131212.4]
  assign regs_306_reset = io_reset; // @[:@131213.4 RegFile.scala 76:16:@131220.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@131219.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@131223.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@131217.4]
  assign regs_307_clock = clock; // @[:@131226.4]
  assign regs_307_reset = io_reset; // @[:@131227.4 RegFile.scala 76:16:@131234.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@131233.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@131237.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@131231.4]
  assign regs_308_clock = clock; // @[:@131240.4]
  assign regs_308_reset = io_reset; // @[:@131241.4 RegFile.scala 76:16:@131248.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@131247.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@131251.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@131245.4]
  assign regs_309_clock = clock; // @[:@131254.4]
  assign regs_309_reset = io_reset; // @[:@131255.4 RegFile.scala 76:16:@131262.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@131261.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@131265.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@131259.4]
  assign regs_310_clock = clock; // @[:@131268.4]
  assign regs_310_reset = io_reset; // @[:@131269.4 RegFile.scala 76:16:@131276.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@131275.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@131279.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@131273.4]
  assign regs_311_clock = clock; // @[:@131282.4]
  assign regs_311_reset = io_reset; // @[:@131283.4 RegFile.scala 76:16:@131290.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@131289.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@131293.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@131287.4]
  assign regs_312_clock = clock; // @[:@131296.4]
  assign regs_312_reset = io_reset; // @[:@131297.4 RegFile.scala 76:16:@131304.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@131303.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@131307.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@131301.4]
  assign regs_313_clock = clock; // @[:@131310.4]
  assign regs_313_reset = io_reset; // @[:@131311.4 RegFile.scala 76:16:@131318.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@131317.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@131321.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@131315.4]
  assign regs_314_clock = clock; // @[:@131324.4]
  assign regs_314_reset = io_reset; // @[:@131325.4 RegFile.scala 76:16:@131332.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@131331.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@131335.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@131329.4]
  assign regs_315_clock = clock; // @[:@131338.4]
  assign regs_315_reset = io_reset; // @[:@131339.4 RegFile.scala 76:16:@131346.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@131345.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@131349.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@131343.4]
  assign regs_316_clock = clock; // @[:@131352.4]
  assign regs_316_reset = io_reset; // @[:@131353.4 RegFile.scala 76:16:@131360.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@131359.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@131363.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@131357.4]
  assign regs_317_clock = clock; // @[:@131366.4]
  assign regs_317_reset = io_reset; // @[:@131367.4 RegFile.scala 76:16:@131374.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@131373.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@131377.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@131371.4]
  assign regs_318_clock = clock; // @[:@131380.4]
  assign regs_318_reset = io_reset; // @[:@131381.4 RegFile.scala 76:16:@131388.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@131387.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@131391.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@131385.4]
  assign regs_319_clock = clock; // @[:@131394.4]
  assign regs_319_reset = io_reset; // @[:@131395.4 RegFile.scala 76:16:@131402.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@131401.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@131405.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@131399.4]
  assign regs_320_clock = clock; // @[:@131408.4]
  assign regs_320_reset = io_reset; // @[:@131409.4 RegFile.scala 76:16:@131416.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@131415.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@131419.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@131413.4]
  assign regs_321_clock = clock; // @[:@131422.4]
  assign regs_321_reset = io_reset; // @[:@131423.4 RegFile.scala 76:16:@131430.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@131429.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@131433.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@131427.4]
  assign regs_322_clock = clock; // @[:@131436.4]
  assign regs_322_reset = io_reset; // @[:@131437.4 RegFile.scala 76:16:@131444.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@131443.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@131447.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@131441.4]
  assign regs_323_clock = clock; // @[:@131450.4]
  assign regs_323_reset = io_reset; // @[:@131451.4 RegFile.scala 76:16:@131458.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@131457.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@131461.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@131455.4]
  assign regs_324_clock = clock; // @[:@131464.4]
  assign regs_324_reset = io_reset; // @[:@131465.4 RegFile.scala 76:16:@131472.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@131471.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@131475.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@131469.4]
  assign regs_325_clock = clock; // @[:@131478.4]
  assign regs_325_reset = io_reset; // @[:@131479.4 RegFile.scala 76:16:@131486.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@131485.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@131489.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@131483.4]
  assign regs_326_clock = clock; // @[:@131492.4]
  assign regs_326_reset = io_reset; // @[:@131493.4 RegFile.scala 76:16:@131500.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@131499.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@131503.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@131497.4]
  assign regs_327_clock = clock; // @[:@131506.4]
  assign regs_327_reset = io_reset; // @[:@131507.4 RegFile.scala 76:16:@131514.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@131513.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@131517.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@131511.4]
  assign regs_328_clock = clock; // @[:@131520.4]
  assign regs_328_reset = io_reset; // @[:@131521.4 RegFile.scala 76:16:@131528.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@131527.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@131531.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@131525.4]
  assign regs_329_clock = clock; // @[:@131534.4]
  assign regs_329_reset = io_reset; // @[:@131535.4 RegFile.scala 76:16:@131542.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@131541.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@131545.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@131539.4]
  assign regs_330_clock = clock; // @[:@131548.4]
  assign regs_330_reset = io_reset; // @[:@131549.4 RegFile.scala 76:16:@131556.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@131555.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@131559.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@131553.4]
  assign regs_331_clock = clock; // @[:@131562.4]
  assign regs_331_reset = io_reset; // @[:@131563.4 RegFile.scala 76:16:@131570.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@131569.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@131573.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@131567.4]
  assign regs_332_clock = clock; // @[:@131576.4]
  assign regs_332_reset = io_reset; // @[:@131577.4 RegFile.scala 76:16:@131584.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@131583.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@131587.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@131581.4]
  assign regs_333_clock = clock; // @[:@131590.4]
  assign regs_333_reset = io_reset; // @[:@131591.4 RegFile.scala 76:16:@131598.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@131597.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@131601.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@131595.4]
  assign regs_334_clock = clock; // @[:@131604.4]
  assign regs_334_reset = io_reset; // @[:@131605.4 RegFile.scala 76:16:@131612.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@131611.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@131615.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@131609.4]
  assign regs_335_clock = clock; // @[:@131618.4]
  assign regs_335_reset = io_reset; // @[:@131619.4 RegFile.scala 76:16:@131626.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@131625.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@131629.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@131623.4]
  assign regs_336_clock = clock; // @[:@131632.4]
  assign regs_336_reset = io_reset; // @[:@131633.4 RegFile.scala 76:16:@131640.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@131639.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@131643.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@131637.4]
  assign regs_337_clock = clock; // @[:@131646.4]
  assign regs_337_reset = io_reset; // @[:@131647.4 RegFile.scala 76:16:@131654.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@131653.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@131657.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@131651.4]
  assign regs_338_clock = clock; // @[:@131660.4]
  assign regs_338_reset = io_reset; // @[:@131661.4 RegFile.scala 76:16:@131668.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@131667.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@131671.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@131665.4]
  assign regs_339_clock = clock; // @[:@131674.4]
  assign regs_339_reset = io_reset; // @[:@131675.4 RegFile.scala 76:16:@131682.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@131681.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@131685.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@131679.4]
  assign regs_340_clock = clock; // @[:@131688.4]
  assign regs_340_reset = io_reset; // @[:@131689.4 RegFile.scala 76:16:@131696.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@131695.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@131699.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@131693.4]
  assign regs_341_clock = clock; // @[:@131702.4]
  assign regs_341_reset = io_reset; // @[:@131703.4 RegFile.scala 76:16:@131710.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@131709.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@131713.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@131707.4]
  assign regs_342_clock = clock; // @[:@131716.4]
  assign regs_342_reset = io_reset; // @[:@131717.4 RegFile.scala 76:16:@131724.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@131723.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@131727.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@131721.4]
  assign regs_343_clock = clock; // @[:@131730.4]
  assign regs_343_reset = io_reset; // @[:@131731.4 RegFile.scala 76:16:@131738.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@131737.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@131741.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@131735.4]
  assign regs_344_clock = clock; // @[:@131744.4]
  assign regs_344_reset = io_reset; // @[:@131745.4 RegFile.scala 76:16:@131752.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@131751.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@131755.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@131749.4]
  assign regs_345_clock = clock; // @[:@131758.4]
  assign regs_345_reset = io_reset; // @[:@131759.4 RegFile.scala 76:16:@131766.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@131765.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@131769.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@131763.4]
  assign regs_346_clock = clock; // @[:@131772.4]
  assign regs_346_reset = io_reset; // @[:@131773.4 RegFile.scala 76:16:@131780.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@131779.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@131783.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@131777.4]
  assign regs_347_clock = clock; // @[:@131786.4]
  assign regs_347_reset = io_reset; // @[:@131787.4 RegFile.scala 76:16:@131794.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@131793.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@131797.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@131791.4]
  assign regs_348_clock = clock; // @[:@131800.4]
  assign regs_348_reset = io_reset; // @[:@131801.4 RegFile.scala 76:16:@131808.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@131807.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@131811.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@131805.4]
  assign regs_349_clock = clock; // @[:@131814.4]
  assign regs_349_reset = io_reset; // @[:@131815.4 RegFile.scala 76:16:@131822.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@131821.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@131825.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@131819.4]
  assign regs_350_clock = clock; // @[:@131828.4]
  assign regs_350_reset = io_reset; // @[:@131829.4 RegFile.scala 76:16:@131836.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@131835.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@131839.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@131833.4]
  assign regs_351_clock = clock; // @[:@131842.4]
  assign regs_351_reset = io_reset; // @[:@131843.4 RegFile.scala 76:16:@131850.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@131849.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@131853.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@131847.4]
  assign regs_352_clock = clock; // @[:@131856.4]
  assign regs_352_reset = io_reset; // @[:@131857.4 RegFile.scala 76:16:@131864.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@131863.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@131867.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@131861.4]
  assign regs_353_clock = clock; // @[:@131870.4]
  assign regs_353_reset = io_reset; // @[:@131871.4 RegFile.scala 76:16:@131878.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@131877.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@131881.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@131875.4]
  assign regs_354_clock = clock; // @[:@131884.4]
  assign regs_354_reset = io_reset; // @[:@131885.4 RegFile.scala 76:16:@131892.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@131891.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@131895.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@131889.4]
  assign regs_355_clock = clock; // @[:@131898.4]
  assign regs_355_reset = io_reset; // @[:@131899.4 RegFile.scala 76:16:@131906.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@131905.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@131909.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@131903.4]
  assign regs_356_clock = clock; // @[:@131912.4]
  assign regs_356_reset = io_reset; // @[:@131913.4 RegFile.scala 76:16:@131920.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@131919.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@131923.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@131917.4]
  assign regs_357_clock = clock; // @[:@131926.4]
  assign regs_357_reset = io_reset; // @[:@131927.4 RegFile.scala 76:16:@131934.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@131933.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@131937.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@131931.4]
  assign regs_358_clock = clock; // @[:@131940.4]
  assign regs_358_reset = io_reset; // @[:@131941.4 RegFile.scala 76:16:@131948.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@131947.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@131951.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@131945.4]
  assign regs_359_clock = clock; // @[:@131954.4]
  assign regs_359_reset = io_reset; // @[:@131955.4 RegFile.scala 76:16:@131962.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@131961.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@131965.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@131959.4]
  assign regs_360_clock = clock; // @[:@131968.4]
  assign regs_360_reset = io_reset; // @[:@131969.4 RegFile.scala 76:16:@131976.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@131975.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@131979.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@131973.4]
  assign regs_361_clock = clock; // @[:@131982.4]
  assign regs_361_reset = io_reset; // @[:@131983.4 RegFile.scala 76:16:@131990.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@131989.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@131993.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@131987.4]
  assign regs_362_clock = clock; // @[:@131996.4]
  assign regs_362_reset = io_reset; // @[:@131997.4 RegFile.scala 76:16:@132004.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@132003.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@132007.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@132001.4]
  assign regs_363_clock = clock; // @[:@132010.4]
  assign regs_363_reset = io_reset; // @[:@132011.4 RegFile.scala 76:16:@132018.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@132017.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@132021.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@132015.4]
  assign regs_364_clock = clock; // @[:@132024.4]
  assign regs_364_reset = io_reset; // @[:@132025.4 RegFile.scala 76:16:@132032.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@132031.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@132035.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@132029.4]
  assign regs_365_clock = clock; // @[:@132038.4]
  assign regs_365_reset = io_reset; // @[:@132039.4 RegFile.scala 76:16:@132046.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@132045.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@132049.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@132043.4]
  assign regs_366_clock = clock; // @[:@132052.4]
  assign regs_366_reset = io_reset; // @[:@132053.4 RegFile.scala 76:16:@132060.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@132059.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@132063.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@132057.4]
  assign regs_367_clock = clock; // @[:@132066.4]
  assign regs_367_reset = io_reset; // @[:@132067.4 RegFile.scala 76:16:@132074.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@132073.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@132077.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@132071.4]
  assign regs_368_clock = clock; // @[:@132080.4]
  assign regs_368_reset = io_reset; // @[:@132081.4 RegFile.scala 76:16:@132088.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@132087.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@132091.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@132085.4]
  assign regs_369_clock = clock; // @[:@132094.4]
  assign regs_369_reset = io_reset; // @[:@132095.4 RegFile.scala 76:16:@132102.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@132101.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@132105.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@132099.4]
  assign regs_370_clock = clock; // @[:@132108.4]
  assign regs_370_reset = io_reset; // @[:@132109.4 RegFile.scala 76:16:@132116.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@132115.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@132119.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@132113.4]
  assign regs_371_clock = clock; // @[:@132122.4]
  assign regs_371_reset = io_reset; // @[:@132123.4 RegFile.scala 76:16:@132130.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@132129.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@132133.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@132127.4]
  assign regs_372_clock = clock; // @[:@132136.4]
  assign regs_372_reset = io_reset; // @[:@132137.4 RegFile.scala 76:16:@132144.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@132143.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@132147.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@132141.4]
  assign regs_373_clock = clock; // @[:@132150.4]
  assign regs_373_reset = io_reset; // @[:@132151.4 RegFile.scala 76:16:@132158.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@132157.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@132161.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@132155.4]
  assign regs_374_clock = clock; // @[:@132164.4]
  assign regs_374_reset = io_reset; // @[:@132165.4 RegFile.scala 76:16:@132172.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@132171.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@132175.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@132169.4]
  assign regs_375_clock = clock; // @[:@132178.4]
  assign regs_375_reset = io_reset; // @[:@132179.4 RegFile.scala 76:16:@132186.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@132185.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@132189.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@132183.4]
  assign regs_376_clock = clock; // @[:@132192.4]
  assign regs_376_reset = io_reset; // @[:@132193.4 RegFile.scala 76:16:@132200.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@132199.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@132203.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@132197.4]
  assign regs_377_clock = clock; // @[:@132206.4]
  assign regs_377_reset = io_reset; // @[:@132207.4 RegFile.scala 76:16:@132214.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@132213.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@132217.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@132211.4]
  assign regs_378_clock = clock; // @[:@132220.4]
  assign regs_378_reset = io_reset; // @[:@132221.4 RegFile.scala 76:16:@132228.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@132227.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@132231.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@132225.4]
  assign regs_379_clock = clock; // @[:@132234.4]
  assign regs_379_reset = io_reset; // @[:@132235.4 RegFile.scala 76:16:@132242.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@132241.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@132245.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@132239.4]
  assign regs_380_clock = clock; // @[:@132248.4]
  assign regs_380_reset = io_reset; // @[:@132249.4 RegFile.scala 76:16:@132256.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@132255.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@132259.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@132253.4]
  assign regs_381_clock = clock; // @[:@132262.4]
  assign regs_381_reset = io_reset; // @[:@132263.4 RegFile.scala 76:16:@132270.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@132269.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@132273.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@132267.4]
  assign regs_382_clock = clock; // @[:@132276.4]
  assign regs_382_reset = io_reset; // @[:@132277.4 RegFile.scala 76:16:@132284.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@132283.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@132287.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@132281.4]
  assign regs_383_clock = clock; // @[:@132290.4]
  assign regs_383_reset = io_reset; // @[:@132291.4 RegFile.scala 76:16:@132298.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@132297.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@132301.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@132295.4]
  assign regs_384_clock = clock; // @[:@132304.4]
  assign regs_384_reset = io_reset; // @[:@132305.4 RegFile.scala 76:16:@132312.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@132311.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@132315.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@132309.4]
  assign regs_385_clock = clock; // @[:@132318.4]
  assign regs_385_reset = io_reset; // @[:@132319.4 RegFile.scala 76:16:@132326.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@132325.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@132329.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@132323.4]
  assign regs_386_clock = clock; // @[:@132332.4]
  assign regs_386_reset = io_reset; // @[:@132333.4 RegFile.scala 76:16:@132340.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@132339.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@132343.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@132337.4]
  assign regs_387_clock = clock; // @[:@132346.4]
  assign regs_387_reset = io_reset; // @[:@132347.4 RegFile.scala 76:16:@132354.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@132353.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@132357.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@132351.4]
  assign regs_388_clock = clock; // @[:@132360.4]
  assign regs_388_reset = io_reset; // @[:@132361.4 RegFile.scala 76:16:@132368.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@132367.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@132371.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@132365.4]
  assign regs_389_clock = clock; // @[:@132374.4]
  assign regs_389_reset = io_reset; // @[:@132375.4 RegFile.scala 76:16:@132382.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@132381.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@132385.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@132379.4]
  assign regs_390_clock = clock; // @[:@132388.4]
  assign regs_390_reset = io_reset; // @[:@132389.4 RegFile.scala 76:16:@132396.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@132395.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@132399.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@132393.4]
  assign regs_391_clock = clock; // @[:@132402.4]
  assign regs_391_reset = io_reset; // @[:@132403.4 RegFile.scala 76:16:@132410.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@132409.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@132413.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@132407.4]
  assign regs_392_clock = clock; // @[:@132416.4]
  assign regs_392_reset = io_reset; // @[:@132417.4 RegFile.scala 76:16:@132424.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@132423.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@132427.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@132421.4]
  assign regs_393_clock = clock; // @[:@132430.4]
  assign regs_393_reset = io_reset; // @[:@132431.4 RegFile.scala 76:16:@132438.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@132437.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@132441.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@132435.4]
  assign regs_394_clock = clock; // @[:@132444.4]
  assign regs_394_reset = io_reset; // @[:@132445.4 RegFile.scala 76:16:@132452.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@132451.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@132455.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@132449.4]
  assign regs_395_clock = clock; // @[:@132458.4]
  assign regs_395_reset = io_reset; // @[:@132459.4 RegFile.scala 76:16:@132466.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@132465.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@132469.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@132463.4]
  assign regs_396_clock = clock; // @[:@132472.4]
  assign regs_396_reset = io_reset; // @[:@132473.4 RegFile.scala 76:16:@132480.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@132479.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@132483.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@132477.4]
  assign regs_397_clock = clock; // @[:@132486.4]
  assign regs_397_reset = io_reset; // @[:@132487.4 RegFile.scala 76:16:@132494.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@132493.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@132497.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@132491.4]
  assign regs_398_clock = clock; // @[:@132500.4]
  assign regs_398_reset = io_reset; // @[:@132501.4 RegFile.scala 76:16:@132508.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@132507.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@132511.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@132505.4]
  assign regs_399_clock = clock; // @[:@132514.4]
  assign regs_399_reset = io_reset; // @[:@132515.4 RegFile.scala 76:16:@132522.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@132521.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@132525.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@132519.4]
  assign regs_400_clock = clock; // @[:@132528.4]
  assign regs_400_reset = io_reset; // @[:@132529.4 RegFile.scala 76:16:@132536.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@132535.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@132539.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@132533.4]
  assign regs_401_clock = clock; // @[:@132542.4]
  assign regs_401_reset = io_reset; // @[:@132543.4 RegFile.scala 76:16:@132550.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@132549.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@132553.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@132547.4]
  assign regs_402_clock = clock; // @[:@132556.4]
  assign regs_402_reset = io_reset; // @[:@132557.4 RegFile.scala 76:16:@132564.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@132563.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@132567.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@132561.4]
  assign regs_403_clock = clock; // @[:@132570.4]
  assign regs_403_reset = io_reset; // @[:@132571.4 RegFile.scala 76:16:@132578.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@132577.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@132581.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@132575.4]
  assign regs_404_clock = clock; // @[:@132584.4]
  assign regs_404_reset = io_reset; // @[:@132585.4 RegFile.scala 76:16:@132592.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@132591.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@132595.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@132589.4]
  assign regs_405_clock = clock; // @[:@132598.4]
  assign regs_405_reset = io_reset; // @[:@132599.4 RegFile.scala 76:16:@132606.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@132605.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@132609.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@132603.4]
  assign regs_406_clock = clock; // @[:@132612.4]
  assign regs_406_reset = io_reset; // @[:@132613.4 RegFile.scala 76:16:@132620.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@132619.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@132623.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@132617.4]
  assign regs_407_clock = clock; // @[:@132626.4]
  assign regs_407_reset = io_reset; // @[:@132627.4 RegFile.scala 76:16:@132634.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@132633.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@132637.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@132631.4]
  assign regs_408_clock = clock; // @[:@132640.4]
  assign regs_408_reset = io_reset; // @[:@132641.4 RegFile.scala 76:16:@132648.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@132647.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@132651.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@132645.4]
  assign regs_409_clock = clock; // @[:@132654.4]
  assign regs_409_reset = io_reset; // @[:@132655.4 RegFile.scala 76:16:@132662.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@132661.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@132665.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@132659.4]
  assign regs_410_clock = clock; // @[:@132668.4]
  assign regs_410_reset = io_reset; // @[:@132669.4 RegFile.scala 76:16:@132676.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@132675.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@132679.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@132673.4]
  assign regs_411_clock = clock; // @[:@132682.4]
  assign regs_411_reset = io_reset; // @[:@132683.4 RegFile.scala 76:16:@132690.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@132689.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@132693.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@132687.4]
  assign regs_412_clock = clock; // @[:@132696.4]
  assign regs_412_reset = io_reset; // @[:@132697.4 RegFile.scala 76:16:@132704.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@132703.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@132707.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@132701.4]
  assign regs_413_clock = clock; // @[:@132710.4]
  assign regs_413_reset = io_reset; // @[:@132711.4 RegFile.scala 76:16:@132718.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@132717.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@132721.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@132715.4]
  assign regs_414_clock = clock; // @[:@132724.4]
  assign regs_414_reset = io_reset; // @[:@132725.4 RegFile.scala 76:16:@132732.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@132731.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@132735.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@132729.4]
  assign regs_415_clock = clock; // @[:@132738.4]
  assign regs_415_reset = io_reset; // @[:@132739.4 RegFile.scala 76:16:@132746.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@132745.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@132749.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@132743.4]
  assign regs_416_clock = clock; // @[:@132752.4]
  assign regs_416_reset = io_reset; // @[:@132753.4 RegFile.scala 76:16:@132760.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@132759.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@132763.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@132757.4]
  assign regs_417_clock = clock; // @[:@132766.4]
  assign regs_417_reset = io_reset; // @[:@132767.4 RegFile.scala 76:16:@132774.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@132773.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@132777.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@132771.4]
  assign regs_418_clock = clock; // @[:@132780.4]
  assign regs_418_reset = io_reset; // @[:@132781.4 RegFile.scala 76:16:@132788.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@132787.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@132791.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@132785.4]
  assign regs_419_clock = clock; // @[:@132794.4]
  assign regs_419_reset = io_reset; // @[:@132795.4 RegFile.scala 76:16:@132802.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@132801.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@132805.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@132799.4]
  assign regs_420_clock = clock; // @[:@132808.4]
  assign regs_420_reset = io_reset; // @[:@132809.4 RegFile.scala 76:16:@132816.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@132815.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@132819.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@132813.4]
  assign regs_421_clock = clock; // @[:@132822.4]
  assign regs_421_reset = io_reset; // @[:@132823.4 RegFile.scala 76:16:@132830.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@132829.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@132833.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@132827.4]
  assign regs_422_clock = clock; // @[:@132836.4]
  assign regs_422_reset = io_reset; // @[:@132837.4 RegFile.scala 76:16:@132844.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@132843.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@132847.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@132841.4]
  assign regs_423_clock = clock; // @[:@132850.4]
  assign regs_423_reset = io_reset; // @[:@132851.4 RegFile.scala 76:16:@132858.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@132857.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@132861.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@132855.4]
  assign regs_424_clock = clock; // @[:@132864.4]
  assign regs_424_reset = io_reset; // @[:@132865.4 RegFile.scala 76:16:@132872.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@132871.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@132875.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@132869.4]
  assign regs_425_clock = clock; // @[:@132878.4]
  assign regs_425_reset = io_reset; // @[:@132879.4 RegFile.scala 76:16:@132886.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@132885.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@132889.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@132883.4]
  assign regs_426_clock = clock; // @[:@132892.4]
  assign regs_426_reset = io_reset; // @[:@132893.4 RegFile.scala 76:16:@132900.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@132899.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@132903.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@132897.4]
  assign regs_427_clock = clock; // @[:@132906.4]
  assign regs_427_reset = io_reset; // @[:@132907.4 RegFile.scala 76:16:@132914.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@132913.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@132917.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@132911.4]
  assign regs_428_clock = clock; // @[:@132920.4]
  assign regs_428_reset = io_reset; // @[:@132921.4 RegFile.scala 76:16:@132928.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@132927.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@132931.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@132925.4]
  assign regs_429_clock = clock; // @[:@132934.4]
  assign regs_429_reset = io_reset; // @[:@132935.4 RegFile.scala 76:16:@132942.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@132941.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@132945.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@132939.4]
  assign regs_430_clock = clock; // @[:@132948.4]
  assign regs_430_reset = io_reset; // @[:@132949.4 RegFile.scala 76:16:@132956.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@132955.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@132959.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@132953.4]
  assign regs_431_clock = clock; // @[:@132962.4]
  assign regs_431_reset = io_reset; // @[:@132963.4 RegFile.scala 76:16:@132970.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@132969.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@132973.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@132967.4]
  assign regs_432_clock = clock; // @[:@132976.4]
  assign regs_432_reset = io_reset; // @[:@132977.4 RegFile.scala 76:16:@132984.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@132983.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@132987.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@132981.4]
  assign regs_433_clock = clock; // @[:@132990.4]
  assign regs_433_reset = io_reset; // @[:@132991.4 RegFile.scala 76:16:@132998.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@132997.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@133001.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@132995.4]
  assign regs_434_clock = clock; // @[:@133004.4]
  assign regs_434_reset = io_reset; // @[:@133005.4 RegFile.scala 76:16:@133012.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@133011.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@133015.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@133009.4]
  assign regs_435_clock = clock; // @[:@133018.4]
  assign regs_435_reset = io_reset; // @[:@133019.4 RegFile.scala 76:16:@133026.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@133025.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@133029.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@133023.4]
  assign regs_436_clock = clock; // @[:@133032.4]
  assign regs_436_reset = io_reset; // @[:@133033.4 RegFile.scala 76:16:@133040.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@133039.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@133043.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@133037.4]
  assign regs_437_clock = clock; // @[:@133046.4]
  assign regs_437_reset = io_reset; // @[:@133047.4 RegFile.scala 76:16:@133054.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@133053.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@133057.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@133051.4]
  assign regs_438_clock = clock; // @[:@133060.4]
  assign regs_438_reset = io_reset; // @[:@133061.4 RegFile.scala 76:16:@133068.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@133067.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@133071.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@133065.4]
  assign regs_439_clock = clock; // @[:@133074.4]
  assign regs_439_reset = io_reset; // @[:@133075.4 RegFile.scala 76:16:@133082.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@133081.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@133085.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@133079.4]
  assign regs_440_clock = clock; // @[:@133088.4]
  assign regs_440_reset = io_reset; // @[:@133089.4 RegFile.scala 76:16:@133096.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@133095.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@133099.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@133093.4]
  assign regs_441_clock = clock; // @[:@133102.4]
  assign regs_441_reset = io_reset; // @[:@133103.4 RegFile.scala 76:16:@133110.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@133109.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@133113.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@133107.4]
  assign regs_442_clock = clock; // @[:@133116.4]
  assign regs_442_reset = io_reset; // @[:@133117.4 RegFile.scala 76:16:@133124.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@133123.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@133127.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@133121.4]
  assign regs_443_clock = clock; // @[:@133130.4]
  assign regs_443_reset = io_reset; // @[:@133131.4 RegFile.scala 76:16:@133138.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@133137.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@133141.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@133135.4]
  assign regs_444_clock = clock; // @[:@133144.4]
  assign regs_444_reset = io_reset; // @[:@133145.4 RegFile.scala 76:16:@133152.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@133151.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@133155.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@133149.4]
  assign regs_445_clock = clock; // @[:@133158.4]
  assign regs_445_reset = io_reset; // @[:@133159.4 RegFile.scala 76:16:@133166.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@133165.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@133169.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@133163.4]
  assign regs_446_clock = clock; // @[:@133172.4]
  assign regs_446_reset = io_reset; // @[:@133173.4 RegFile.scala 76:16:@133180.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@133179.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@133183.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@133177.4]
  assign regs_447_clock = clock; // @[:@133186.4]
  assign regs_447_reset = io_reset; // @[:@133187.4 RegFile.scala 76:16:@133194.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@133193.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@133197.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@133191.4]
  assign regs_448_clock = clock; // @[:@133200.4]
  assign regs_448_reset = io_reset; // @[:@133201.4 RegFile.scala 76:16:@133208.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@133207.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@133211.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@133205.4]
  assign regs_449_clock = clock; // @[:@133214.4]
  assign regs_449_reset = io_reset; // @[:@133215.4 RegFile.scala 76:16:@133222.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@133221.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@133225.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@133219.4]
  assign regs_450_clock = clock; // @[:@133228.4]
  assign regs_450_reset = io_reset; // @[:@133229.4 RegFile.scala 76:16:@133236.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@133235.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@133239.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@133233.4]
  assign regs_451_clock = clock; // @[:@133242.4]
  assign regs_451_reset = io_reset; // @[:@133243.4 RegFile.scala 76:16:@133250.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@133249.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@133253.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@133247.4]
  assign regs_452_clock = clock; // @[:@133256.4]
  assign regs_452_reset = io_reset; // @[:@133257.4 RegFile.scala 76:16:@133264.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@133263.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@133267.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@133261.4]
  assign regs_453_clock = clock; // @[:@133270.4]
  assign regs_453_reset = io_reset; // @[:@133271.4 RegFile.scala 76:16:@133278.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@133277.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@133281.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@133275.4]
  assign regs_454_clock = clock; // @[:@133284.4]
  assign regs_454_reset = io_reset; // @[:@133285.4 RegFile.scala 76:16:@133292.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@133291.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@133295.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@133289.4]
  assign regs_455_clock = clock; // @[:@133298.4]
  assign regs_455_reset = io_reset; // @[:@133299.4 RegFile.scala 76:16:@133306.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@133305.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@133309.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@133303.4]
  assign regs_456_clock = clock; // @[:@133312.4]
  assign regs_456_reset = io_reset; // @[:@133313.4 RegFile.scala 76:16:@133320.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@133319.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@133323.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@133317.4]
  assign regs_457_clock = clock; // @[:@133326.4]
  assign regs_457_reset = io_reset; // @[:@133327.4 RegFile.scala 76:16:@133334.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@133333.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@133337.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@133331.4]
  assign regs_458_clock = clock; // @[:@133340.4]
  assign regs_458_reset = io_reset; // @[:@133341.4 RegFile.scala 76:16:@133348.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@133347.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@133351.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@133345.4]
  assign regs_459_clock = clock; // @[:@133354.4]
  assign regs_459_reset = io_reset; // @[:@133355.4 RegFile.scala 76:16:@133362.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@133361.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@133365.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@133359.4]
  assign regs_460_clock = clock; // @[:@133368.4]
  assign regs_460_reset = io_reset; // @[:@133369.4 RegFile.scala 76:16:@133376.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@133375.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@133379.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@133373.4]
  assign regs_461_clock = clock; // @[:@133382.4]
  assign regs_461_reset = io_reset; // @[:@133383.4 RegFile.scala 76:16:@133390.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@133389.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@133393.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@133387.4]
  assign regs_462_clock = clock; // @[:@133396.4]
  assign regs_462_reset = io_reset; // @[:@133397.4 RegFile.scala 76:16:@133404.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@133403.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@133407.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@133401.4]
  assign regs_463_clock = clock; // @[:@133410.4]
  assign regs_463_reset = io_reset; // @[:@133411.4 RegFile.scala 76:16:@133418.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@133417.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@133421.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@133415.4]
  assign regs_464_clock = clock; // @[:@133424.4]
  assign regs_464_reset = io_reset; // @[:@133425.4 RegFile.scala 76:16:@133432.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@133431.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@133435.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@133429.4]
  assign regs_465_clock = clock; // @[:@133438.4]
  assign regs_465_reset = io_reset; // @[:@133439.4 RegFile.scala 76:16:@133446.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@133445.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@133449.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@133443.4]
  assign regs_466_clock = clock; // @[:@133452.4]
  assign regs_466_reset = io_reset; // @[:@133453.4 RegFile.scala 76:16:@133460.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@133459.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@133463.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@133457.4]
  assign regs_467_clock = clock; // @[:@133466.4]
  assign regs_467_reset = io_reset; // @[:@133467.4 RegFile.scala 76:16:@133474.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@133473.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@133477.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@133471.4]
  assign regs_468_clock = clock; // @[:@133480.4]
  assign regs_468_reset = io_reset; // @[:@133481.4 RegFile.scala 76:16:@133488.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@133487.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@133491.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@133485.4]
  assign regs_469_clock = clock; // @[:@133494.4]
  assign regs_469_reset = io_reset; // @[:@133495.4 RegFile.scala 76:16:@133502.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@133501.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@133505.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@133499.4]
  assign regs_470_clock = clock; // @[:@133508.4]
  assign regs_470_reset = io_reset; // @[:@133509.4 RegFile.scala 76:16:@133516.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@133515.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@133519.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@133513.4]
  assign regs_471_clock = clock; // @[:@133522.4]
  assign regs_471_reset = io_reset; // @[:@133523.4 RegFile.scala 76:16:@133530.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@133529.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@133533.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@133527.4]
  assign regs_472_clock = clock; // @[:@133536.4]
  assign regs_472_reset = io_reset; // @[:@133537.4 RegFile.scala 76:16:@133544.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@133543.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@133547.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@133541.4]
  assign regs_473_clock = clock; // @[:@133550.4]
  assign regs_473_reset = io_reset; // @[:@133551.4 RegFile.scala 76:16:@133558.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@133557.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@133561.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@133555.4]
  assign regs_474_clock = clock; // @[:@133564.4]
  assign regs_474_reset = io_reset; // @[:@133565.4 RegFile.scala 76:16:@133572.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@133571.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@133575.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@133569.4]
  assign regs_475_clock = clock; // @[:@133578.4]
  assign regs_475_reset = io_reset; // @[:@133579.4 RegFile.scala 76:16:@133586.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@133585.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@133589.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@133583.4]
  assign regs_476_clock = clock; // @[:@133592.4]
  assign regs_476_reset = io_reset; // @[:@133593.4 RegFile.scala 76:16:@133600.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@133599.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@133603.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@133597.4]
  assign regs_477_clock = clock; // @[:@133606.4]
  assign regs_477_reset = io_reset; // @[:@133607.4 RegFile.scala 76:16:@133614.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@133613.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@133617.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@133611.4]
  assign regs_478_clock = clock; // @[:@133620.4]
  assign regs_478_reset = io_reset; // @[:@133621.4 RegFile.scala 76:16:@133628.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@133627.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@133631.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@133625.4]
  assign regs_479_clock = clock; // @[:@133634.4]
  assign regs_479_reset = io_reset; // @[:@133635.4 RegFile.scala 76:16:@133642.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@133641.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@133645.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@133639.4]
  assign regs_480_clock = clock; // @[:@133648.4]
  assign regs_480_reset = io_reset; // @[:@133649.4 RegFile.scala 76:16:@133656.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@133655.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@133659.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@133653.4]
  assign regs_481_clock = clock; // @[:@133662.4]
  assign regs_481_reset = io_reset; // @[:@133663.4 RegFile.scala 76:16:@133670.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@133669.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@133673.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@133667.4]
  assign regs_482_clock = clock; // @[:@133676.4]
  assign regs_482_reset = io_reset; // @[:@133677.4 RegFile.scala 76:16:@133684.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@133683.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@133687.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@133681.4]
  assign regs_483_clock = clock; // @[:@133690.4]
  assign regs_483_reset = io_reset; // @[:@133691.4 RegFile.scala 76:16:@133698.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@133697.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@133701.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@133695.4]
  assign regs_484_clock = clock; // @[:@133704.4]
  assign regs_484_reset = io_reset; // @[:@133705.4 RegFile.scala 76:16:@133712.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@133711.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@133715.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@133709.4]
  assign regs_485_clock = clock; // @[:@133718.4]
  assign regs_485_reset = io_reset; // @[:@133719.4 RegFile.scala 76:16:@133726.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@133725.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@133729.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@133723.4]
  assign regs_486_clock = clock; // @[:@133732.4]
  assign regs_486_reset = io_reset; // @[:@133733.4 RegFile.scala 76:16:@133740.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@133739.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@133743.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@133737.4]
  assign regs_487_clock = clock; // @[:@133746.4]
  assign regs_487_reset = io_reset; // @[:@133747.4 RegFile.scala 76:16:@133754.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@133753.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@133757.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@133751.4]
  assign regs_488_clock = clock; // @[:@133760.4]
  assign regs_488_reset = io_reset; // @[:@133761.4 RegFile.scala 76:16:@133768.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@133767.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@133771.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@133765.4]
  assign regs_489_clock = clock; // @[:@133774.4]
  assign regs_489_reset = io_reset; // @[:@133775.4 RegFile.scala 76:16:@133782.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@133781.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@133785.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@133779.4]
  assign regs_490_clock = clock; // @[:@133788.4]
  assign regs_490_reset = io_reset; // @[:@133789.4 RegFile.scala 76:16:@133796.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@133795.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@133799.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@133793.4]
  assign regs_491_clock = clock; // @[:@133802.4]
  assign regs_491_reset = io_reset; // @[:@133803.4 RegFile.scala 76:16:@133810.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@133809.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@133813.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@133807.4]
  assign regs_492_clock = clock; // @[:@133816.4]
  assign regs_492_reset = io_reset; // @[:@133817.4 RegFile.scala 76:16:@133824.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@133823.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@133827.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@133821.4]
  assign regs_493_clock = clock; // @[:@133830.4]
  assign regs_493_reset = io_reset; // @[:@133831.4 RegFile.scala 76:16:@133838.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@133837.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@133841.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@133835.4]
  assign regs_494_clock = clock; // @[:@133844.4]
  assign regs_494_reset = io_reset; // @[:@133845.4 RegFile.scala 76:16:@133852.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@133851.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@133855.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@133849.4]
  assign regs_495_clock = clock; // @[:@133858.4]
  assign regs_495_reset = io_reset; // @[:@133859.4 RegFile.scala 76:16:@133866.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@133865.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@133869.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@133863.4]
  assign regs_496_clock = clock; // @[:@133872.4]
  assign regs_496_reset = io_reset; // @[:@133873.4 RegFile.scala 76:16:@133880.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@133879.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@133883.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@133877.4]
  assign regs_497_clock = clock; // @[:@133886.4]
  assign regs_497_reset = io_reset; // @[:@133887.4 RegFile.scala 76:16:@133894.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@133893.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@133897.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@133891.4]
  assign regs_498_clock = clock; // @[:@133900.4]
  assign regs_498_reset = io_reset; // @[:@133901.4 RegFile.scala 76:16:@133908.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@133907.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@133911.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@133905.4]
  assign regs_499_clock = clock; // @[:@133914.4]
  assign regs_499_reset = io_reset; // @[:@133915.4 RegFile.scala 76:16:@133922.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@133921.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@133925.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@133919.4]
  assign regs_500_clock = clock; // @[:@133928.4]
  assign regs_500_reset = io_reset; // @[:@133929.4 RegFile.scala 76:16:@133936.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@133935.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@133939.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@133933.4]
  assign regs_501_clock = clock; // @[:@133942.4]
  assign regs_501_reset = io_reset; // @[:@133943.4 RegFile.scala 76:16:@133950.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@133949.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@133953.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@133947.4]
  assign regs_502_clock = clock; // @[:@133956.4]
  assign regs_502_reset = io_reset; // @[:@133957.4 RegFile.scala 76:16:@133964.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@133963.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@133967.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@133961.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@134476.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@134477.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@134478.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@134479.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@134480.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@134481.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@134482.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@134483.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@134484.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@134485.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@134486.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@134487.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@134488.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@134489.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@134490.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@134491.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@134492.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@134493.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@134494.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@134495.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@134496.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@134497.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@134498.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@134499.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@134500.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@134501.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@134502.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@134503.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@134504.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@134505.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@134506.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@134507.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@134508.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@134509.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@134510.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@134511.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@134512.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@134513.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@134514.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@134515.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@134516.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@134517.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@134518.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@134519.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@134520.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@134521.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@134522.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@134523.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@134524.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@134525.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@134526.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@134527.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@134528.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@134529.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@134530.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@134531.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@134532.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@134533.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@134534.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@134535.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@134536.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@134537.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@134538.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@134539.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@134540.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@134541.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@134542.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@134543.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@134544.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@134545.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@134546.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@134547.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@134548.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@134549.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@134550.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@134551.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@134552.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@134553.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@134554.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@134555.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@134556.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@134557.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@134558.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@134559.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@134560.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@134561.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@134562.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@134563.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@134564.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@134565.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@134566.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@134567.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@134568.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@134569.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@134570.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@134571.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@134572.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@134573.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@134574.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@134575.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@134576.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@134577.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@134578.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@134579.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@134580.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@134581.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@134582.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@134583.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@134584.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@134585.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@134586.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@134587.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@134588.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@134589.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@134590.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@134591.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@134592.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@134593.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@134594.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@134595.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@134596.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@134597.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@134598.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@134599.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@134600.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@134601.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@134602.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@134603.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@134604.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@134605.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@134606.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@134607.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@134608.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@134609.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@134610.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@134611.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@134612.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@134613.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@134614.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@134615.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@134616.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@134617.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@134618.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@134619.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@134620.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@134621.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@134622.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@134623.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@134624.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@134625.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@134626.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@134627.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@134628.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@134629.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@134630.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@134631.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@134632.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@134633.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@134634.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@134635.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@134636.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@134637.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@134638.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@134639.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@134640.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@134641.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@134642.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@134643.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@134644.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@134645.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@134646.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@134647.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@134648.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@134649.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@134650.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@134651.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@134652.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@134653.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@134654.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@134655.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@134656.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@134657.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@134658.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@134659.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@134660.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@134661.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@134662.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@134663.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@134664.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@134665.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@134666.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@134667.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@134668.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@134669.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@134670.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@134671.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@134672.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@134673.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@134674.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@134675.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@134676.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@134677.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@134678.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@134679.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@134680.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@134681.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@134682.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@134683.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@134684.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@134685.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@134686.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@134687.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@134688.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@134689.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@134690.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@134691.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@134692.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@134693.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@134694.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@134695.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@134696.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@134697.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@134698.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@134699.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@134700.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@134701.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@134702.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@134703.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@134704.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@134705.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@134706.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@134707.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@134708.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@134709.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@134710.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@134711.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@134712.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@134713.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@134714.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@134715.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@134716.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@134717.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@134718.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@134719.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@134720.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@134721.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@134722.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@134723.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@134724.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@134725.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@134726.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@134727.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@134728.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@134729.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@134730.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@134731.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@134732.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@134733.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@134734.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@134735.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@134736.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@134737.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@134738.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@134739.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@134740.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@134741.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@134742.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@134743.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@134744.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@134745.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@134746.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@134747.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@134748.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@134749.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@134750.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@134751.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@134752.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@134753.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@134754.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@134755.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@134756.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@134757.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@134758.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@134759.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@134760.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@134761.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@134762.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@134763.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@134764.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@134765.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@134766.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@134767.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@134768.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@134769.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@134770.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@134771.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@134772.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@134773.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@134774.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@134775.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@134776.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@134777.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@134778.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@134779.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@134780.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@134781.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@134782.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@134783.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@134784.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@134785.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@134786.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@134787.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@134788.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@134789.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@134790.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@134791.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@134792.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@134793.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@134794.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@134795.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@134796.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@134797.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@134798.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@134799.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@134800.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@134801.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@134802.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@134803.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@134804.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@134805.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@134806.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@134807.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@134808.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@134809.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@134810.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@134811.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@134812.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@134813.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@134814.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@134815.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@134816.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@134817.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@134818.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@134819.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@134820.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@134821.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@134822.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@134823.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@134824.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@134825.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@134826.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@134827.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@134828.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@134829.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@134830.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@134831.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@134832.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@134833.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@134834.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@134835.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@134836.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@134837.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@134838.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@134839.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@134840.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@134841.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@134842.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@134843.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@134844.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@134845.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@134846.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@134847.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@134848.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@134849.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@134850.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@134851.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@134852.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@134853.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@134854.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@134855.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@134856.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@134857.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@134858.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@134859.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@134860.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@134861.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@134862.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@134863.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@134864.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@134865.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@134866.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@134867.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@134868.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@134869.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@134870.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@134871.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@134872.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@134873.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@134874.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@134875.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@134876.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@134877.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@134878.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@134879.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@134880.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@134881.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@134882.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@134883.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@134884.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@134885.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@134886.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@134887.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@134888.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@134889.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@134890.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@134891.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@134892.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@134893.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@134894.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@134895.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@134896.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@134897.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@134898.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@134899.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@134900.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@134901.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@134902.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@134903.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@134904.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@134905.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@134906.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@134907.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@134908.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@134909.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@134910.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@134911.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@134912.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@134913.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@134914.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@134915.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@134916.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@134917.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@134918.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@134919.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@134920.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@134921.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@134922.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@134923.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@134924.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@134925.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@134926.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@134927.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@134928.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@134929.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@134930.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@134931.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@134932.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@134933.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@134934.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@134935.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@134936.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@134937.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@134938.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@134939.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@134940.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@134941.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@134942.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@134943.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@134944.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@134945.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@134946.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@134947.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@134948.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@134949.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@134950.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@134951.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@134952.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@134953.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@134954.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@134955.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@134956.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@134957.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@134958.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@134959.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@134960.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@134961.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@134962.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@134963.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@134964.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@134965.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@134966.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@134967.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@134968.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@134969.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@134970.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@134971.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@134972.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@134973.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@134974.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@134975.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@134976.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@134977.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@134978.4]
  assign rport_io_sel = io_raddr[8:0]; // @[RegFile.scala 106:18:@134979.4]
endmodule
module RetimeWrapper_836( // @[:@135003.2]
  input         clock, // @[:@135004.4]
  input         reset, // @[:@135005.4]
  input  [39:0] io_in, // @[:@135006.4]
  output [39:0] io_out // @[:@135006.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@135008.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@135008.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@135008.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@135008.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@135008.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@135008.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@135008.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@135021.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@135020.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@135019.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@135018.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@135017.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@135015.4]
endmodule
module FringeFF_503( // @[:@135023.2]
  input         clock, // @[:@135024.4]
  input         reset, // @[:@135025.4]
  input  [39:0] io_in, // @[:@135026.4]
  output [39:0] io_out, // @[:@135026.4]
  input         io_enable // @[:@135026.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@135029.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@135029.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@135029.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@135029.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@135034.4 package.scala 96:25:@135035.4]
  RetimeWrapper_836 RetimeWrapper ( // @[package.scala 93:22:@135029.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@135034.4 package.scala 96:25:@135035.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@135046.4]
  assign RetimeWrapper_clock = clock; // @[:@135030.4]
  assign RetimeWrapper_reset = reset; // @[:@135031.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@135032.4]
endmodule
module FringeCounter( // @[:@135048.2]
  input   clock, // @[:@135049.4]
  input   reset, // @[:@135050.4]
  input   io_enable, // @[:@135051.4]
  output  io_done // @[:@135051.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@135053.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@135053.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@135053.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@135053.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@135053.4]
  wire [40:0] count; // @[Cat.scala 30:58:@135060.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@135061.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@135062.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@135063.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@135065.4]
  FringeFF_503 reg$ ( // @[FringeCounter.scala 24:19:@135053.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@135060.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@135061.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@135062.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@135063.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@135065.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@135076.4]
  assign reg$_clock = clock; // @[:@135054.4]
  assign reg$_reset = reset; // @[:@135055.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@135067.6 FringeCounter.scala 37:15:@135070.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@135058.4]
endmodule
module FringeFF_504( // @[:@135110.2]
  input   clock, // @[:@135111.4]
  input   reset, // @[:@135112.4]
  input   io_in, // @[:@135113.4]
  input   io_reset, // @[:@135113.4]
  output  io_out, // @[:@135113.4]
  input   io_enable // @[:@135113.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@135116.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@135116.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@135116.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@135116.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@135116.4]
  wire  _T_18; // @[package.scala 96:25:@135121.4 package.scala 96:25:@135122.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@135127.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@135116.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@135121.4 package.scala 96:25:@135122.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@135127.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@135133.4]
  assign RetimeWrapper_clock = clock; // @[:@135117.4]
  assign RetimeWrapper_reset = reset; // @[:@135118.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@135120.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@135119.4]
endmodule
module Depulser( // @[:@135135.2]
  input   clock, // @[:@135136.4]
  input   reset, // @[:@135137.4]
  input   io_in, // @[:@135138.4]
  input   io_rst, // @[:@135138.4]
  output  io_out // @[:@135138.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@135140.4]
  wire  r_reset; // @[Depulser.scala 14:17:@135140.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@135140.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@135140.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@135140.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@135140.4]
  FringeFF_504 r ( // @[Depulser.scala 14:17:@135140.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@135149.4]
  assign r_clock = clock; // @[:@135141.4]
  assign r_reset = reset; // @[:@135142.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@135144.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@135148.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@135147.4]
endmodule
module Fringe( // @[:@135151.2]
  input         clock, // @[:@135152.4]
  input         reset, // @[:@135153.4]
  input  [31:0] io_raddr, // @[:@135154.4]
  input         io_wen, // @[:@135154.4]
  input  [31:0] io_waddr, // @[:@135154.4]
  input  [63:0] io_wdata, // @[:@135154.4]
  output [63:0] io_rdata, // @[:@135154.4]
  output        io_enable, // @[:@135154.4]
  input         io_done, // @[:@135154.4]
  output        io_reset, // @[:@135154.4]
  output [63:0] io_argIns_0, // @[:@135154.4]
  output [63:0] io_argIns_1, // @[:@135154.4]
  input         io_argOuts_0_valid, // @[:@135154.4]
  input  [63:0] io_argOuts_0_bits, // @[:@135154.4]
  output        io_memStreams_stores_0_cmd_ready, // @[:@135154.4]
  input         io_memStreams_stores_0_cmd_valid, // @[:@135154.4]
  input  [63:0] io_memStreams_stores_0_cmd_bits_addr, // @[:@135154.4]
  input  [31:0] io_memStreams_stores_0_cmd_bits_size, // @[:@135154.4]
  output        io_memStreams_stores_0_data_ready, // @[:@135154.4]
  input         io_memStreams_stores_0_data_valid, // @[:@135154.4]
  input  [31:0] io_memStreams_stores_0_data_bits_wdata_0, // @[:@135154.4]
  input         io_memStreams_stores_0_data_bits_wstrb, // @[:@135154.4]
  input         io_memStreams_stores_0_wresp_ready, // @[:@135154.4]
  output        io_memStreams_stores_0_wresp_valid, // @[:@135154.4]
  output        io_memStreams_stores_0_wresp_bits, // @[:@135154.4]
  input         io_dram_0_cmd_ready, // @[:@135154.4]
  output        io_dram_0_cmd_valid, // @[:@135154.4]
  output [63:0] io_dram_0_cmd_bits_addr, // @[:@135154.4]
  output [31:0] io_dram_0_cmd_bits_size, // @[:@135154.4]
  output        io_dram_0_cmd_bits_isWr, // @[:@135154.4]
  output [31:0] io_dram_0_cmd_bits_tag, // @[:@135154.4]
  input         io_dram_0_wdata_ready, // @[:@135154.4]
  output        io_dram_0_wdata_valid, // @[:@135154.4]
  output [31:0] io_dram_0_wdata_bits_wdata_0, // @[:@135154.4]
  output [31:0] io_dram_0_wdata_bits_wdata_1, // @[:@135154.4]
  output [31:0] io_dram_0_wdata_bits_wdata_2, // @[:@135154.4]
  output [31:0] io_dram_0_wdata_bits_wdata_3, // @[:@135154.4]
  output [31:0] io_dram_0_wdata_bits_wdata_4, // @[:@135154.4]
  output [31:0] io_dram_0_wdata_bits_wdata_5, // @[:@135154.4]
  output [31:0] io_dram_0_wdata_bits_wdata_6, // @[:@135154.4]
  output [31:0] io_dram_0_wdata_bits_wdata_7, // @[:@135154.4]
  output [31:0] io_dram_0_wdata_bits_wdata_8, // @[:@135154.4]
  output [31:0] io_dram_0_wdata_bits_wdata_9, // @[:@135154.4]
  output [31:0] io_dram_0_wdata_bits_wdata_10, // @[:@135154.4]
  output [31:0] io_dram_0_wdata_bits_wdata_11, // @[:@135154.4]
  output [31:0] io_dram_0_wdata_bits_wdata_12, // @[:@135154.4]
  output [31:0] io_dram_0_wdata_bits_wdata_13, // @[:@135154.4]
  output [31:0] io_dram_0_wdata_bits_wdata_14, // @[:@135154.4]
  output [31:0] io_dram_0_wdata_bits_wdata_15, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_0, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_1, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_2, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_3, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_4, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_5, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_6, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_7, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_8, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_9, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_10, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_11, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_12, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_13, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_14, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_15, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_16, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_17, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_18, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_19, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_20, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_21, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_22, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_23, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_24, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_25, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_26, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_27, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_28, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_29, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_30, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_31, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_32, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_33, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_34, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_35, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_36, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_37, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_38, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_39, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_40, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_41, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_42, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_43, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_44, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_45, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_46, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_47, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_48, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_49, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_50, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_51, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_52, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_53, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_54, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_55, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_56, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_57, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_58, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_59, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_60, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_61, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_62, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wstrb_63, // @[:@135154.4]
  output        io_dram_0_wdata_bits_wlast, // @[:@135154.4]
  output        io_dram_0_rresp_ready, // @[:@135154.4]
  output        io_dram_0_wresp_ready, // @[:@135154.4]
  input         io_dram_0_wresp_valid, // @[:@135154.4]
  input  [31:0] io_dram_0_wresp_bits_tag, // @[:@135154.4]
  input         io_dram_1_cmd_ready, // @[:@135154.4]
  output        io_dram_1_cmd_valid, // @[:@135154.4]
  output [63:0] io_dram_1_cmd_bits_addr, // @[:@135154.4]
  output [31:0] io_dram_1_cmd_bits_size, // @[:@135154.4]
  output        io_dram_1_cmd_bits_isWr, // @[:@135154.4]
  output [31:0] io_dram_1_cmd_bits_tag, // @[:@135154.4]
  input         io_dram_1_wdata_ready, // @[:@135154.4]
  output        io_dram_1_wdata_valid, // @[:@135154.4]
  output [31:0] io_dram_1_wdata_bits_wdata_0, // @[:@135154.4]
  output [31:0] io_dram_1_wdata_bits_wdata_1, // @[:@135154.4]
  output [31:0] io_dram_1_wdata_bits_wdata_2, // @[:@135154.4]
  output [31:0] io_dram_1_wdata_bits_wdata_3, // @[:@135154.4]
  output [31:0] io_dram_1_wdata_bits_wdata_4, // @[:@135154.4]
  output [31:0] io_dram_1_wdata_bits_wdata_5, // @[:@135154.4]
  output [31:0] io_dram_1_wdata_bits_wdata_6, // @[:@135154.4]
  output [31:0] io_dram_1_wdata_bits_wdata_7, // @[:@135154.4]
  output [31:0] io_dram_1_wdata_bits_wdata_8, // @[:@135154.4]
  output [31:0] io_dram_1_wdata_bits_wdata_9, // @[:@135154.4]
  output [31:0] io_dram_1_wdata_bits_wdata_10, // @[:@135154.4]
  output [31:0] io_dram_1_wdata_bits_wdata_11, // @[:@135154.4]
  output [31:0] io_dram_1_wdata_bits_wdata_12, // @[:@135154.4]
  output [31:0] io_dram_1_wdata_bits_wdata_13, // @[:@135154.4]
  output [31:0] io_dram_1_wdata_bits_wdata_14, // @[:@135154.4]
  output [31:0] io_dram_1_wdata_bits_wdata_15, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_0, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_1, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_2, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_3, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_4, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_5, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_6, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_7, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_8, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_9, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_10, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_11, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_12, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_13, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_14, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_15, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_16, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_17, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_18, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_19, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_20, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_21, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_22, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_23, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_24, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_25, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_26, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_27, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_28, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_29, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_30, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_31, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_32, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_33, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_34, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_35, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_36, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_37, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_38, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_39, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_40, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_41, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_42, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_43, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_44, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_45, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_46, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_47, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_48, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_49, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_50, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_51, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_52, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_53, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_54, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_55, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_56, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_57, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_58, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_59, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_60, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_61, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_62, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wstrb_63, // @[:@135154.4]
  output        io_dram_1_wdata_bits_wlast, // @[:@135154.4]
  output        io_dram_1_rresp_ready, // @[:@135154.4]
  output        io_dram_1_wresp_ready, // @[:@135154.4]
  input         io_dram_1_wresp_valid, // @[:@135154.4]
  input  [31:0] io_dram_1_wresp_bits_tag, // @[:@135154.4]
  input         io_dram_2_cmd_ready, // @[:@135154.4]
  output        io_dram_2_cmd_valid, // @[:@135154.4]
  output [63:0] io_dram_2_cmd_bits_addr, // @[:@135154.4]
  output [31:0] io_dram_2_cmd_bits_size, // @[:@135154.4]
  output        io_dram_2_cmd_bits_isWr, // @[:@135154.4]
  output [31:0] io_dram_2_cmd_bits_tag, // @[:@135154.4]
  input         io_dram_2_wdata_ready, // @[:@135154.4]
  output        io_dram_2_wdata_valid, // @[:@135154.4]
  output [31:0] io_dram_2_wdata_bits_wdata_0, // @[:@135154.4]
  output [31:0] io_dram_2_wdata_bits_wdata_1, // @[:@135154.4]
  output [31:0] io_dram_2_wdata_bits_wdata_2, // @[:@135154.4]
  output [31:0] io_dram_2_wdata_bits_wdata_3, // @[:@135154.4]
  output [31:0] io_dram_2_wdata_bits_wdata_4, // @[:@135154.4]
  output [31:0] io_dram_2_wdata_bits_wdata_5, // @[:@135154.4]
  output [31:0] io_dram_2_wdata_bits_wdata_6, // @[:@135154.4]
  output [31:0] io_dram_2_wdata_bits_wdata_7, // @[:@135154.4]
  output [31:0] io_dram_2_wdata_bits_wdata_8, // @[:@135154.4]
  output [31:0] io_dram_2_wdata_bits_wdata_9, // @[:@135154.4]
  output [31:0] io_dram_2_wdata_bits_wdata_10, // @[:@135154.4]
  output [31:0] io_dram_2_wdata_bits_wdata_11, // @[:@135154.4]
  output [31:0] io_dram_2_wdata_bits_wdata_12, // @[:@135154.4]
  output [31:0] io_dram_2_wdata_bits_wdata_13, // @[:@135154.4]
  output [31:0] io_dram_2_wdata_bits_wdata_14, // @[:@135154.4]
  output [31:0] io_dram_2_wdata_bits_wdata_15, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_0, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_1, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_2, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_3, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_4, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_5, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_6, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_7, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_8, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_9, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_10, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_11, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_12, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_13, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_14, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_15, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_16, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_17, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_18, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_19, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_20, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_21, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_22, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_23, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_24, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_25, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_26, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_27, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_28, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_29, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_30, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_31, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_32, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_33, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_34, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_35, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_36, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_37, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_38, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_39, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_40, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_41, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_42, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_43, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_44, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_45, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_46, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_47, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_48, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_49, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_50, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_51, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_52, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_53, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_54, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_55, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_56, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_57, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_58, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_59, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_60, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_61, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_62, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wstrb_63, // @[:@135154.4]
  output        io_dram_2_wdata_bits_wlast, // @[:@135154.4]
  output        io_dram_2_rresp_ready, // @[:@135154.4]
  output        io_dram_2_wresp_ready, // @[:@135154.4]
  input         io_dram_2_wresp_valid, // @[:@135154.4]
  input  [31:0] io_dram_2_wresp_bits_tag, // @[:@135154.4]
  input         io_dram_3_cmd_ready, // @[:@135154.4]
  output        io_dram_3_cmd_valid, // @[:@135154.4]
  output [63:0] io_dram_3_cmd_bits_addr, // @[:@135154.4]
  output [31:0] io_dram_3_cmd_bits_size, // @[:@135154.4]
  output        io_dram_3_cmd_bits_isWr, // @[:@135154.4]
  output [31:0] io_dram_3_cmd_bits_tag, // @[:@135154.4]
  input         io_dram_3_wdata_ready, // @[:@135154.4]
  output        io_dram_3_wdata_valid, // @[:@135154.4]
  output [31:0] io_dram_3_wdata_bits_wdata_0, // @[:@135154.4]
  output [31:0] io_dram_3_wdata_bits_wdata_1, // @[:@135154.4]
  output [31:0] io_dram_3_wdata_bits_wdata_2, // @[:@135154.4]
  output [31:0] io_dram_3_wdata_bits_wdata_3, // @[:@135154.4]
  output [31:0] io_dram_3_wdata_bits_wdata_4, // @[:@135154.4]
  output [31:0] io_dram_3_wdata_bits_wdata_5, // @[:@135154.4]
  output [31:0] io_dram_3_wdata_bits_wdata_6, // @[:@135154.4]
  output [31:0] io_dram_3_wdata_bits_wdata_7, // @[:@135154.4]
  output [31:0] io_dram_3_wdata_bits_wdata_8, // @[:@135154.4]
  output [31:0] io_dram_3_wdata_bits_wdata_9, // @[:@135154.4]
  output [31:0] io_dram_3_wdata_bits_wdata_10, // @[:@135154.4]
  output [31:0] io_dram_3_wdata_bits_wdata_11, // @[:@135154.4]
  output [31:0] io_dram_3_wdata_bits_wdata_12, // @[:@135154.4]
  output [31:0] io_dram_3_wdata_bits_wdata_13, // @[:@135154.4]
  output [31:0] io_dram_3_wdata_bits_wdata_14, // @[:@135154.4]
  output [31:0] io_dram_3_wdata_bits_wdata_15, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_0, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_1, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_2, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_3, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_4, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_5, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_6, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_7, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_8, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_9, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_10, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_11, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_12, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_13, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_14, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_15, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_16, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_17, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_18, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_19, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_20, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_21, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_22, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_23, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_24, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_25, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_26, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_27, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_28, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_29, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_30, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_31, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_32, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_33, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_34, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_35, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_36, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_37, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_38, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_39, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_40, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_41, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_42, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_43, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_44, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_45, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_46, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_47, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_48, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_49, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_50, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_51, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_52, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_53, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_54, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_55, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_56, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_57, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_58, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_59, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_60, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_61, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_62, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wstrb_63, // @[:@135154.4]
  output        io_dram_3_wdata_bits_wlast, // @[:@135154.4]
  output        io_dram_3_rresp_ready, // @[:@135154.4]
  output        io_dram_3_wresp_ready, // @[:@135154.4]
  input         io_dram_3_wresp_valid, // @[:@135154.4]
  input  [31:0] io_dram_3_wresp_bits_tag, // @[:@135154.4]
  input         io_heap_0_req_valid, // @[:@135154.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@135154.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@135154.4]
  output        io_heap_0_resp_valid, // @[:@135154.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@135154.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@135154.4]
);
  wire  dramArbs_0_clock; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_reset; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_enable; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_app_stores_0_cmd_valid; // @[Fringe.scala 91:25:@135160.4]
  wire [63:0] dramArbs_0_io_app_stores_0_cmd_bits_addr; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_app_stores_0_cmd_bits_size; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_app_stores_0_data_valid; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_app_stores_0_data_bits_wdata_0; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_app_stores_0_data_bits_wstrb; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_app_stores_0_wresp_ready; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_cmd_ready; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 91:25:@135160.4]
  wire [63:0] dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_ready; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_0_io_dram_wresp_valid; // @[Fringe.scala 91:25:@135160.4]
  wire [31:0] dramArbs_0_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@135160.4]
  wire  dramArbs_1_clock; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_reset; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_enable; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_cmd_ready; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 91:25:@136153.4]
  wire [63:0] dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_ready; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_1_io_dram_wresp_valid; // @[Fringe.scala 91:25:@136153.4]
  wire [31:0] dramArbs_1_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@136153.4]
  wire  dramArbs_2_clock; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_reset; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_enable; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_cmd_ready; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 91:25:@137113.4]
  wire [63:0] dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_ready; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_2_io_dram_wresp_valid; // @[Fringe.scala 91:25:@137113.4]
  wire [31:0] dramArbs_2_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@137113.4]
  wire  dramArbs_3_clock; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_reset; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_enable; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_cmd_ready; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 91:25:@138073.4]
  wire [63:0] dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_ready; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 91:25:@138073.4]
  wire  dramArbs_3_io_dram_wresp_valid; // @[Fringe.scala 91:25:@138073.4]
  wire [31:0] dramArbs_3_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@138073.4]
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@139033.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@139033.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@139033.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@139033.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@139033.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@139033.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@139033.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@139033.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@139033.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@139033.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@139033.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@139033.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@139042.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@139042.4]
  wire [31:0] regs_io_raddr; // @[Fringe.scala 116:20:@139042.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@139042.4]
  wire [31:0] regs_io_waddr; // @[Fringe.scala 116:20:@139042.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@139042.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@139042.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@139042.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@139042.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@139042.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@139042.4]
  wire [63:0] regs_io_argIns_3; // @[Fringe.scala 116:20:@139042.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@139042.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@139042.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@139042.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@139042.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@141092.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@141092.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@141092.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@141092.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@141111.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@141111.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@141111.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@141111.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@141111.4]
  wire [63:0] _T_1020; // @[:@141069.4 :@141070.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@141071.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@141073.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@141075.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@141077.4]
  wire  _T_1025; // @[Fringe.scala 134:28:@141079.4]
  wire  _T_1029; // @[Fringe.scala 134:42:@141081.4]
  wire  _T_1030; // @[Fringe.scala 135:27:@141083.4]
  wire [63:0] _T_1040; // @[Fringe.scala 156:22:@141119.4]
  reg  _T_1047; // @[package.scala 152:20:@141122.4]
  reg [31:0] _RAND_0;
  wire  _T_1048; // @[package.scala 153:13:@141124.4]
  wire  _T_1049; // @[package.scala 153:8:@141125.4]
  wire  _T_1052; // @[Fringe.scala 160:55:@141129.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@141130.4]
  wire  _T_1055; // @[Fringe.scala 161:58:@141133.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@141134.4]
  wire [1:0] _T_1059; // @[Fringe.scala 162:57:@141136.4]
  wire [1:0] _T_1061; // @[Fringe.scala 162:34:@141137.4]
  wire [63:0] _T_1063; // @[Fringe.scala 163:30:@141139.4]
  wire [1:0] _T_1064; // @[Fringe.scala 171:37:@141142.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@141121.4 Fringe.scala 163:24:@141140.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@141121.4 Fringe.scala 162:28:@141138.4]
  wire [61:0] _T_1065; // @[Fringe.scala 171:37:@141143.4]
  wire  alloc; // @[Fringe.scala 202:38:@142773.4]
  wire  dealloc; // @[Fringe.scala 203:40:@142774.4]
  wire  _T_1569; // @[Fringe.scala 204:37:@142775.4]
  reg  _T_1572; // @[package.scala 152:20:@142776.4]
  reg [31:0] _RAND_1;
  wire  _T_1573; // @[package.scala 153:13:@142778.4]
  DRAMArbiter dramArbs_0 ( // @[Fringe.scala 91:25:@135160.4]
    .clock(dramArbs_0_clock),
    .reset(dramArbs_0_reset),
    .io_enable(dramArbs_0_io_enable),
    .io_app_stores_0_cmd_ready(dramArbs_0_io_app_stores_0_cmd_ready),
    .io_app_stores_0_cmd_valid(dramArbs_0_io_app_stores_0_cmd_valid),
    .io_app_stores_0_cmd_bits_addr(dramArbs_0_io_app_stores_0_cmd_bits_addr),
    .io_app_stores_0_cmd_bits_size(dramArbs_0_io_app_stores_0_cmd_bits_size),
    .io_app_stores_0_data_ready(dramArbs_0_io_app_stores_0_data_ready),
    .io_app_stores_0_data_valid(dramArbs_0_io_app_stores_0_data_valid),
    .io_app_stores_0_data_bits_wdata_0(dramArbs_0_io_app_stores_0_data_bits_wdata_0),
    .io_app_stores_0_data_bits_wstrb(dramArbs_0_io_app_stores_0_data_bits_wstrb),
    .io_app_stores_0_wresp_ready(dramArbs_0_io_app_stores_0_wresp_ready),
    .io_app_stores_0_wresp_valid(dramArbs_0_io_app_stores_0_wresp_valid),
    .io_app_stores_0_wresp_bits(dramArbs_0_io_app_stores_0_wresp_bits),
    .io_dram_cmd_ready(dramArbs_0_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_0_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_0_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_0_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_0_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_0_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_0_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_0_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_0_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_0_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_0_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_0_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_0_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_0_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_0_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_0_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_0_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_0_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_0_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_0_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_0_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_0_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_0_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_0_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_0_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_0_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_0_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_0_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_0_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_0_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_0_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_0_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_0_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_0_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_0_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_0_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_0_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_0_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_0_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_0_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_0_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_0_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_0_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_0_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_0_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_0_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_0_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_0_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_0_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_0_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_0_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_0_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_0_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_0_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_0_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_0_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_0_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_0_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_0_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_0_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_0_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_0_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_0_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_0_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_0_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_0_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_0_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_0_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_0_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_0_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_0_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_0_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_0_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_0_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_0_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_0_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_0_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_0_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_0_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_0_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_0_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_0_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_0_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_0_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_0_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_0_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_0_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_0_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_0_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_0_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_0_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_0_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_0_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_1 ( // @[Fringe.scala 91:25:@136153.4]
    .clock(dramArbs_1_clock),
    .reset(dramArbs_1_reset),
    .io_enable(dramArbs_1_io_enable),
    .io_dram_cmd_ready(dramArbs_1_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_1_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_1_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_1_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_1_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_1_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_1_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_1_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_1_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_1_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_1_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_1_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_1_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_1_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_1_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_1_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_1_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_1_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_1_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_1_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_1_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_1_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_1_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_1_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_1_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_1_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_1_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_1_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_1_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_1_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_1_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_1_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_1_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_1_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_1_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_1_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_1_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_1_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_1_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_1_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_1_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_1_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_1_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_1_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_1_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_1_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_1_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_1_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_1_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_1_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_1_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_1_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_1_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_1_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_1_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_1_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_1_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_1_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_1_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_1_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_1_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_1_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_1_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_1_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_1_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_1_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_1_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_1_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_1_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_1_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_1_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_1_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_1_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_1_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_1_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_1_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_1_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_1_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_1_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_1_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_1_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_1_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_1_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_1_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_1_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_1_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_1_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_1_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_1_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_1_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_1_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_1_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_1_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_2 ( // @[Fringe.scala 91:25:@137113.4]
    .clock(dramArbs_2_clock),
    .reset(dramArbs_2_reset),
    .io_enable(dramArbs_2_io_enable),
    .io_dram_cmd_ready(dramArbs_2_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_2_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_2_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_2_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_2_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_2_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_2_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_2_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_2_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_2_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_2_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_2_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_2_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_2_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_2_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_2_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_2_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_2_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_2_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_2_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_2_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_2_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_2_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_2_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_2_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_2_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_2_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_2_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_2_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_2_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_2_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_2_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_2_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_2_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_2_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_2_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_2_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_2_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_2_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_2_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_2_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_2_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_2_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_2_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_2_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_2_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_2_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_2_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_2_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_2_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_2_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_2_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_2_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_2_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_2_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_2_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_2_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_2_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_2_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_2_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_2_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_2_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_2_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_2_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_2_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_2_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_2_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_2_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_2_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_2_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_2_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_2_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_2_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_2_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_2_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_2_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_2_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_2_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_2_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_2_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_2_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_2_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_2_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_2_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_2_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_2_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_2_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_2_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_2_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_2_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_2_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_2_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_2_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_3 ( // @[Fringe.scala 91:25:@138073.4]
    .clock(dramArbs_3_clock),
    .reset(dramArbs_3_reset),
    .io_enable(dramArbs_3_io_enable),
    .io_dram_cmd_ready(dramArbs_3_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_3_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_3_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_3_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_3_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_3_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_3_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_3_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_3_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_3_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_3_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_3_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_3_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_3_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_3_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_3_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_3_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_3_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_3_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_3_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_3_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_3_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_3_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_3_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_3_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_3_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_3_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_3_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_3_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_3_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_3_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_3_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_3_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_3_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_3_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_3_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_3_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_3_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_3_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_3_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_3_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_3_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_3_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_3_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_3_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_3_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_3_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_3_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_3_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_3_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_3_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_3_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_3_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_3_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_3_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_3_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_3_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_3_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_3_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_3_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_3_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_3_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_3_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_3_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_3_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_3_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_3_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_3_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_3_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_3_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_3_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_3_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_3_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_3_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_3_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_3_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_3_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_3_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_3_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_3_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_3_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_3_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_3_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_3_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_3_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_3_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_3_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_3_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_3_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_3_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_3_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_3_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_3_io_dram_wresp_bits_tag)
  );
  DRAMHeap heap ( // @[Fringe.scala 107:20:@139033.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@139042.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argIns_3(regs_io_argIns_3),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@141092.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@141111.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_1020 = regs_io_argIns_1; // @[:@141069.4 :@141070.4]
  assign curStatus_done = _T_1020[0]; // @[Fringe.scala 133:45:@141071.4]
  assign curStatus_timeout = _T_1020[1]; // @[Fringe.scala 133:45:@141073.4]
  assign curStatus_allocDealloc = _T_1020[4:2]; // @[Fringe.scala 133:45:@141075.4]
  assign curStatus_sizeAddr = _T_1020[63:5]; // @[Fringe.scala 133:45:@141077.4]
  assign _T_1025 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@141079.4]
  assign _T_1029 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@141081.4]
  assign _T_1030 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@141083.4]
  assign _T_1040 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@141119.4]
  assign _T_1048 = _T_1047 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@141124.4]
  assign _T_1049 = heap_io_host_0_req_valid & _T_1048; // @[package.scala 153:8:@141125.4]
  assign _T_1052 = _T_1025 & depulser_io_out; // @[Fringe.scala 160:55:@141129.4]
  assign status_bits_done = depulser_io_out ? _T_1052 : curStatus_done; // @[Fringe.scala 160:26:@141130.4]
  assign _T_1055 = _T_1025 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@141133.4]
  assign status_bits_timeout = depulser_io_out ? _T_1055 : curStatus_timeout; // @[Fringe.scala 161:29:@141134.4]
  assign _T_1059 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@141136.4]
  assign _T_1061 = heap_io_host_0_req_valid ? _T_1059 : 2'h0; // @[Fringe.scala 162:34:@141137.4]
  assign _T_1063 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@141139.4]
  assign _T_1064 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@141142.4]
  assign status_bits_sizeAddr = _T_1063[58:0]; // @[Fringe.scala 158:20:@141121.4 Fringe.scala 163:24:@141140.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_1061}; // @[Fringe.scala 158:20:@141121.4 Fringe.scala 162:28:@141138.4]
  assign _T_1065 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@141143.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@142773.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@142774.4]
  assign _T_1569 = alloc | dealloc; // @[Fringe.scala 204:37:@142775.4]
  assign _T_1573 = _T_1572 ^ _T_1569; // @[package.scala 153:13:@142778.4]
  assign io_rdata = regs_io_rdata; // @[Fringe.scala 125:14:@141067.4]
  assign io_enable = _T_1025 & _T_1029; // @[Fringe.scala 136:13:@141087.4]
  assign io_reset = _T_1030 | reset; // @[Fringe.scala 137:12:@141088.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@141109.4]
  assign io_argIns_1 = regs_io_argIns_3; // @[Fringe.scala 151:51:@141110.4]
  assign io_memStreams_stores_0_cmd_ready = dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 101:72:@136079.4]
  assign io_memStreams_stores_0_data_ready = dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 101:72:@136075.4]
  assign io_memStreams_stores_0_wresp_valid = dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 101:72:@136070.4]
  assign io_memStreams_stores_0_wresp_bits = dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 101:72:@136069.4]
  assign io_dram_0_cmd_valid = dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 195:72:@142271.4]
  assign io_dram_0_cmd_bits_addr = dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@142270.4]
  assign io_dram_0_cmd_bits_size = dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@142269.4]
  assign io_dram_0_cmd_bits_isWr = dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@142267.4]
  assign io_dram_0_cmd_bits_tag = dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@142266.4]
  assign io_dram_0_wdata_valid = dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 195:72:@142264.4]
  assign io_dram_0_wdata_bits_wdata_0 = dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@142248.4]
  assign io_dram_0_wdata_bits_wdata_1 = dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@142249.4]
  assign io_dram_0_wdata_bits_wdata_2 = dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@142250.4]
  assign io_dram_0_wdata_bits_wdata_3 = dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@142251.4]
  assign io_dram_0_wdata_bits_wdata_4 = dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@142252.4]
  assign io_dram_0_wdata_bits_wdata_5 = dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@142253.4]
  assign io_dram_0_wdata_bits_wdata_6 = dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@142254.4]
  assign io_dram_0_wdata_bits_wdata_7 = dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@142255.4]
  assign io_dram_0_wdata_bits_wdata_8 = dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@142256.4]
  assign io_dram_0_wdata_bits_wdata_9 = dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@142257.4]
  assign io_dram_0_wdata_bits_wdata_10 = dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@142258.4]
  assign io_dram_0_wdata_bits_wdata_11 = dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@142259.4]
  assign io_dram_0_wdata_bits_wdata_12 = dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@142260.4]
  assign io_dram_0_wdata_bits_wdata_13 = dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@142261.4]
  assign io_dram_0_wdata_bits_wdata_14 = dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@142262.4]
  assign io_dram_0_wdata_bits_wdata_15 = dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@142263.4]
  assign io_dram_0_wdata_bits_wstrb_0 = dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@142184.4]
  assign io_dram_0_wdata_bits_wstrb_1 = dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@142185.4]
  assign io_dram_0_wdata_bits_wstrb_2 = dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@142186.4]
  assign io_dram_0_wdata_bits_wstrb_3 = dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@142187.4]
  assign io_dram_0_wdata_bits_wstrb_4 = dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@142188.4]
  assign io_dram_0_wdata_bits_wstrb_5 = dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@142189.4]
  assign io_dram_0_wdata_bits_wstrb_6 = dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@142190.4]
  assign io_dram_0_wdata_bits_wstrb_7 = dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@142191.4]
  assign io_dram_0_wdata_bits_wstrb_8 = dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@142192.4]
  assign io_dram_0_wdata_bits_wstrb_9 = dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@142193.4]
  assign io_dram_0_wdata_bits_wstrb_10 = dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@142194.4]
  assign io_dram_0_wdata_bits_wstrb_11 = dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@142195.4]
  assign io_dram_0_wdata_bits_wstrb_12 = dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@142196.4]
  assign io_dram_0_wdata_bits_wstrb_13 = dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@142197.4]
  assign io_dram_0_wdata_bits_wstrb_14 = dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@142198.4]
  assign io_dram_0_wdata_bits_wstrb_15 = dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@142199.4]
  assign io_dram_0_wdata_bits_wstrb_16 = dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@142200.4]
  assign io_dram_0_wdata_bits_wstrb_17 = dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@142201.4]
  assign io_dram_0_wdata_bits_wstrb_18 = dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@142202.4]
  assign io_dram_0_wdata_bits_wstrb_19 = dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@142203.4]
  assign io_dram_0_wdata_bits_wstrb_20 = dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@142204.4]
  assign io_dram_0_wdata_bits_wstrb_21 = dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@142205.4]
  assign io_dram_0_wdata_bits_wstrb_22 = dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@142206.4]
  assign io_dram_0_wdata_bits_wstrb_23 = dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@142207.4]
  assign io_dram_0_wdata_bits_wstrb_24 = dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@142208.4]
  assign io_dram_0_wdata_bits_wstrb_25 = dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@142209.4]
  assign io_dram_0_wdata_bits_wstrb_26 = dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@142210.4]
  assign io_dram_0_wdata_bits_wstrb_27 = dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@142211.4]
  assign io_dram_0_wdata_bits_wstrb_28 = dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@142212.4]
  assign io_dram_0_wdata_bits_wstrb_29 = dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@142213.4]
  assign io_dram_0_wdata_bits_wstrb_30 = dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@142214.4]
  assign io_dram_0_wdata_bits_wstrb_31 = dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@142215.4]
  assign io_dram_0_wdata_bits_wstrb_32 = dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@142216.4]
  assign io_dram_0_wdata_bits_wstrb_33 = dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@142217.4]
  assign io_dram_0_wdata_bits_wstrb_34 = dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@142218.4]
  assign io_dram_0_wdata_bits_wstrb_35 = dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@142219.4]
  assign io_dram_0_wdata_bits_wstrb_36 = dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@142220.4]
  assign io_dram_0_wdata_bits_wstrb_37 = dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@142221.4]
  assign io_dram_0_wdata_bits_wstrb_38 = dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@142222.4]
  assign io_dram_0_wdata_bits_wstrb_39 = dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@142223.4]
  assign io_dram_0_wdata_bits_wstrb_40 = dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@142224.4]
  assign io_dram_0_wdata_bits_wstrb_41 = dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@142225.4]
  assign io_dram_0_wdata_bits_wstrb_42 = dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@142226.4]
  assign io_dram_0_wdata_bits_wstrb_43 = dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@142227.4]
  assign io_dram_0_wdata_bits_wstrb_44 = dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@142228.4]
  assign io_dram_0_wdata_bits_wstrb_45 = dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@142229.4]
  assign io_dram_0_wdata_bits_wstrb_46 = dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@142230.4]
  assign io_dram_0_wdata_bits_wstrb_47 = dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@142231.4]
  assign io_dram_0_wdata_bits_wstrb_48 = dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@142232.4]
  assign io_dram_0_wdata_bits_wstrb_49 = dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@142233.4]
  assign io_dram_0_wdata_bits_wstrb_50 = dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@142234.4]
  assign io_dram_0_wdata_bits_wstrb_51 = dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@142235.4]
  assign io_dram_0_wdata_bits_wstrb_52 = dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@142236.4]
  assign io_dram_0_wdata_bits_wstrb_53 = dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@142237.4]
  assign io_dram_0_wdata_bits_wstrb_54 = dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@142238.4]
  assign io_dram_0_wdata_bits_wstrb_55 = dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@142239.4]
  assign io_dram_0_wdata_bits_wstrb_56 = dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@142240.4]
  assign io_dram_0_wdata_bits_wstrb_57 = dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@142241.4]
  assign io_dram_0_wdata_bits_wstrb_58 = dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@142242.4]
  assign io_dram_0_wdata_bits_wstrb_59 = dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@142243.4]
  assign io_dram_0_wdata_bits_wstrb_60 = dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@142244.4]
  assign io_dram_0_wdata_bits_wstrb_61 = dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@142245.4]
  assign io_dram_0_wdata_bits_wstrb_62 = dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@142246.4]
  assign io_dram_0_wdata_bits_wstrb_63 = dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@142247.4]
  assign io_dram_0_wdata_bits_wlast = dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@142183.4]
  assign io_dram_0_rresp_ready = dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 195:72:@142182.4]
  assign io_dram_0_wresp_ready = dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 195:72:@142163.4]
  assign io_dram_1_cmd_valid = dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 195:72:@142383.4]
  assign io_dram_1_cmd_bits_addr = dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@142382.4]
  assign io_dram_1_cmd_bits_size = dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@142381.4]
  assign io_dram_1_cmd_bits_isWr = dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@142379.4]
  assign io_dram_1_cmd_bits_tag = dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@142378.4]
  assign io_dram_1_wdata_valid = dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 195:72:@142376.4]
  assign io_dram_1_wdata_bits_wdata_0 = dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@142360.4]
  assign io_dram_1_wdata_bits_wdata_1 = dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@142361.4]
  assign io_dram_1_wdata_bits_wdata_2 = dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@142362.4]
  assign io_dram_1_wdata_bits_wdata_3 = dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@142363.4]
  assign io_dram_1_wdata_bits_wdata_4 = dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@142364.4]
  assign io_dram_1_wdata_bits_wdata_5 = dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@142365.4]
  assign io_dram_1_wdata_bits_wdata_6 = dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@142366.4]
  assign io_dram_1_wdata_bits_wdata_7 = dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@142367.4]
  assign io_dram_1_wdata_bits_wdata_8 = dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@142368.4]
  assign io_dram_1_wdata_bits_wdata_9 = dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@142369.4]
  assign io_dram_1_wdata_bits_wdata_10 = dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@142370.4]
  assign io_dram_1_wdata_bits_wdata_11 = dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@142371.4]
  assign io_dram_1_wdata_bits_wdata_12 = dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@142372.4]
  assign io_dram_1_wdata_bits_wdata_13 = dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@142373.4]
  assign io_dram_1_wdata_bits_wdata_14 = dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@142374.4]
  assign io_dram_1_wdata_bits_wdata_15 = dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@142375.4]
  assign io_dram_1_wdata_bits_wstrb_0 = dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@142296.4]
  assign io_dram_1_wdata_bits_wstrb_1 = dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@142297.4]
  assign io_dram_1_wdata_bits_wstrb_2 = dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@142298.4]
  assign io_dram_1_wdata_bits_wstrb_3 = dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@142299.4]
  assign io_dram_1_wdata_bits_wstrb_4 = dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@142300.4]
  assign io_dram_1_wdata_bits_wstrb_5 = dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@142301.4]
  assign io_dram_1_wdata_bits_wstrb_6 = dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@142302.4]
  assign io_dram_1_wdata_bits_wstrb_7 = dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@142303.4]
  assign io_dram_1_wdata_bits_wstrb_8 = dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@142304.4]
  assign io_dram_1_wdata_bits_wstrb_9 = dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@142305.4]
  assign io_dram_1_wdata_bits_wstrb_10 = dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@142306.4]
  assign io_dram_1_wdata_bits_wstrb_11 = dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@142307.4]
  assign io_dram_1_wdata_bits_wstrb_12 = dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@142308.4]
  assign io_dram_1_wdata_bits_wstrb_13 = dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@142309.4]
  assign io_dram_1_wdata_bits_wstrb_14 = dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@142310.4]
  assign io_dram_1_wdata_bits_wstrb_15 = dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@142311.4]
  assign io_dram_1_wdata_bits_wstrb_16 = dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@142312.4]
  assign io_dram_1_wdata_bits_wstrb_17 = dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@142313.4]
  assign io_dram_1_wdata_bits_wstrb_18 = dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@142314.4]
  assign io_dram_1_wdata_bits_wstrb_19 = dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@142315.4]
  assign io_dram_1_wdata_bits_wstrb_20 = dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@142316.4]
  assign io_dram_1_wdata_bits_wstrb_21 = dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@142317.4]
  assign io_dram_1_wdata_bits_wstrb_22 = dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@142318.4]
  assign io_dram_1_wdata_bits_wstrb_23 = dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@142319.4]
  assign io_dram_1_wdata_bits_wstrb_24 = dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@142320.4]
  assign io_dram_1_wdata_bits_wstrb_25 = dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@142321.4]
  assign io_dram_1_wdata_bits_wstrb_26 = dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@142322.4]
  assign io_dram_1_wdata_bits_wstrb_27 = dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@142323.4]
  assign io_dram_1_wdata_bits_wstrb_28 = dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@142324.4]
  assign io_dram_1_wdata_bits_wstrb_29 = dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@142325.4]
  assign io_dram_1_wdata_bits_wstrb_30 = dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@142326.4]
  assign io_dram_1_wdata_bits_wstrb_31 = dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@142327.4]
  assign io_dram_1_wdata_bits_wstrb_32 = dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@142328.4]
  assign io_dram_1_wdata_bits_wstrb_33 = dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@142329.4]
  assign io_dram_1_wdata_bits_wstrb_34 = dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@142330.4]
  assign io_dram_1_wdata_bits_wstrb_35 = dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@142331.4]
  assign io_dram_1_wdata_bits_wstrb_36 = dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@142332.4]
  assign io_dram_1_wdata_bits_wstrb_37 = dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@142333.4]
  assign io_dram_1_wdata_bits_wstrb_38 = dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@142334.4]
  assign io_dram_1_wdata_bits_wstrb_39 = dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@142335.4]
  assign io_dram_1_wdata_bits_wstrb_40 = dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@142336.4]
  assign io_dram_1_wdata_bits_wstrb_41 = dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@142337.4]
  assign io_dram_1_wdata_bits_wstrb_42 = dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@142338.4]
  assign io_dram_1_wdata_bits_wstrb_43 = dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@142339.4]
  assign io_dram_1_wdata_bits_wstrb_44 = dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@142340.4]
  assign io_dram_1_wdata_bits_wstrb_45 = dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@142341.4]
  assign io_dram_1_wdata_bits_wstrb_46 = dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@142342.4]
  assign io_dram_1_wdata_bits_wstrb_47 = dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@142343.4]
  assign io_dram_1_wdata_bits_wstrb_48 = dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@142344.4]
  assign io_dram_1_wdata_bits_wstrb_49 = dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@142345.4]
  assign io_dram_1_wdata_bits_wstrb_50 = dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@142346.4]
  assign io_dram_1_wdata_bits_wstrb_51 = dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@142347.4]
  assign io_dram_1_wdata_bits_wstrb_52 = dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@142348.4]
  assign io_dram_1_wdata_bits_wstrb_53 = dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@142349.4]
  assign io_dram_1_wdata_bits_wstrb_54 = dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@142350.4]
  assign io_dram_1_wdata_bits_wstrb_55 = dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@142351.4]
  assign io_dram_1_wdata_bits_wstrb_56 = dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@142352.4]
  assign io_dram_1_wdata_bits_wstrb_57 = dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@142353.4]
  assign io_dram_1_wdata_bits_wstrb_58 = dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@142354.4]
  assign io_dram_1_wdata_bits_wstrb_59 = dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@142355.4]
  assign io_dram_1_wdata_bits_wstrb_60 = dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@142356.4]
  assign io_dram_1_wdata_bits_wstrb_61 = dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@142357.4]
  assign io_dram_1_wdata_bits_wstrb_62 = dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@142358.4]
  assign io_dram_1_wdata_bits_wstrb_63 = dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@142359.4]
  assign io_dram_1_wdata_bits_wlast = dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@142295.4]
  assign io_dram_1_rresp_ready = dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 195:72:@142294.4]
  assign io_dram_1_wresp_ready = dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 195:72:@142275.4]
  assign io_dram_2_cmd_valid = dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 195:72:@142495.4]
  assign io_dram_2_cmd_bits_addr = dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@142494.4]
  assign io_dram_2_cmd_bits_size = dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@142493.4]
  assign io_dram_2_cmd_bits_isWr = dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@142491.4]
  assign io_dram_2_cmd_bits_tag = dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@142490.4]
  assign io_dram_2_wdata_valid = dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 195:72:@142488.4]
  assign io_dram_2_wdata_bits_wdata_0 = dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@142472.4]
  assign io_dram_2_wdata_bits_wdata_1 = dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@142473.4]
  assign io_dram_2_wdata_bits_wdata_2 = dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@142474.4]
  assign io_dram_2_wdata_bits_wdata_3 = dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@142475.4]
  assign io_dram_2_wdata_bits_wdata_4 = dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@142476.4]
  assign io_dram_2_wdata_bits_wdata_5 = dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@142477.4]
  assign io_dram_2_wdata_bits_wdata_6 = dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@142478.4]
  assign io_dram_2_wdata_bits_wdata_7 = dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@142479.4]
  assign io_dram_2_wdata_bits_wdata_8 = dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@142480.4]
  assign io_dram_2_wdata_bits_wdata_9 = dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@142481.4]
  assign io_dram_2_wdata_bits_wdata_10 = dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@142482.4]
  assign io_dram_2_wdata_bits_wdata_11 = dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@142483.4]
  assign io_dram_2_wdata_bits_wdata_12 = dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@142484.4]
  assign io_dram_2_wdata_bits_wdata_13 = dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@142485.4]
  assign io_dram_2_wdata_bits_wdata_14 = dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@142486.4]
  assign io_dram_2_wdata_bits_wdata_15 = dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@142487.4]
  assign io_dram_2_wdata_bits_wstrb_0 = dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@142408.4]
  assign io_dram_2_wdata_bits_wstrb_1 = dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@142409.4]
  assign io_dram_2_wdata_bits_wstrb_2 = dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@142410.4]
  assign io_dram_2_wdata_bits_wstrb_3 = dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@142411.4]
  assign io_dram_2_wdata_bits_wstrb_4 = dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@142412.4]
  assign io_dram_2_wdata_bits_wstrb_5 = dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@142413.4]
  assign io_dram_2_wdata_bits_wstrb_6 = dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@142414.4]
  assign io_dram_2_wdata_bits_wstrb_7 = dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@142415.4]
  assign io_dram_2_wdata_bits_wstrb_8 = dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@142416.4]
  assign io_dram_2_wdata_bits_wstrb_9 = dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@142417.4]
  assign io_dram_2_wdata_bits_wstrb_10 = dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@142418.4]
  assign io_dram_2_wdata_bits_wstrb_11 = dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@142419.4]
  assign io_dram_2_wdata_bits_wstrb_12 = dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@142420.4]
  assign io_dram_2_wdata_bits_wstrb_13 = dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@142421.4]
  assign io_dram_2_wdata_bits_wstrb_14 = dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@142422.4]
  assign io_dram_2_wdata_bits_wstrb_15 = dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@142423.4]
  assign io_dram_2_wdata_bits_wstrb_16 = dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@142424.4]
  assign io_dram_2_wdata_bits_wstrb_17 = dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@142425.4]
  assign io_dram_2_wdata_bits_wstrb_18 = dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@142426.4]
  assign io_dram_2_wdata_bits_wstrb_19 = dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@142427.4]
  assign io_dram_2_wdata_bits_wstrb_20 = dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@142428.4]
  assign io_dram_2_wdata_bits_wstrb_21 = dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@142429.4]
  assign io_dram_2_wdata_bits_wstrb_22 = dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@142430.4]
  assign io_dram_2_wdata_bits_wstrb_23 = dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@142431.4]
  assign io_dram_2_wdata_bits_wstrb_24 = dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@142432.4]
  assign io_dram_2_wdata_bits_wstrb_25 = dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@142433.4]
  assign io_dram_2_wdata_bits_wstrb_26 = dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@142434.4]
  assign io_dram_2_wdata_bits_wstrb_27 = dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@142435.4]
  assign io_dram_2_wdata_bits_wstrb_28 = dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@142436.4]
  assign io_dram_2_wdata_bits_wstrb_29 = dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@142437.4]
  assign io_dram_2_wdata_bits_wstrb_30 = dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@142438.4]
  assign io_dram_2_wdata_bits_wstrb_31 = dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@142439.4]
  assign io_dram_2_wdata_bits_wstrb_32 = dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@142440.4]
  assign io_dram_2_wdata_bits_wstrb_33 = dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@142441.4]
  assign io_dram_2_wdata_bits_wstrb_34 = dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@142442.4]
  assign io_dram_2_wdata_bits_wstrb_35 = dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@142443.4]
  assign io_dram_2_wdata_bits_wstrb_36 = dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@142444.4]
  assign io_dram_2_wdata_bits_wstrb_37 = dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@142445.4]
  assign io_dram_2_wdata_bits_wstrb_38 = dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@142446.4]
  assign io_dram_2_wdata_bits_wstrb_39 = dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@142447.4]
  assign io_dram_2_wdata_bits_wstrb_40 = dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@142448.4]
  assign io_dram_2_wdata_bits_wstrb_41 = dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@142449.4]
  assign io_dram_2_wdata_bits_wstrb_42 = dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@142450.4]
  assign io_dram_2_wdata_bits_wstrb_43 = dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@142451.4]
  assign io_dram_2_wdata_bits_wstrb_44 = dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@142452.4]
  assign io_dram_2_wdata_bits_wstrb_45 = dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@142453.4]
  assign io_dram_2_wdata_bits_wstrb_46 = dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@142454.4]
  assign io_dram_2_wdata_bits_wstrb_47 = dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@142455.4]
  assign io_dram_2_wdata_bits_wstrb_48 = dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@142456.4]
  assign io_dram_2_wdata_bits_wstrb_49 = dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@142457.4]
  assign io_dram_2_wdata_bits_wstrb_50 = dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@142458.4]
  assign io_dram_2_wdata_bits_wstrb_51 = dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@142459.4]
  assign io_dram_2_wdata_bits_wstrb_52 = dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@142460.4]
  assign io_dram_2_wdata_bits_wstrb_53 = dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@142461.4]
  assign io_dram_2_wdata_bits_wstrb_54 = dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@142462.4]
  assign io_dram_2_wdata_bits_wstrb_55 = dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@142463.4]
  assign io_dram_2_wdata_bits_wstrb_56 = dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@142464.4]
  assign io_dram_2_wdata_bits_wstrb_57 = dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@142465.4]
  assign io_dram_2_wdata_bits_wstrb_58 = dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@142466.4]
  assign io_dram_2_wdata_bits_wstrb_59 = dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@142467.4]
  assign io_dram_2_wdata_bits_wstrb_60 = dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@142468.4]
  assign io_dram_2_wdata_bits_wstrb_61 = dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@142469.4]
  assign io_dram_2_wdata_bits_wstrb_62 = dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@142470.4]
  assign io_dram_2_wdata_bits_wstrb_63 = dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@142471.4]
  assign io_dram_2_wdata_bits_wlast = dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@142407.4]
  assign io_dram_2_rresp_ready = dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 195:72:@142406.4]
  assign io_dram_2_wresp_ready = dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 195:72:@142387.4]
  assign io_dram_3_cmd_valid = dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 195:72:@142607.4]
  assign io_dram_3_cmd_bits_addr = dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@142606.4]
  assign io_dram_3_cmd_bits_size = dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@142605.4]
  assign io_dram_3_cmd_bits_isWr = dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@142603.4]
  assign io_dram_3_cmd_bits_tag = dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@142602.4]
  assign io_dram_3_wdata_valid = dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 195:72:@142600.4]
  assign io_dram_3_wdata_bits_wdata_0 = dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@142584.4]
  assign io_dram_3_wdata_bits_wdata_1 = dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@142585.4]
  assign io_dram_3_wdata_bits_wdata_2 = dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@142586.4]
  assign io_dram_3_wdata_bits_wdata_3 = dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@142587.4]
  assign io_dram_3_wdata_bits_wdata_4 = dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@142588.4]
  assign io_dram_3_wdata_bits_wdata_5 = dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@142589.4]
  assign io_dram_3_wdata_bits_wdata_6 = dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@142590.4]
  assign io_dram_3_wdata_bits_wdata_7 = dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@142591.4]
  assign io_dram_3_wdata_bits_wdata_8 = dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@142592.4]
  assign io_dram_3_wdata_bits_wdata_9 = dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@142593.4]
  assign io_dram_3_wdata_bits_wdata_10 = dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@142594.4]
  assign io_dram_3_wdata_bits_wdata_11 = dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@142595.4]
  assign io_dram_3_wdata_bits_wdata_12 = dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@142596.4]
  assign io_dram_3_wdata_bits_wdata_13 = dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@142597.4]
  assign io_dram_3_wdata_bits_wdata_14 = dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@142598.4]
  assign io_dram_3_wdata_bits_wdata_15 = dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@142599.4]
  assign io_dram_3_wdata_bits_wstrb_0 = dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@142520.4]
  assign io_dram_3_wdata_bits_wstrb_1 = dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@142521.4]
  assign io_dram_3_wdata_bits_wstrb_2 = dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@142522.4]
  assign io_dram_3_wdata_bits_wstrb_3 = dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@142523.4]
  assign io_dram_3_wdata_bits_wstrb_4 = dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@142524.4]
  assign io_dram_3_wdata_bits_wstrb_5 = dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@142525.4]
  assign io_dram_3_wdata_bits_wstrb_6 = dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@142526.4]
  assign io_dram_3_wdata_bits_wstrb_7 = dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@142527.4]
  assign io_dram_3_wdata_bits_wstrb_8 = dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@142528.4]
  assign io_dram_3_wdata_bits_wstrb_9 = dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@142529.4]
  assign io_dram_3_wdata_bits_wstrb_10 = dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@142530.4]
  assign io_dram_3_wdata_bits_wstrb_11 = dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@142531.4]
  assign io_dram_3_wdata_bits_wstrb_12 = dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@142532.4]
  assign io_dram_3_wdata_bits_wstrb_13 = dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@142533.4]
  assign io_dram_3_wdata_bits_wstrb_14 = dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@142534.4]
  assign io_dram_3_wdata_bits_wstrb_15 = dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@142535.4]
  assign io_dram_3_wdata_bits_wstrb_16 = dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@142536.4]
  assign io_dram_3_wdata_bits_wstrb_17 = dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@142537.4]
  assign io_dram_3_wdata_bits_wstrb_18 = dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@142538.4]
  assign io_dram_3_wdata_bits_wstrb_19 = dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@142539.4]
  assign io_dram_3_wdata_bits_wstrb_20 = dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@142540.4]
  assign io_dram_3_wdata_bits_wstrb_21 = dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@142541.4]
  assign io_dram_3_wdata_bits_wstrb_22 = dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@142542.4]
  assign io_dram_3_wdata_bits_wstrb_23 = dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@142543.4]
  assign io_dram_3_wdata_bits_wstrb_24 = dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@142544.4]
  assign io_dram_3_wdata_bits_wstrb_25 = dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@142545.4]
  assign io_dram_3_wdata_bits_wstrb_26 = dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@142546.4]
  assign io_dram_3_wdata_bits_wstrb_27 = dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@142547.4]
  assign io_dram_3_wdata_bits_wstrb_28 = dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@142548.4]
  assign io_dram_3_wdata_bits_wstrb_29 = dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@142549.4]
  assign io_dram_3_wdata_bits_wstrb_30 = dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@142550.4]
  assign io_dram_3_wdata_bits_wstrb_31 = dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@142551.4]
  assign io_dram_3_wdata_bits_wstrb_32 = dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@142552.4]
  assign io_dram_3_wdata_bits_wstrb_33 = dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@142553.4]
  assign io_dram_3_wdata_bits_wstrb_34 = dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@142554.4]
  assign io_dram_3_wdata_bits_wstrb_35 = dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@142555.4]
  assign io_dram_3_wdata_bits_wstrb_36 = dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@142556.4]
  assign io_dram_3_wdata_bits_wstrb_37 = dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@142557.4]
  assign io_dram_3_wdata_bits_wstrb_38 = dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@142558.4]
  assign io_dram_3_wdata_bits_wstrb_39 = dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@142559.4]
  assign io_dram_3_wdata_bits_wstrb_40 = dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@142560.4]
  assign io_dram_3_wdata_bits_wstrb_41 = dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@142561.4]
  assign io_dram_3_wdata_bits_wstrb_42 = dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@142562.4]
  assign io_dram_3_wdata_bits_wstrb_43 = dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@142563.4]
  assign io_dram_3_wdata_bits_wstrb_44 = dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@142564.4]
  assign io_dram_3_wdata_bits_wstrb_45 = dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@142565.4]
  assign io_dram_3_wdata_bits_wstrb_46 = dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@142566.4]
  assign io_dram_3_wdata_bits_wstrb_47 = dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@142567.4]
  assign io_dram_3_wdata_bits_wstrb_48 = dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@142568.4]
  assign io_dram_3_wdata_bits_wstrb_49 = dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@142569.4]
  assign io_dram_3_wdata_bits_wstrb_50 = dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@142570.4]
  assign io_dram_3_wdata_bits_wstrb_51 = dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@142571.4]
  assign io_dram_3_wdata_bits_wstrb_52 = dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@142572.4]
  assign io_dram_3_wdata_bits_wstrb_53 = dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@142573.4]
  assign io_dram_3_wdata_bits_wstrb_54 = dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@142574.4]
  assign io_dram_3_wdata_bits_wstrb_55 = dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@142575.4]
  assign io_dram_3_wdata_bits_wstrb_56 = dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@142576.4]
  assign io_dram_3_wdata_bits_wstrb_57 = dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@142577.4]
  assign io_dram_3_wdata_bits_wstrb_58 = dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@142578.4]
  assign io_dram_3_wdata_bits_wstrb_59 = dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@142579.4]
  assign io_dram_3_wdata_bits_wstrb_60 = dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@142580.4]
  assign io_dram_3_wdata_bits_wstrb_61 = dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@142581.4]
  assign io_dram_3_wdata_bits_wstrb_62 = dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@142582.4]
  assign io_dram_3_wdata_bits_wstrb_63 = dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@142583.4]
  assign io_dram_3_wdata_bits_wlast = dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@142519.4]
  assign io_dram_3_rresp_ready = dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 195:72:@142518.4]
  assign io_dram_3_wresp_ready = dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 195:72:@142499.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@139038.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@139037.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@139036.4]
  assign dramArbs_0_clock = clock; // @[:@135161.4]
  assign dramArbs_0_reset = _T_1030 | reset; // @[:@135162.4 Fringe.scala 187:30:@142153.4]
  assign dramArbs_0_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@142157.4]
  assign dramArbs_0_io_app_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[Fringe.scala 101:72:@136078.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[Fringe.scala 101:72:@136077.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[Fringe.scala 101:72:@136076.4]
  assign dramArbs_0_io_app_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[Fringe.scala 101:72:@136074.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[Fringe.scala 101:72:@136073.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[Fringe.scala 101:72:@136072.4]
  assign dramArbs_0_io_app_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[Fringe.scala 101:72:@136071.4]
  assign dramArbs_0_io_dram_cmd_ready = io_dram_0_cmd_ready; // @[Fringe.scala 195:72:@142272.4]
  assign dramArbs_0_io_dram_wdata_ready = io_dram_0_wdata_ready; // @[Fringe.scala 195:72:@142265.4]
  assign dramArbs_0_io_dram_wresp_valid = io_dram_0_wresp_valid; // @[Fringe.scala 195:72:@142162.4]
  assign dramArbs_0_io_dram_wresp_bits_tag = io_dram_0_wresp_bits_tag; // @[Fringe.scala 195:72:@142161.4]
  assign dramArbs_1_clock = clock; // @[:@136154.4]
  assign dramArbs_1_reset = _T_1030 | reset; // @[:@136155.4 Fringe.scala 187:30:@142154.4]
  assign dramArbs_1_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@142158.4]
  assign dramArbs_1_io_dram_cmd_ready = io_dram_1_cmd_ready; // @[Fringe.scala 195:72:@142384.4]
  assign dramArbs_1_io_dram_wdata_ready = io_dram_1_wdata_ready; // @[Fringe.scala 195:72:@142377.4]
  assign dramArbs_1_io_dram_wresp_valid = io_dram_1_wresp_valid; // @[Fringe.scala 195:72:@142274.4]
  assign dramArbs_1_io_dram_wresp_bits_tag = io_dram_1_wresp_bits_tag; // @[Fringe.scala 195:72:@142273.4]
  assign dramArbs_2_clock = clock; // @[:@137114.4]
  assign dramArbs_2_reset = _T_1030 | reset; // @[:@137115.4 Fringe.scala 187:30:@142155.4]
  assign dramArbs_2_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@142159.4]
  assign dramArbs_2_io_dram_cmd_ready = io_dram_2_cmd_ready; // @[Fringe.scala 195:72:@142496.4]
  assign dramArbs_2_io_dram_wdata_ready = io_dram_2_wdata_ready; // @[Fringe.scala 195:72:@142489.4]
  assign dramArbs_2_io_dram_wresp_valid = io_dram_2_wresp_valid; // @[Fringe.scala 195:72:@142386.4]
  assign dramArbs_2_io_dram_wresp_bits_tag = io_dram_2_wresp_bits_tag; // @[Fringe.scala 195:72:@142385.4]
  assign dramArbs_3_clock = clock; // @[:@138074.4]
  assign dramArbs_3_reset = _T_1030 | reset; // @[:@138075.4 Fringe.scala 187:30:@142156.4]
  assign dramArbs_3_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@142160.4]
  assign dramArbs_3_io_dram_cmd_ready = io_dram_3_cmd_ready; // @[Fringe.scala 195:72:@142608.4]
  assign dramArbs_3_io_dram_wdata_ready = io_dram_3_wdata_ready; // @[Fringe.scala 195:72:@142601.4]
  assign dramArbs_3_io_dram_wresp_valid = io_dram_3_wresp_valid; // @[Fringe.scala 195:72:@142498.4]
  assign dramArbs_3_io_dram_wresp_bits_tag = io_dram_3_wresp_bits_tag; // @[Fringe.scala 195:72:@142497.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@139041.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@139040.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@139039.4]
  assign heap_io_host_0_resp_valid = _T_1569 & _T_1573; // @[Fringe.scala 204:22:@142780.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@142781.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@142782.4]
  assign regs_clock = clock; // @[:@139043.4]
  assign regs_reset = reset; // @[:@139044.4 Fringe.scala 139:14:@141091.4]
  assign regs_io_raddr = io_raddr; // @[Fringe.scala 118:17:@141063.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@141065.4]
  assign regs_io_waddr = io_waddr; // @[Fringe.scala 119:17:@141064.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@141066.4]
  assign regs_io_reset = _T_1030 | reset; // @[Fringe.scala 138:17:@141089.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_1049; // @[Fringe.scala 170:23:@141141.4]
  assign regs_io_argOuts_0_bits = {_T_1065,_T_1064}; // @[Fringe.scala 171:22:@141145.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@141148.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@141147.4]
  assign timeoutCtr_clock = clock; // @[:@141093.4]
  assign timeoutCtr_reset = reset; // @[:@141094.4]
  assign timeoutCtr_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 149:24:@141108.4]
  assign depulser_clock = clock; // @[:@141112.4]
  assign depulser_reset = reset; // @[:@141113.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@141118.4]
  assign depulser_io_rst = _T_1040[0]; // @[Fringe.scala 156:19:@141120.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1047 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1572 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1047 <= 1'h0;
    end else begin
      _T_1047 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1572 <= 1'h0;
    end else begin
      _T_1572 <= _T_1569;
    end
  end
endmodule
module AXI4LiteToRFBridge( // @[:@142797.2]
  input         clock, // @[:@142798.4]
  input         reset, // @[:@142799.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@142800.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@142800.4]
  input         io_S_AXI_AWVALID, // @[:@142800.4]
  output        io_S_AXI_AWREADY, // @[:@142800.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@142800.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@142800.4]
  input         io_S_AXI_ARVALID, // @[:@142800.4]
  output        io_S_AXI_ARREADY, // @[:@142800.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@142800.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@142800.4]
  input         io_S_AXI_WVALID, // @[:@142800.4]
  output        io_S_AXI_WREADY, // @[:@142800.4]
  output [31:0] io_S_AXI_RDATA, // @[:@142800.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@142800.4]
  output        io_S_AXI_RVALID, // @[:@142800.4]
  input         io_S_AXI_RREADY, // @[:@142800.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@142800.4]
  output        io_S_AXI_BVALID, // @[:@142800.4]
  input         io_S_AXI_BREADY, // @[:@142800.4]
  output [31:0] io_raddr, // @[:@142800.4]
  output        io_wen, // @[:@142800.4]
  output [31:0] io_waddr, // @[:@142800.4]
  output [31:0] io_wdata, // @[:@142800.4]
  input  [31:0] io_rdata // @[:@142800.4]
);
  wire [31:0] d_rf_rdata; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire [31:0] d_rf_wdata; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire [31:0] d_rf_waddr; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire  d_rf_wen; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire [31:0] d_rf_raddr; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire  d_S_AXI_ARESETN; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire  d_S_AXI_ACLK; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire [31:0] d_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire [2:0] d_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire  d_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire  d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire [31:0] d_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire [2:0] d_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire  d_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire  d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire [31:0] d_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire [3:0] d_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire  d_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire  d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire [31:0] d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire [1:0] d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire  d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire  d_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire [1:0] d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire  d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  wire  d_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
  AXI4LiteToRFBridgeVerilog d ( // @[AXI4LiteToRFBridge.scala 36:17:@142802.4]
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 38:14:@142826.4]
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 38:14:@142822.4]
  assign io_S_AXI_WREADY = d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 38:14:@142818.4]
  assign io_S_AXI_RDATA = d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 38:14:@142817.4]
  assign io_S_AXI_RRESP = d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 38:14:@142816.4]
  assign io_S_AXI_RVALID = d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 38:14:@142815.4]
  assign io_S_AXI_BRESP = d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 38:14:@142813.4]
  assign io_S_AXI_BVALID = d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 38:14:@142812.4]
  assign io_raddr = d_rf_raddr; // @[AXI4LiteToRFBridge.scala 42:12:@142834.4]
  assign io_wen = d_rf_wen; // @[AXI4LiteToRFBridge.scala 45:12:@142837.4]
  assign io_waddr = d_rf_waddr; // @[AXI4LiteToRFBridge.scala 43:12:@142835.4]
  assign io_wdata = d_rf_wdata; // @[AXI4LiteToRFBridge.scala 44:12:@142836.4]
  assign d_rf_rdata = io_rdata; // @[AXI4LiteToRFBridge.scala 46:17:@142838.4]
  assign d_S_AXI_ARESETN = ~ reset; // @[AXI4LiteToRFBridge.scala 40:22:@142833.4]
  assign d_S_AXI_ACLK = clock; // @[AXI4LiteToRFBridge.scala 39:19:@142830.4]
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 38:14:@142829.4]
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 38:14:@142828.4]
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 38:14:@142827.4]
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 38:14:@142825.4]
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 38:14:@142824.4]
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 38:14:@142823.4]
  assign d_S_AXI_WDATA = io_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 38:14:@142821.4]
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 38:14:@142820.4]
  assign d_S_AXI_WVALID = io_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 38:14:@142819.4]
  assign d_S_AXI_RREADY = io_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 38:14:@142814.4]
  assign d_S_AXI_BREADY = io_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 38:14:@142811.4]
endmodule
module MAGToAXI4Bridge( // @[:@142840.2]
  output         io_in_cmd_ready, // @[:@142843.4]
  input          io_in_cmd_valid, // @[:@142843.4]
  input  [63:0]  io_in_cmd_bits_addr, // @[:@142843.4]
  input  [31:0]  io_in_cmd_bits_size, // @[:@142843.4]
  input          io_in_cmd_bits_isWr, // @[:@142843.4]
  input  [31:0]  io_in_cmd_bits_tag, // @[:@142843.4]
  output         io_in_wdata_ready, // @[:@142843.4]
  input          io_in_wdata_valid, // @[:@142843.4]
  input  [31:0]  io_in_wdata_bits_wdata_0, // @[:@142843.4]
  input  [31:0]  io_in_wdata_bits_wdata_1, // @[:@142843.4]
  input  [31:0]  io_in_wdata_bits_wdata_2, // @[:@142843.4]
  input  [31:0]  io_in_wdata_bits_wdata_3, // @[:@142843.4]
  input  [31:0]  io_in_wdata_bits_wdata_4, // @[:@142843.4]
  input  [31:0]  io_in_wdata_bits_wdata_5, // @[:@142843.4]
  input  [31:0]  io_in_wdata_bits_wdata_6, // @[:@142843.4]
  input  [31:0]  io_in_wdata_bits_wdata_7, // @[:@142843.4]
  input  [31:0]  io_in_wdata_bits_wdata_8, // @[:@142843.4]
  input  [31:0]  io_in_wdata_bits_wdata_9, // @[:@142843.4]
  input  [31:0]  io_in_wdata_bits_wdata_10, // @[:@142843.4]
  input  [31:0]  io_in_wdata_bits_wdata_11, // @[:@142843.4]
  input  [31:0]  io_in_wdata_bits_wdata_12, // @[:@142843.4]
  input  [31:0]  io_in_wdata_bits_wdata_13, // @[:@142843.4]
  input  [31:0]  io_in_wdata_bits_wdata_14, // @[:@142843.4]
  input  [31:0]  io_in_wdata_bits_wdata_15, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_0, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_1, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_2, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_3, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_4, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_5, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_6, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_7, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_8, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_9, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_10, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_11, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_12, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_13, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_14, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_15, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_16, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_17, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_18, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_19, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_20, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_21, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_22, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_23, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_24, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_25, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_26, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_27, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_28, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_29, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_30, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_31, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_32, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_33, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_34, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_35, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_36, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_37, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_38, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_39, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_40, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_41, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_42, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_43, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_44, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_45, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_46, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_47, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_48, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_49, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_50, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_51, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_52, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_53, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_54, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_55, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_56, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_57, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_58, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_59, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_60, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_61, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_62, // @[:@142843.4]
  input          io_in_wdata_bits_wstrb_63, // @[:@142843.4]
  input          io_in_wdata_bits_wlast, // @[:@142843.4]
  input          io_in_rresp_ready, // @[:@142843.4]
  input          io_in_wresp_ready, // @[:@142843.4]
  output         io_in_wresp_valid, // @[:@142843.4]
  output [31:0]  io_in_wresp_bits_tag, // @[:@142843.4]
  output [31:0]  io_M_AXI_AWID, // @[:@142843.4]
  output [31:0]  io_M_AXI_AWADDR, // @[:@142843.4]
  output [7:0]   io_M_AXI_AWLEN, // @[:@142843.4]
  output         io_M_AXI_AWVALID, // @[:@142843.4]
  input          io_M_AXI_AWREADY, // @[:@142843.4]
  output [31:0]  io_M_AXI_ARID, // @[:@142843.4]
  output [31:0]  io_M_AXI_ARADDR, // @[:@142843.4]
  output [7:0]   io_M_AXI_ARLEN, // @[:@142843.4]
  output         io_M_AXI_ARVALID, // @[:@142843.4]
  input          io_M_AXI_ARREADY, // @[:@142843.4]
  output [511:0] io_M_AXI_WDATA, // @[:@142843.4]
  output [63:0]  io_M_AXI_WSTRB, // @[:@142843.4]
  output         io_M_AXI_WLAST, // @[:@142843.4]
  output         io_M_AXI_WVALID, // @[:@142843.4]
  input          io_M_AXI_WREADY, // @[:@142843.4]
  output         io_M_AXI_RREADY, // @[:@142843.4]
  input  [31:0]  io_M_AXI_BID, // @[:@142843.4]
  input          io_M_AXI_BVALID, // @[:@142843.4]
  output         io_M_AXI_BREADY // @[:@142843.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@143000.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@143001.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@143002.4]
  wire  _T_228; // @[MAGToAXI4Bridge.scala 35:42:@143010.4]
  wire [319:0] _T_250; // @[Cat.scala 30:58:@143037.4]
  wire [479:0] _T_255; // @[Cat.scala 30:58:@143042.4]
  wire [9:0] _T_265; // @[Cat.scala 30:58:@143053.4]
  wire [18:0] _T_274; // @[Cat.scala 30:58:@143062.4]
  wire [27:0] _T_283; // @[Cat.scala 30:58:@143071.4]
  wire [36:0] _T_292; // @[Cat.scala 30:58:@143080.4]
  wire [45:0] _T_301; // @[Cat.scala 30:58:@143089.4]
  wire [54:0] _T_310; // @[Cat.scala 30:58:@143098.4]
  wire [62:0] _T_318; // @[Cat.scala 30:58:@143106.4]
  assign _T_218 = io_in_cmd_bits_size - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@143000.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@143001.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@143002.4]
  assign _T_228 = io_in_cmd_bits_isWr == 1'h0; // @[MAGToAXI4Bridge.scala 35:42:@143010.4]
  assign _T_250 = {io_in_wdata_bits_wdata_15,io_in_wdata_bits_wdata_14,io_in_wdata_bits_wdata_13,io_in_wdata_bits_wdata_12,io_in_wdata_bits_wdata_11,io_in_wdata_bits_wdata_10,io_in_wdata_bits_wdata_9,io_in_wdata_bits_wdata_8,io_in_wdata_bits_wdata_7,io_in_wdata_bits_wdata_6}; // @[Cat.scala 30:58:@143037.4]
  assign _T_255 = {_T_250,io_in_wdata_bits_wdata_5,io_in_wdata_bits_wdata_4,io_in_wdata_bits_wdata_3,io_in_wdata_bits_wdata_2,io_in_wdata_bits_wdata_1}; // @[Cat.scala 30:58:@143042.4]
  assign _T_265 = {io_in_wdata_bits_wstrb_63,io_in_wdata_bits_wstrb_62,io_in_wdata_bits_wstrb_61,io_in_wdata_bits_wstrb_60,io_in_wdata_bits_wstrb_59,io_in_wdata_bits_wstrb_58,io_in_wdata_bits_wstrb_57,io_in_wdata_bits_wstrb_56,io_in_wdata_bits_wstrb_55,io_in_wdata_bits_wstrb_54}; // @[Cat.scala 30:58:@143053.4]
  assign _T_274 = {_T_265,io_in_wdata_bits_wstrb_53,io_in_wdata_bits_wstrb_52,io_in_wdata_bits_wstrb_51,io_in_wdata_bits_wstrb_50,io_in_wdata_bits_wstrb_49,io_in_wdata_bits_wstrb_48,io_in_wdata_bits_wstrb_47,io_in_wdata_bits_wstrb_46,io_in_wdata_bits_wstrb_45}; // @[Cat.scala 30:58:@143062.4]
  assign _T_283 = {_T_274,io_in_wdata_bits_wstrb_44,io_in_wdata_bits_wstrb_43,io_in_wdata_bits_wstrb_42,io_in_wdata_bits_wstrb_41,io_in_wdata_bits_wstrb_40,io_in_wdata_bits_wstrb_39,io_in_wdata_bits_wstrb_38,io_in_wdata_bits_wstrb_37,io_in_wdata_bits_wstrb_36}; // @[Cat.scala 30:58:@143071.4]
  assign _T_292 = {_T_283,io_in_wdata_bits_wstrb_35,io_in_wdata_bits_wstrb_34,io_in_wdata_bits_wstrb_33,io_in_wdata_bits_wstrb_32,io_in_wdata_bits_wstrb_31,io_in_wdata_bits_wstrb_30,io_in_wdata_bits_wstrb_29,io_in_wdata_bits_wstrb_28,io_in_wdata_bits_wstrb_27}; // @[Cat.scala 30:58:@143080.4]
  assign _T_301 = {_T_292,io_in_wdata_bits_wstrb_26,io_in_wdata_bits_wstrb_25,io_in_wdata_bits_wstrb_24,io_in_wdata_bits_wstrb_23,io_in_wdata_bits_wstrb_22,io_in_wdata_bits_wstrb_21,io_in_wdata_bits_wstrb_20,io_in_wdata_bits_wstrb_19,io_in_wdata_bits_wstrb_18}; // @[Cat.scala 30:58:@143089.4]
  assign _T_310 = {_T_301,io_in_wdata_bits_wstrb_17,io_in_wdata_bits_wstrb_16,io_in_wdata_bits_wstrb_15,io_in_wdata_bits_wstrb_14,io_in_wdata_bits_wstrb_13,io_in_wdata_bits_wstrb_12,io_in_wdata_bits_wstrb_11,io_in_wdata_bits_wstrb_10,io_in_wdata_bits_wstrb_9}; // @[Cat.scala 30:58:@143098.4]
  assign _T_318 = {_T_310,io_in_wdata_bits_wstrb_8,io_in_wdata_bits_wstrb_7,io_in_wdata_bits_wstrb_6,io_in_wdata_bits_wstrb_5,io_in_wdata_bits_wstrb_4,io_in_wdata_bits_wstrb_3,io_in_wdata_bits_wstrb_2,io_in_wdata_bits_wstrb_1}; // @[Cat.scala 30:58:@143106.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? io_M_AXI_AWREADY : io_M_AXI_ARREADY; // @[MAGToAXI4Bridge.scala 36:21:@143014.4]
  assign io_in_wdata_ready = io_M_AXI_WREADY; // @[MAGToAXI4Bridge.scala 56:21:@143111.4]
  assign io_in_wresp_valid = io_M_AXI_BVALID; // @[MAGToAXI4Bridge.scala 71:21:@143164.4]
  assign io_in_wresp_bits_tag = io_M_AXI_BID; // @[MAGToAXI4Bridge.scala 74:24:@143166.4]
  assign io_M_AXI_AWID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 39:21:@143015.4]
  assign io_M_AXI_AWADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 40:21:@143016.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@143020.4]
  assign io_M_AXI_AWVALID = io_in_cmd_valid & io_in_cmd_bits_isWr; // @[MAGToAXI4Bridge.scala 49:21:@143028.4]
  assign io_M_AXI_ARID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 25:21:@142998.4]
  assign io_M_AXI_ARADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 26:21:@142999.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@143003.4]
  assign io_M_AXI_ARVALID = io_in_cmd_valid & _T_228; // @[MAGToAXI4Bridge.scala 35:21:@143012.4]
  assign io_M_AXI_WDATA = {_T_255,io_in_wdata_bits_wdata_0}; // @[MAGToAXI4Bridge.scala 52:21:@143044.4]
  assign io_M_AXI_WSTRB = {_T_318,io_in_wdata_bits_wstrb_0}; // @[MAGToAXI4Bridge.scala 53:21:@143108.4]
  assign io_M_AXI_WLAST = io_in_wdata_bits_wlast; // @[MAGToAXI4Bridge.scala 54:21:@143109.4]
  assign io_M_AXI_WVALID = io_in_wdata_valid; // @[MAGToAXI4Bridge.scala 55:21:@143110.4]
  assign io_M_AXI_RREADY = io_in_rresp_ready; // @[MAGToAXI4Bridge.scala 64:19:@143161.4]
  assign io_M_AXI_BREADY = io_in_wresp_ready; // @[MAGToAXI4Bridge.scala 67:19:@143162.4]
endmodule
module FringeZynq( // @[:@144152.2]
  input          clock, // @[:@144153.4]
  input          reset, // @[:@144154.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@144155.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@144155.4]
  input          io_S_AXI_AWVALID, // @[:@144155.4]
  output         io_S_AXI_AWREADY, // @[:@144155.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@144155.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@144155.4]
  input          io_S_AXI_ARVALID, // @[:@144155.4]
  output         io_S_AXI_ARREADY, // @[:@144155.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@144155.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@144155.4]
  input          io_S_AXI_WVALID, // @[:@144155.4]
  output         io_S_AXI_WREADY, // @[:@144155.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@144155.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@144155.4]
  output         io_S_AXI_RVALID, // @[:@144155.4]
  input          io_S_AXI_RREADY, // @[:@144155.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@144155.4]
  output         io_S_AXI_BVALID, // @[:@144155.4]
  input          io_S_AXI_BREADY, // @[:@144155.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@144155.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@144155.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@144155.4]
  output         io_M_AXI_0_AWVALID, // @[:@144155.4]
  input          io_M_AXI_0_AWREADY, // @[:@144155.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@144155.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@144155.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@144155.4]
  output         io_M_AXI_0_ARVALID, // @[:@144155.4]
  input          io_M_AXI_0_ARREADY, // @[:@144155.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@144155.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@144155.4]
  output         io_M_AXI_0_WLAST, // @[:@144155.4]
  output         io_M_AXI_0_WVALID, // @[:@144155.4]
  input          io_M_AXI_0_WREADY, // @[:@144155.4]
  output         io_M_AXI_0_RREADY, // @[:@144155.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@144155.4]
  input          io_M_AXI_0_BVALID, // @[:@144155.4]
  output         io_M_AXI_0_BREADY, // @[:@144155.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@144155.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@144155.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@144155.4]
  output         io_M_AXI_1_AWVALID, // @[:@144155.4]
  input          io_M_AXI_1_AWREADY, // @[:@144155.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@144155.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@144155.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@144155.4]
  output         io_M_AXI_1_ARVALID, // @[:@144155.4]
  input          io_M_AXI_1_ARREADY, // @[:@144155.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@144155.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@144155.4]
  output         io_M_AXI_1_WLAST, // @[:@144155.4]
  output         io_M_AXI_1_WVALID, // @[:@144155.4]
  input          io_M_AXI_1_WREADY, // @[:@144155.4]
  output         io_M_AXI_1_RREADY, // @[:@144155.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@144155.4]
  input          io_M_AXI_1_BVALID, // @[:@144155.4]
  output         io_M_AXI_1_BREADY, // @[:@144155.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@144155.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@144155.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@144155.4]
  output         io_M_AXI_2_AWVALID, // @[:@144155.4]
  input          io_M_AXI_2_AWREADY, // @[:@144155.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@144155.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@144155.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@144155.4]
  output         io_M_AXI_2_ARVALID, // @[:@144155.4]
  input          io_M_AXI_2_ARREADY, // @[:@144155.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@144155.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@144155.4]
  output         io_M_AXI_2_WLAST, // @[:@144155.4]
  output         io_M_AXI_2_WVALID, // @[:@144155.4]
  input          io_M_AXI_2_WREADY, // @[:@144155.4]
  output         io_M_AXI_2_RREADY, // @[:@144155.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@144155.4]
  input          io_M_AXI_2_BVALID, // @[:@144155.4]
  output         io_M_AXI_2_BREADY, // @[:@144155.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@144155.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@144155.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@144155.4]
  output         io_M_AXI_3_AWVALID, // @[:@144155.4]
  input          io_M_AXI_3_AWREADY, // @[:@144155.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@144155.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@144155.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@144155.4]
  output         io_M_AXI_3_ARVALID, // @[:@144155.4]
  input          io_M_AXI_3_ARREADY, // @[:@144155.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@144155.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@144155.4]
  output         io_M_AXI_3_WLAST, // @[:@144155.4]
  output         io_M_AXI_3_WVALID, // @[:@144155.4]
  input          io_M_AXI_3_WREADY, // @[:@144155.4]
  output         io_M_AXI_3_RREADY, // @[:@144155.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@144155.4]
  input          io_M_AXI_3_BVALID, // @[:@144155.4]
  output         io_M_AXI_3_BREADY, // @[:@144155.4]
  output         io_enable, // @[:@144155.4]
  input          io_done, // @[:@144155.4]
  output         io_reset, // @[:@144155.4]
  output [63:0]  io_argIns_0, // @[:@144155.4]
  output [63:0]  io_argIns_1, // @[:@144155.4]
  input          io_argOuts_0_valid, // @[:@144155.4]
  input  [63:0]  io_argOuts_0_bits, // @[:@144155.4]
  output         io_memStreams_stores_0_cmd_ready, // @[:@144155.4]
  input          io_memStreams_stores_0_cmd_valid, // @[:@144155.4]
  input  [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@144155.4]
  input  [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@144155.4]
  output         io_memStreams_stores_0_data_ready, // @[:@144155.4]
  input          io_memStreams_stores_0_data_valid, // @[:@144155.4]
  input  [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@144155.4]
  input          io_memStreams_stores_0_data_bits_wstrb, // @[:@144155.4]
  input          io_memStreams_stores_0_wresp_ready, // @[:@144155.4]
  output         io_memStreams_stores_0_wresp_valid, // @[:@144155.4]
  output         io_memStreams_stores_0_wresp_bits, // @[:@144155.4]
  input          io_heap_0_req_valid, // @[:@144155.4]
  input          io_heap_0_req_bits_allocDealloc, // @[:@144155.4]
  input  [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@144155.4]
  output         io_heap_0_resp_valid, // @[:@144155.4]
  output         io_heap_0_resp_bits_allocDealloc, // @[:@144155.4]
  output [63:0]  io_heap_0_resp_bits_sizeAddr // @[:@144155.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_raddr; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_wen; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_waddr; // @[FringeZynq.scala 69:28:@144626.4]
  wire [63:0] fringeCommon_io_wdata; // @[FringeZynq.scala 69:28:@144626.4]
  wire [63:0] fringeCommon_io_rdata; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 69:28:@144626.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 69:28:@144626.4]
  wire [63:0] fringeCommon_io_argIns_1; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 69:28:@144626.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 69:28:@144626.4]
  wire [63:0] fringeCommon_io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_cmd_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 69:28:@144626.4]
  wire [63:0] fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_0_wresp_valid; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_0_wresp_bits_tag; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_cmd_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 69:28:@144626.4]
  wire [63:0] fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_1_wresp_valid; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_1_wresp_bits_tag; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_cmd_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 69:28:@144626.4]
  wire [63:0] fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_2_wresp_valid; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_2_wresp_bits_tag; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_cmd_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 69:28:@144626.4]
  wire [63:0] fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_dram_3_wresp_valid; // @[FringeZynq.scala 69:28:@144626.4]
  wire [31:0] fringeCommon_io_dram_3_wresp_bits_tag; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_heap_0_req_valid; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 69:28:@144626.4]
  wire [63:0] fringeCommon_io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 69:28:@144626.4]
  wire  fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 69:28:@144626.4]
  wire [63:0] fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 69:28:@144626.4]
  wire  AXI4LiteToRFBridge_clock; // @[FringeZynq.scala 90:31:@145532.4]
  wire  AXI4LiteToRFBridge_reset; // @[FringeZynq.scala 90:31:@145532.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_AWADDR; // @[FringeZynq.scala 90:31:@145532.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_AWPROT; // @[FringeZynq.scala 90:31:@145532.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWVALID; // @[FringeZynq.scala 90:31:@145532.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 90:31:@145532.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_ARADDR; // @[FringeZynq.scala 90:31:@145532.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_ARPROT; // @[FringeZynq.scala 90:31:@145532.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARVALID; // @[FringeZynq.scala 90:31:@145532.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 90:31:@145532.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_WDATA; // @[FringeZynq.scala 90:31:@145532.4]
  wire [3:0] AXI4LiteToRFBridge_io_S_AXI_WSTRB; // @[FringeZynq.scala 90:31:@145532.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WVALID; // @[FringeZynq.scala 90:31:@145532.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 90:31:@145532.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 90:31:@145532.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 90:31:@145532.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 90:31:@145532.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RREADY; // @[FringeZynq.scala 90:31:@145532.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 90:31:@145532.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 90:31:@145532.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BREADY; // @[FringeZynq.scala 90:31:@145532.4]
  wire [31:0] AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 90:31:@145532.4]
  wire  AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 90:31:@145532.4]
  wire [31:0] AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 90:31:@145532.4]
  wire [31:0] AXI4LiteToRFBridge_io_wdata; // @[FringeZynq.scala 90:31:@145532.4]
  wire [31:0] AXI4LiteToRFBridge_io_rdata; // @[FringeZynq.scala 90:31:@145532.4]
  wire  MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@145682.4]
  wire [63:0] MAGToAXI4Bridge_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@145682.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@145682.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@145682.4]
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@145682.4]
  wire [63:0] MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@145682.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@145682.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@145838.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@145838.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@145838.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@145838.4]
  wire [511:0] MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@145838.4]
  wire [63:0] MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@145838.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@145838.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@145994.4]
  wire [63:0] MAGToAXI4Bridge_2_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@145994.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@145994.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@145994.4]
  wire [511:0] MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@145994.4]
  wire [63:0] MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@145994.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@145994.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@146150.4]
  wire [63:0] MAGToAXI4Bridge_3_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@146150.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@146150.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@146150.4]
  wire [511:0] MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@146150.4]
  wire [63:0] MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@146150.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@146150.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@146150.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 69:28:@144626.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argIns_1(fringeCommon_io_argIns_1),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(fringeCommon_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(fringeCommon_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(fringeCommon_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(fringeCommon_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(fringeCommon_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(fringeCommon_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(fringeCommon_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(fringeCommon_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(fringeCommon_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(fringeCommon_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(fringeCommon_io_memStreams_stores_0_wresp_bits),
    .io_dram_0_cmd_ready(fringeCommon_io_dram_0_cmd_ready),
    .io_dram_0_cmd_valid(fringeCommon_io_dram_0_cmd_valid),
    .io_dram_0_cmd_bits_addr(fringeCommon_io_dram_0_cmd_bits_addr),
    .io_dram_0_cmd_bits_size(fringeCommon_io_dram_0_cmd_bits_size),
    .io_dram_0_cmd_bits_isWr(fringeCommon_io_dram_0_cmd_bits_isWr),
    .io_dram_0_cmd_bits_tag(fringeCommon_io_dram_0_cmd_bits_tag),
    .io_dram_0_wdata_ready(fringeCommon_io_dram_0_wdata_ready),
    .io_dram_0_wdata_valid(fringeCommon_io_dram_0_wdata_valid),
    .io_dram_0_wdata_bits_wdata_0(fringeCommon_io_dram_0_wdata_bits_wdata_0),
    .io_dram_0_wdata_bits_wdata_1(fringeCommon_io_dram_0_wdata_bits_wdata_1),
    .io_dram_0_wdata_bits_wdata_2(fringeCommon_io_dram_0_wdata_bits_wdata_2),
    .io_dram_0_wdata_bits_wdata_3(fringeCommon_io_dram_0_wdata_bits_wdata_3),
    .io_dram_0_wdata_bits_wdata_4(fringeCommon_io_dram_0_wdata_bits_wdata_4),
    .io_dram_0_wdata_bits_wdata_5(fringeCommon_io_dram_0_wdata_bits_wdata_5),
    .io_dram_0_wdata_bits_wdata_6(fringeCommon_io_dram_0_wdata_bits_wdata_6),
    .io_dram_0_wdata_bits_wdata_7(fringeCommon_io_dram_0_wdata_bits_wdata_7),
    .io_dram_0_wdata_bits_wdata_8(fringeCommon_io_dram_0_wdata_bits_wdata_8),
    .io_dram_0_wdata_bits_wdata_9(fringeCommon_io_dram_0_wdata_bits_wdata_9),
    .io_dram_0_wdata_bits_wdata_10(fringeCommon_io_dram_0_wdata_bits_wdata_10),
    .io_dram_0_wdata_bits_wdata_11(fringeCommon_io_dram_0_wdata_bits_wdata_11),
    .io_dram_0_wdata_bits_wdata_12(fringeCommon_io_dram_0_wdata_bits_wdata_12),
    .io_dram_0_wdata_bits_wdata_13(fringeCommon_io_dram_0_wdata_bits_wdata_13),
    .io_dram_0_wdata_bits_wdata_14(fringeCommon_io_dram_0_wdata_bits_wdata_14),
    .io_dram_0_wdata_bits_wdata_15(fringeCommon_io_dram_0_wdata_bits_wdata_15),
    .io_dram_0_wdata_bits_wstrb_0(fringeCommon_io_dram_0_wdata_bits_wstrb_0),
    .io_dram_0_wdata_bits_wstrb_1(fringeCommon_io_dram_0_wdata_bits_wstrb_1),
    .io_dram_0_wdata_bits_wstrb_2(fringeCommon_io_dram_0_wdata_bits_wstrb_2),
    .io_dram_0_wdata_bits_wstrb_3(fringeCommon_io_dram_0_wdata_bits_wstrb_3),
    .io_dram_0_wdata_bits_wstrb_4(fringeCommon_io_dram_0_wdata_bits_wstrb_4),
    .io_dram_0_wdata_bits_wstrb_5(fringeCommon_io_dram_0_wdata_bits_wstrb_5),
    .io_dram_0_wdata_bits_wstrb_6(fringeCommon_io_dram_0_wdata_bits_wstrb_6),
    .io_dram_0_wdata_bits_wstrb_7(fringeCommon_io_dram_0_wdata_bits_wstrb_7),
    .io_dram_0_wdata_bits_wstrb_8(fringeCommon_io_dram_0_wdata_bits_wstrb_8),
    .io_dram_0_wdata_bits_wstrb_9(fringeCommon_io_dram_0_wdata_bits_wstrb_9),
    .io_dram_0_wdata_bits_wstrb_10(fringeCommon_io_dram_0_wdata_bits_wstrb_10),
    .io_dram_0_wdata_bits_wstrb_11(fringeCommon_io_dram_0_wdata_bits_wstrb_11),
    .io_dram_0_wdata_bits_wstrb_12(fringeCommon_io_dram_0_wdata_bits_wstrb_12),
    .io_dram_0_wdata_bits_wstrb_13(fringeCommon_io_dram_0_wdata_bits_wstrb_13),
    .io_dram_0_wdata_bits_wstrb_14(fringeCommon_io_dram_0_wdata_bits_wstrb_14),
    .io_dram_0_wdata_bits_wstrb_15(fringeCommon_io_dram_0_wdata_bits_wstrb_15),
    .io_dram_0_wdata_bits_wstrb_16(fringeCommon_io_dram_0_wdata_bits_wstrb_16),
    .io_dram_0_wdata_bits_wstrb_17(fringeCommon_io_dram_0_wdata_bits_wstrb_17),
    .io_dram_0_wdata_bits_wstrb_18(fringeCommon_io_dram_0_wdata_bits_wstrb_18),
    .io_dram_0_wdata_bits_wstrb_19(fringeCommon_io_dram_0_wdata_bits_wstrb_19),
    .io_dram_0_wdata_bits_wstrb_20(fringeCommon_io_dram_0_wdata_bits_wstrb_20),
    .io_dram_0_wdata_bits_wstrb_21(fringeCommon_io_dram_0_wdata_bits_wstrb_21),
    .io_dram_0_wdata_bits_wstrb_22(fringeCommon_io_dram_0_wdata_bits_wstrb_22),
    .io_dram_0_wdata_bits_wstrb_23(fringeCommon_io_dram_0_wdata_bits_wstrb_23),
    .io_dram_0_wdata_bits_wstrb_24(fringeCommon_io_dram_0_wdata_bits_wstrb_24),
    .io_dram_0_wdata_bits_wstrb_25(fringeCommon_io_dram_0_wdata_bits_wstrb_25),
    .io_dram_0_wdata_bits_wstrb_26(fringeCommon_io_dram_0_wdata_bits_wstrb_26),
    .io_dram_0_wdata_bits_wstrb_27(fringeCommon_io_dram_0_wdata_bits_wstrb_27),
    .io_dram_0_wdata_bits_wstrb_28(fringeCommon_io_dram_0_wdata_bits_wstrb_28),
    .io_dram_0_wdata_bits_wstrb_29(fringeCommon_io_dram_0_wdata_bits_wstrb_29),
    .io_dram_0_wdata_bits_wstrb_30(fringeCommon_io_dram_0_wdata_bits_wstrb_30),
    .io_dram_0_wdata_bits_wstrb_31(fringeCommon_io_dram_0_wdata_bits_wstrb_31),
    .io_dram_0_wdata_bits_wstrb_32(fringeCommon_io_dram_0_wdata_bits_wstrb_32),
    .io_dram_0_wdata_bits_wstrb_33(fringeCommon_io_dram_0_wdata_bits_wstrb_33),
    .io_dram_0_wdata_bits_wstrb_34(fringeCommon_io_dram_0_wdata_bits_wstrb_34),
    .io_dram_0_wdata_bits_wstrb_35(fringeCommon_io_dram_0_wdata_bits_wstrb_35),
    .io_dram_0_wdata_bits_wstrb_36(fringeCommon_io_dram_0_wdata_bits_wstrb_36),
    .io_dram_0_wdata_bits_wstrb_37(fringeCommon_io_dram_0_wdata_bits_wstrb_37),
    .io_dram_0_wdata_bits_wstrb_38(fringeCommon_io_dram_0_wdata_bits_wstrb_38),
    .io_dram_0_wdata_bits_wstrb_39(fringeCommon_io_dram_0_wdata_bits_wstrb_39),
    .io_dram_0_wdata_bits_wstrb_40(fringeCommon_io_dram_0_wdata_bits_wstrb_40),
    .io_dram_0_wdata_bits_wstrb_41(fringeCommon_io_dram_0_wdata_bits_wstrb_41),
    .io_dram_0_wdata_bits_wstrb_42(fringeCommon_io_dram_0_wdata_bits_wstrb_42),
    .io_dram_0_wdata_bits_wstrb_43(fringeCommon_io_dram_0_wdata_bits_wstrb_43),
    .io_dram_0_wdata_bits_wstrb_44(fringeCommon_io_dram_0_wdata_bits_wstrb_44),
    .io_dram_0_wdata_bits_wstrb_45(fringeCommon_io_dram_0_wdata_bits_wstrb_45),
    .io_dram_0_wdata_bits_wstrb_46(fringeCommon_io_dram_0_wdata_bits_wstrb_46),
    .io_dram_0_wdata_bits_wstrb_47(fringeCommon_io_dram_0_wdata_bits_wstrb_47),
    .io_dram_0_wdata_bits_wstrb_48(fringeCommon_io_dram_0_wdata_bits_wstrb_48),
    .io_dram_0_wdata_bits_wstrb_49(fringeCommon_io_dram_0_wdata_bits_wstrb_49),
    .io_dram_0_wdata_bits_wstrb_50(fringeCommon_io_dram_0_wdata_bits_wstrb_50),
    .io_dram_0_wdata_bits_wstrb_51(fringeCommon_io_dram_0_wdata_bits_wstrb_51),
    .io_dram_0_wdata_bits_wstrb_52(fringeCommon_io_dram_0_wdata_bits_wstrb_52),
    .io_dram_0_wdata_bits_wstrb_53(fringeCommon_io_dram_0_wdata_bits_wstrb_53),
    .io_dram_0_wdata_bits_wstrb_54(fringeCommon_io_dram_0_wdata_bits_wstrb_54),
    .io_dram_0_wdata_bits_wstrb_55(fringeCommon_io_dram_0_wdata_bits_wstrb_55),
    .io_dram_0_wdata_bits_wstrb_56(fringeCommon_io_dram_0_wdata_bits_wstrb_56),
    .io_dram_0_wdata_bits_wstrb_57(fringeCommon_io_dram_0_wdata_bits_wstrb_57),
    .io_dram_0_wdata_bits_wstrb_58(fringeCommon_io_dram_0_wdata_bits_wstrb_58),
    .io_dram_0_wdata_bits_wstrb_59(fringeCommon_io_dram_0_wdata_bits_wstrb_59),
    .io_dram_0_wdata_bits_wstrb_60(fringeCommon_io_dram_0_wdata_bits_wstrb_60),
    .io_dram_0_wdata_bits_wstrb_61(fringeCommon_io_dram_0_wdata_bits_wstrb_61),
    .io_dram_0_wdata_bits_wstrb_62(fringeCommon_io_dram_0_wdata_bits_wstrb_62),
    .io_dram_0_wdata_bits_wstrb_63(fringeCommon_io_dram_0_wdata_bits_wstrb_63),
    .io_dram_0_wdata_bits_wlast(fringeCommon_io_dram_0_wdata_bits_wlast),
    .io_dram_0_rresp_ready(fringeCommon_io_dram_0_rresp_ready),
    .io_dram_0_wresp_ready(fringeCommon_io_dram_0_wresp_ready),
    .io_dram_0_wresp_valid(fringeCommon_io_dram_0_wresp_valid),
    .io_dram_0_wresp_bits_tag(fringeCommon_io_dram_0_wresp_bits_tag),
    .io_dram_1_cmd_ready(fringeCommon_io_dram_1_cmd_ready),
    .io_dram_1_cmd_valid(fringeCommon_io_dram_1_cmd_valid),
    .io_dram_1_cmd_bits_addr(fringeCommon_io_dram_1_cmd_bits_addr),
    .io_dram_1_cmd_bits_size(fringeCommon_io_dram_1_cmd_bits_size),
    .io_dram_1_cmd_bits_isWr(fringeCommon_io_dram_1_cmd_bits_isWr),
    .io_dram_1_cmd_bits_tag(fringeCommon_io_dram_1_cmd_bits_tag),
    .io_dram_1_wdata_ready(fringeCommon_io_dram_1_wdata_ready),
    .io_dram_1_wdata_valid(fringeCommon_io_dram_1_wdata_valid),
    .io_dram_1_wdata_bits_wdata_0(fringeCommon_io_dram_1_wdata_bits_wdata_0),
    .io_dram_1_wdata_bits_wdata_1(fringeCommon_io_dram_1_wdata_bits_wdata_1),
    .io_dram_1_wdata_bits_wdata_2(fringeCommon_io_dram_1_wdata_bits_wdata_2),
    .io_dram_1_wdata_bits_wdata_3(fringeCommon_io_dram_1_wdata_bits_wdata_3),
    .io_dram_1_wdata_bits_wdata_4(fringeCommon_io_dram_1_wdata_bits_wdata_4),
    .io_dram_1_wdata_bits_wdata_5(fringeCommon_io_dram_1_wdata_bits_wdata_5),
    .io_dram_1_wdata_bits_wdata_6(fringeCommon_io_dram_1_wdata_bits_wdata_6),
    .io_dram_1_wdata_bits_wdata_7(fringeCommon_io_dram_1_wdata_bits_wdata_7),
    .io_dram_1_wdata_bits_wdata_8(fringeCommon_io_dram_1_wdata_bits_wdata_8),
    .io_dram_1_wdata_bits_wdata_9(fringeCommon_io_dram_1_wdata_bits_wdata_9),
    .io_dram_1_wdata_bits_wdata_10(fringeCommon_io_dram_1_wdata_bits_wdata_10),
    .io_dram_1_wdata_bits_wdata_11(fringeCommon_io_dram_1_wdata_bits_wdata_11),
    .io_dram_1_wdata_bits_wdata_12(fringeCommon_io_dram_1_wdata_bits_wdata_12),
    .io_dram_1_wdata_bits_wdata_13(fringeCommon_io_dram_1_wdata_bits_wdata_13),
    .io_dram_1_wdata_bits_wdata_14(fringeCommon_io_dram_1_wdata_bits_wdata_14),
    .io_dram_1_wdata_bits_wdata_15(fringeCommon_io_dram_1_wdata_bits_wdata_15),
    .io_dram_1_wdata_bits_wstrb_0(fringeCommon_io_dram_1_wdata_bits_wstrb_0),
    .io_dram_1_wdata_bits_wstrb_1(fringeCommon_io_dram_1_wdata_bits_wstrb_1),
    .io_dram_1_wdata_bits_wstrb_2(fringeCommon_io_dram_1_wdata_bits_wstrb_2),
    .io_dram_1_wdata_bits_wstrb_3(fringeCommon_io_dram_1_wdata_bits_wstrb_3),
    .io_dram_1_wdata_bits_wstrb_4(fringeCommon_io_dram_1_wdata_bits_wstrb_4),
    .io_dram_1_wdata_bits_wstrb_5(fringeCommon_io_dram_1_wdata_bits_wstrb_5),
    .io_dram_1_wdata_bits_wstrb_6(fringeCommon_io_dram_1_wdata_bits_wstrb_6),
    .io_dram_1_wdata_bits_wstrb_7(fringeCommon_io_dram_1_wdata_bits_wstrb_7),
    .io_dram_1_wdata_bits_wstrb_8(fringeCommon_io_dram_1_wdata_bits_wstrb_8),
    .io_dram_1_wdata_bits_wstrb_9(fringeCommon_io_dram_1_wdata_bits_wstrb_9),
    .io_dram_1_wdata_bits_wstrb_10(fringeCommon_io_dram_1_wdata_bits_wstrb_10),
    .io_dram_1_wdata_bits_wstrb_11(fringeCommon_io_dram_1_wdata_bits_wstrb_11),
    .io_dram_1_wdata_bits_wstrb_12(fringeCommon_io_dram_1_wdata_bits_wstrb_12),
    .io_dram_1_wdata_bits_wstrb_13(fringeCommon_io_dram_1_wdata_bits_wstrb_13),
    .io_dram_1_wdata_bits_wstrb_14(fringeCommon_io_dram_1_wdata_bits_wstrb_14),
    .io_dram_1_wdata_bits_wstrb_15(fringeCommon_io_dram_1_wdata_bits_wstrb_15),
    .io_dram_1_wdata_bits_wstrb_16(fringeCommon_io_dram_1_wdata_bits_wstrb_16),
    .io_dram_1_wdata_bits_wstrb_17(fringeCommon_io_dram_1_wdata_bits_wstrb_17),
    .io_dram_1_wdata_bits_wstrb_18(fringeCommon_io_dram_1_wdata_bits_wstrb_18),
    .io_dram_1_wdata_bits_wstrb_19(fringeCommon_io_dram_1_wdata_bits_wstrb_19),
    .io_dram_1_wdata_bits_wstrb_20(fringeCommon_io_dram_1_wdata_bits_wstrb_20),
    .io_dram_1_wdata_bits_wstrb_21(fringeCommon_io_dram_1_wdata_bits_wstrb_21),
    .io_dram_1_wdata_bits_wstrb_22(fringeCommon_io_dram_1_wdata_bits_wstrb_22),
    .io_dram_1_wdata_bits_wstrb_23(fringeCommon_io_dram_1_wdata_bits_wstrb_23),
    .io_dram_1_wdata_bits_wstrb_24(fringeCommon_io_dram_1_wdata_bits_wstrb_24),
    .io_dram_1_wdata_bits_wstrb_25(fringeCommon_io_dram_1_wdata_bits_wstrb_25),
    .io_dram_1_wdata_bits_wstrb_26(fringeCommon_io_dram_1_wdata_bits_wstrb_26),
    .io_dram_1_wdata_bits_wstrb_27(fringeCommon_io_dram_1_wdata_bits_wstrb_27),
    .io_dram_1_wdata_bits_wstrb_28(fringeCommon_io_dram_1_wdata_bits_wstrb_28),
    .io_dram_1_wdata_bits_wstrb_29(fringeCommon_io_dram_1_wdata_bits_wstrb_29),
    .io_dram_1_wdata_bits_wstrb_30(fringeCommon_io_dram_1_wdata_bits_wstrb_30),
    .io_dram_1_wdata_bits_wstrb_31(fringeCommon_io_dram_1_wdata_bits_wstrb_31),
    .io_dram_1_wdata_bits_wstrb_32(fringeCommon_io_dram_1_wdata_bits_wstrb_32),
    .io_dram_1_wdata_bits_wstrb_33(fringeCommon_io_dram_1_wdata_bits_wstrb_33),
    .io_dram_1_wdata_bits_wstrb_34(fringeCommon_io_dram_1_wdata_bits_wstrb_34),
    .io_dram_1_wdata_bits_wstrb_35(fringeCommon_io_dram_1_wdata_bits_wstrb_35),
    .io_dram_1_wdata_bits_wstrb_36(fringeCommon_io_dram_1_wdata_bits_wstrb_36),
    .io_dram_1_wdata_bits_wstrb_37(fringeCommon_io_dram_1_wdata_bits_wstrb_37),
    .io_dram_1_wdata_bits_wstrb_38(fringeCommon_io_dram_1_wdata_bits_wstrb_38),
    .io_dram_1_wdata_bits_wstrb_39(fringeCommon_io_dram_1_wdata_bits_wstrb_39),
    .io_dram_1_wdata_bits_wstrb_40(fringeCommon_io_dram_1_wdata_bits_wstrb_40),
    .io_dram_1_wdata_bits_wstrb_41(fringeCommon_io_dram_1_wdata_bits_wstrb_41),
    .io_dram_1_wdata_bits_wstrb_42(fringeCommon_io_dram_1_wdata_bits_wstrb_42),
    .io_dram_1_wdata_bits_wstrb_43(fringeCommon_io_dram_1_wdata_bits_wstrb_43),
    .io_dram_1_wdata_bits_wstrb_44(fringeCommon_io_dram_1_wdata_bits_wstrb_44),
    .io_dram_1_wdata_bits_wstrb_45(fringeCommon_io_dram_1_wdata_bits_wstrb_45),
    .io_dram_1_wdata_bits_wstrb_46(fringeCommon_io_dram_1_wdata_bits_wstrb_46),
    .io_dram_1_wdata_bits_wstrb_47(fringeCommon_io_dram_1_wdata_bits_wstrb_47),
    .io_dram_1_wdata_bits_wstrb_48(fringeCommon_io_dram_1_wdata_bits_wstrb_48),
    .io_dram_1_wdata_bits_wstrb_49(fringeCommon_io_dram_1_wdata_bits_wstrb_49),
    .io_dram_1_wdata_bits_wstrb_50(fringeCommon_io_dram_1_wdata_bits_wstrb_50),
    .io_dram_1_wdata_bits_wstrb_51(fringeCommon_io_dram_1_wdata_bits_wstrb_51),
    .io_dram_1_wdata_bits_wstrb_52(fringeCommon_io_dram_1_wdata_bits_wstrb_52),
    .io_dram_1_wdata_bits_wstrb_53(fringeCommon_io_dram_1_wdata_bits_wstrb_53),
    .io_dram_1_wdata_bits_wstrb_54(fringeCommon_io_dram_1_wdata_bits_wstrb_54),
    .io_dram_1_wdata_bits_wstrb_55(fringeCommon_io_dram_1_wdata_bits_wstrb_55),
    .io_dram_1_wdata_bits_wstrb_56(fringeCommon_io_dram_1_wdata_bits_wstrb_56),
    .io_dram_1_wdata_bits_wstrb_57(fringeCommon_io_dram_1_wdata_bits_wstrb_57),
    .io_dram_1_wdata_bits_wstrb_58(fringeCommon_io_dram_1_wdata_bits_wstrb_58),
    .io_dram_1_wdata_bits_wstrb_59(fringeCommon_io_dram_1_wdata_bits_wstrb_59),
    .io_dram_1_wdata_bits_wstrb_60(fringeCommon_io_dram_1_wdata_bits_wstrb_60),
    .io_dram_1_wdata_bits_wstrb_61(fringeCommon_io_dram_1_wdata_bits_wstrb_61),
    .io_dram_1_wdata_bits_wstrb_62(fringeCommon_io_dram_1_wdata_bits_wstrb_62),
    .io_dram_1_wdata_bits_wstrb_63(fringeCommon_io_dram_1_wdata_bits_wstrb_63),
    .io_dram_1_wdata_bits_wlast(fringeCommon_io_dram_1_wdata_bits_wlast),
    .io_dram_1_rresp_ready(fringeCommon_io_dram_1_rresp_ready),
    .io_dram_1_wresp_ready(fringeCommon_io_dram_1_wresp_ready),
    .io_dram_1_wresp_valid(fringeCommon_io_dram_1_wresp_valid),
    .io_dram_1_wresp_bits_tag(fringeCommon_io_dram_1_wresp_bits_tag),
    .io_dram_2_cmd_ready(fringeCommon_io_dram_2_cmd_ready),
    .io_dram_2_cmd_valid(fringeCommon_io_dram_2_cmd_valid),
    .io_dram_2_cmd_bits_addr(fringeCommon_io_dram_2_cmd_bits_addr),
    .io_dram_2_cmd_bits_size(fringeCommon_io_dram_2_cmd_bits_size),
    .io_dram_2_cmd_bits_isWr(fringeCommon_io_dram_2_cmd_bits_isWr),
    .io_dram_2_cmd_bits_tag(fringeCommon_io_dram_2_cmd_bits_tag),
    .io_dram_2_wdata_ready(fringeCommon_io_dram_2_wdata_ready),
    .io_dram_2_wdata_valid(fringeCommon_io_dram_2_wdata_valid),
    .io_dram_2_wdata_bits_wdata_0(fringeCommon_io_dram_2_wdata_bits_wdata_0),
    .io_dram_2_wdata_bits_wdata_1(fringeCommon_io_dram_2_wdata_bits_wdata_1),
    .io_dram_2_wdata_bits_wdata_2(fringeCommon_io_dram_2_wdata_bits_wdata_2),
    .io_dram_2_wdata_bits_wdata_3(fringeCommon_io_dram_2_wdata_bits_wdata_3),
    .io_dram_2_wdata_bits_wdata_4(fringeCommon_io_dram_2_wdata_bits_wdata_4),
    .io_dram_2_wdata_bits_wdata_5(fringeCommon_io_dram_2_wdata_bits_wdata_5),
    .io_dram_2_wdata_bits_wdata_6(fringeCommon_io_dram_2_wdata_bits_wdata_6),
    .io_dram_2_wdata_bits_wdata_7(fringeCommon_io_dram_2_wdata_bits_wdata_7),
    .io_dram_2_wdata_bits_wdata_8(fringeCommon_io_dram_2_wdata_bits_wdata_8),
    .io_dram_2_wdata_bits_wdata_9(fringeCommon_io_dram_2_wdata_bits_wdata_9),
    .io_dram_2_wdata_bits_wdata_10(fringeCommon_io_dram_2_wdata_bits_wdata_10),
    .io_dram_2_wdata_bits_wdata_11(fringeCommon_io_dram_2_wdata_bits_wdata_11),
    .io_dram_2_wdata_bits_wdata_12(fringeCommon_io_dram_2_wdata_bits_wdata_12),
    .io_dram_2_wdata_bits_wdata_13(fringeCommon_io_dram_2_wdata_bits_wdata_13),
    .io_dram_2_wdata_bits_wdata_14(fringeCommon_io_dram_2_wdata_bits_wdata_14),
    .io_dram_2_wdata_bits_wdata_15(fringeCommon_io_dram_2_wdata_bits_wdata_15),
    .io_dram_2_wdata_bits_wstrb_0(fringeCommon_io_dram_2_wdata_bits_wstrb_0),
    .io_dram_2_wdata_bits_wstrb_1(fringeCommon_io_dram_2_wdata_bits_wstrb_1),
    .io_dram_2_wdata_bits_wstrb_2(fringeCommon_io_dram_2_wdata_bits_wstrb_2),
    .io_dram_2_wdata_bits_wstrb_3(fringeCommon_io_dram_2_wdata_bits_wstrb_3),
    .io_dram_2_wdata_bits_wstrb_4(fringeCommon_io_dram_2_wdata_bits_wstrb_4),
    .io_dram_2_wdata_bits_wstrb_5(fringeCommon_io_dram_2_wdata_bits_wstrb_5),
    .io_dram_2_wdata_bits_wstrb_6(fringeCommon_io_dram_2_wdata_bits_wstrb_6),
    .io_dram_2_wdata_bits_wstrb_7(fringeCommon_io_dram_2_wdata_bits_wstrb_7),
    .io_dram_2_wdata_bits_wstrb_8(fringeCommon_io_dram_2_wdata_bits_wstrb_8),
    .io_dram_2_wdata_bits_wstrb_9(fringeCommon_io_dram_2_wdata_bits_wstrb_9),
    .io_dram_2_wdata_bits_wstrb_10(fringeCommon_io_dram_2_wdata_bits_wstrb_10),
    .io_dram_2_wdata_bits_wstrb_11(fringeCommon_io_dram_2_wdata_bits_wstrb_11),
    .io_dram_2_wdata_bits_wstrb_12(fringeCommon_io_dram_2_wdata_bits_wstrb_12),
    .io_dram_2_wdata_bits_wstrb_13(fringeCommon_io_dram_2_wdata_bits_wstrb_13),
    .io_dram_2_wdata_bits_wstrb_14(fringeCommon_io_dram_2_wdata_bits_wstrb_14),
    .io_dram_2_wdata_bits_wstrb_15(fringeCommon_io_dram_2_wdata_bits_wstrb_15),
    .io_dram_2_wdata_bits_wstrb_16(fringeCommon_io_dram_2_wdata_bits_wstrb_16),
    .io_dram_2_wdata_bits_wstrb_17(fringeCommon_io_dram_2_wdata_bits_wstrb_17),
    .io_dram_2_wdata_bits_wstrb_18(fringeCommon_io_dram_2_wdata_bits_wstrb_18),
    .io_dram_2_wdata_bits_wstrb_19(fringeCommon_io_dram_2_wdata_bits_wstrb_19),
    .io_dram_2_wdata_bits_wstrb_20(fringeCommon_io_dram_2_wdata_bits_wstrb_20),
    .io_dram_2_wdata_bits_wstrb_21(fringeCommon_io_dram_2_wdata_bits_wstrb_21),
    .io_dram_2_wdata_bits_wstrb_22(fringeCommon_io_dram_2_wdata_bits_wstrb_22),
    .io_dram_2_wdata_bits_wstrb_23(fringeCommon_io_dram_2_wdata_bits_wstrb_23),
    .io_dram_2_wdata_bits_wstrb_24(fringeCommon_io_dram_2_wdata_bits_wstrb_24),
    .io_dram_2_wdata_bits_wstrb_25(fringeCommon_io_dram_2_wdata_bits_wstrb_25),
    .io_dram_2_wdata_bits_wstrb_26(fringeCommon_io_dram_2_wdata_bits_wstrb_26),
    .io_dram_2_wdata_bits_wstrb_27(fringeCommon_io_dram_2_wdata_bits_wstrb_27),
    .io_dram_2_wdata_bits_wstrb_28(fringeCommon_io_dram_2_wdata_bits_wstrb_28),
    .io_dram_2_wdata_bits_wstrb_29(fringeCommon_io_dram_2_wdata_bits_wstrb_29),
    .io_dram_2_wdata_bits_wstrb_30(fringeCommon_io_dram_2_wdata_bits_wstrb_30),
    .io_dram_2_wdata_bits_wstrb_31(fringeCommon_io_dram_2_wdata_bits_wstrb_31),
    .io_dram_2_wdata_bits_wstrb_32(fringeCommon_io_dram_2_wdata_bits_wstrb_32),
    .io_dram_2_wdata_bits_wstrb_33(fringeCommon_io_dram_2_wdata_bits_wstrb_33),
    .io_dram_2_wdata_bits_wstrb_34(fringeCommon_io_dram_2_wdata_bits_wstrb_34),
    .io_dram_2_wdata_bits_wstrb_35(fringeCommon_io_dram_2_wdata_bits_wstrb_35),
    .io_dram_2_wdata_bits_wstrb_36(fringeCommon_io_dram_2_wdata_bits_wstrb_36),
    .io_dram_2_wdata_bits_wstrb_37(fringeCommon_io_dram_2_wdata_bits_wstrb_37),
    .io_dram_2_wdata_bits_wstrb_38(fringeCommon_io_dram_2_wdata_bits_wstrb_38),
    .io_dram_2_wdata_bits_wstrb_39(fringeCommon_io_dram_2_wdata_bits_wstrb_39),
    .io_dram_2_wdata_bits_wstrb_40(fringeCommon_io_dram_2_wdata_bits_wstrb_40),
    .io_dram_2_wdata_bits_wstrb_41(fringeCommon_io_dram_2_wdata_bits_wstrb_41),
    .io_dram_2_wdata_bits_wstrb_42(fringeCommon_io_dram_2_wdata_bits_wstrb_42),
    .io_dram_2_wdata_bits_wstrb_43(fringeCommon_io_dram_2_wdata_bits_wstrb_43),
    .io_dram_2_wdata_bits_wstrb_44(fringeCommon_io_dram_2_wdata_bits_wstrb_44),
    .io_dram_2_wdata_bits_wstrb_45(fringeCommon_io_dram_2_wdata_bits_wstrb_45),
    .io_dram_2_wdata_bits_wstrb_46(fringeCommon_io_dram_2_wdata_bits_wstrb_46),
    .io_dram_2_wdata_bits_wstrb_47(fringeCommon_io_dram_2_wdata_bits_wstrb_47),
    .io_dram_2_wdata_bits_wstrb_48(fringeCommon_io_dram_2_wdata_bits_wstrb_48),
    .io_dram_2_wdata_bits_wstrb_49(fringeCommon_io_dram_2_wdata_bits_wstrb_49),
    .io_dram_2_wdata_bits_wstrb_50(fringeCommon_io_dram_2_wdata_bits_wstrb_50),
    .io_dram_2_wdata_bits_wstrb_51(fringeCommon_io_dram_2_wdata_bits_wstrb_51),
    .io_dram_2_wdata_bits_wstrb_52(fringeCommon_io_dram_2_wdata_bits_wstrb_52),
    .io_dram_2_wdata_bits_wstrb_53(fringeCommon_io_dram_2_wdata_bits_wstrb_53),
    .io_dram_2_wdata_bits_wstrb_54(fringeCommon_io_dram_2_wdata_bits_wstrb_54),
    .io_dram_2_wdata_bits_wstrb_55(fringeCommon_io_dram_2_wdata_bits_wstrb_55),
    .io_dram_2_wdata_bits_wstrb_56(fringeCommon_io_dram_2_wdata_bits_wstrb_56),
    .io_dram_2_wdata_bits_wstrb_57(fringeCommon_io_dram_2_wdata_bits_wstrb_57),
    .io_dram_2_wdata_bits_wstrb_58(fringeCommon_io_dram_2_wdata_bits_wstrb_58),
    .io_dram_2_wdata_bits_wstrb_59(fringeCommon_io_dram_2_wdata_bits_wstrb_59),
    .io_dram_2_wdata_bits_wstrb_60(fringeCommon_io_dram_2_wdata_bits_wstrb_60),
    .io_dram_2_wdata_bits_wstrb_61(fringeCommon_io_dram_2_wdata_bits_wstrb_61),
    .io_dram_2_wdata_bits_wstrb_62(fringeCommon_io_dram_2_wdata_bits_wstrb_62),
    .io_dram_2_wdata_bits_wstrb_63(fringeCommon_io_dram_2_wdata_bits_wstrb_63),
    .io_dram_2_wdata_bits_wlast(fringeCommon_io_dram_2_wdata_bits_wlast),
    .io_dram_2_rresp_ready(fringeCommon_io_dram_2_rresp_ready),
    .io_dram_2_wresp_ready(fringeCommon_io_dram_2_wresp_ready),
    .io_dram_2_wresp_valid(fringeCommon_io_dram_2_wresp_valid),
    .io_dram_2_wresp_bits_tag(fringeCommon_io_dram_2_wresp_bits_tag),
    .io_dram_3_cmd_ready(fringeCommon_io_dram_3_cmd_ready),
    .io_dram_3_cmd_valid(fringeCommon_io_dram_3_cmd_valid),
    .io_dram_3_cmd_bits_addr(fringeCommon_io_dram_3_cmd_bits_addr),
    .io_dram_3_cmd_bits_size(fringeCommon_io_dram_3_cmd_bits_size),
    .io_dram_3_cmd_bits_isWr(fringeCommon_io_dram_3_cmd_bits_isWr),
    .io_dram_3_cmd_bits_tag(fringeCommon_io_dram_3_cmd_bits_tag),
    .io_dram_3_wdata_ready(fringeCommon_io_dram_3_wdata_ready),
    .io_dram_3_wdata_valid(fringeCommon_io_dram_3_wdata_valid),
    .io_dram_3_wdata_bits_wdata_0(fringeCommon_io_dram_3_wdata_bits_wdata_0),
    .io_dram_3_wdata_bits_wdata_1(fringeCommon_io_dram_3_wdata_bits_wdata_1),
    .io_dram_3_wdata_bits_wdata_2(fringeCommon_io_dram_3_wdata_bits_wdata_2),
    .io_dram_3_wdata_bits_wdata_3(fringeCommon_io_dram_3_wdata_bits_wdata_3),
    .io_dram_3_wdata_bits_wdata_4(fringeCommon_io_dram_3_wdata_bits_wdata_4),
    .io_dram_3_wdata_bits_wdata_5(fringeCommon_io_dram_3_wdata_bits_wdata_5),
    .io_dram_3_wdata_bits_wdata_6(fringeCommon_io_dram_3_wdata_bits_wdata_6),
    .io_dram_3_wdata_bits_wdata_7(fringeCommon_io_dram_3_wdata_bits_wdata_7),
    .io_dram_3_wdata_bits_wdata_8(fringeCommon_io_dram_3_wdata_bits_wdata_8),
    .io_dram_3_wdata_bits_wdata_9(fringeCommon_io_dram_3_wdata_bits_wdata_9),
    .io_dram_3_wdata_bits_wdata_10(fringeCommon_io_dram_3_wdata_bits_wdata_10),
    .io_dram_3_wdata_bits_wdata_11(fringeCommon_io_dram_3_wdata_bits_wdata_11),
    .io_dram_3_wdata_bits_wdata_12(fringeCommon_io_dram_3_wdata_bits_wdata_12),
    .io_dram_3_wdata_bits_wdata_13(fringeCommon_io_dram_3_wdata_bits_wdata_13),
    .io_dram_3_wdata_bits_wdata_14(fringeCommon_io_dram_3_wdata_bits_wdata_14),
    .io_dram_3_wdata_bits_wdata_15(fringeCommon_io_dram_3_wdata_bits_wdata_15),
    .io_dram_3_wdata_bits_wstrb_0(fringeCommon_io_dram_3_wdata_bits_wstrb_0),
    .io_dram_3_wdata_bits_wstrb_1(fringeCommon_io_dram_3_wdata_bits_wstrb_1),
    .io_dram_3_wdata_bits_wstrb_2(fringeCommon_io_dram_3_wdata_bits_wstrb_2),
    .io_dram_3_wdata_bits_wstrb_3(fringeCommon_io_dram_3_wdata_bits_wstrb_3),
    .io_dram_3_wdata_bits_wstrb_4(fringeCommon_io_dram_3_wdata_bits_wstrb_4),
    .io_dram_3_wdata_bits_wstrb_5(fringeCommon_io_dram_3_wdata_bits_wstrb_5),
    .io_dram_3_wdata_bits_wstrb_6(fringeCommon_io_dram_3_wdata_bits_wstrb_6),
    .io_dram_3_wdata_bits_wstrb_7(fringeCommon_io_dram_3_wdata_bits_wstrb_7),
    .io_dram_3_wdata_bits_wstrb_8(fringeCommon_io_dram_3_wdata_bits_wstrb_8),
    .io_dram_3_wdata_bits_wstrb_9(fringeCommon_io_dram_3_wdata_bits_wstrb_9),
    .io_dram_3_wdata_bits_wstrb_10(fringeCommon_io_dram_3_wdata_bits_wstrb_10),
    .io_dram_3_wdata_bits_wstrb_11(fringeCommon_io_dram_3_wdata_bits_wstrb_11),
    .io_dram_3_wdata_bits_wstrb_12(fringeCommon_io_dram_3_wdata_bits_wstrb_12),
    .io_dram_3_wdata_bits_wstrb_13(fringeCommon_io_dram_3_wdata_bits_wstrb_13),
    .io_dram_3_wdata_bits_wstrb_14(fringeCommon_io_dram_3_wdata_bits_wstrb_14),
    .io_dram_3_wdata_bits_wstrb_15(fringeCommon_io_dram_3_wdata_bits_wstrb_15),
    .io_dram_3_wdata_bits_wstrb_16(fringeCommon_io_dram_3_wdata_bits_wstrb_16),
    .io_dram_3_wdata_bits_wstrb_17(fringeCommon_io_dram_3_wdata_bits_wstrb_17),
    .io_dram_3_wdata_bits_wstrb_18(fringeCommon_io_dram_3_wdata_bits_wstrb_18),
    .io_dram_3_wdata_bits_wstrb_19(fringeCommon_io_dram_3_wdata_bits_wstrb_19),
    .io_dram_3_wdata_bits_wstrb_20(fringeCommon_io_dram_3_wdata_bits_wstrb_20),
    .io_dram_3_wdata_bits_wstrb_21(fringeCommon_io_dram_3_wdata_bits_wstrb_21),
    .io_dram_3_wdata_bits_wstrb_22(fringeCommon_io_dram_3_wdata_bits_wstrb_22),
    .io_dram_3_wdata_bits_wstrb_23(fringeCommon_io_dram_3_wdata_bits_wstrb_23),
    .io_dram_3_wdata_bits_wstrb_24(fringeCommon_io_dram_3_wdata_bits_wstrb_24),
    .io_dram_3_wdata_bits_wstrb_25(fringeCommon_io_dram_3_wdata_bits_wstrb_25),
    .io_dram_3_wdata_bits_wstrb_26(fringeCommon_io_dram_3_wdata_bits_wstrb_26),
    .io_dram_3_wdata_bits_wstrb_27(fringeCommon_io_dram_3_wdata_bits_wstrb_27),
    .io_dram_3_wdata_bits_wstrb_28(fringeCommon_io_dram_3_wdata_bits_wstrb_28),
    .io_dram_3_wdata_bits_wstrb_29(fringeCommon_io_dram_3_wdata_bits_wstrb_29),
    .io_dram_3_wdata_bits_wstrb_30(fringeCommon_io_dram_3_wdata_bits_wstrb_30),
    .io_dram_3_wdata_bits_wstrb_31(fringeCommon_io_dram_3_wdata_bits_wstrb_31),
    .io_dram_3_wdata_bits_wstrb_32(fringeCommon_io_dram_3_wdata_bits_wstrb_32),
    .io_dram_3_wdata_bits_wstrb_33(fringeCommon_io_dram_3_wdata_bits_wstrb_33),
    .io_dram_3_wdata_bits_wstrb_34(fringeCommon_io_dram_3_wdata_bits_wstrb_34),
    .io_dram_3_wdata_bits_wstrb_35(fringeCommon_io_dram_3_wdata_bits_wstrb_35),
    .io_dram_3_wdata_bits_wstrb_36(fringeCommon_io_dram_3_wdata_bits_wstrb_36),
    .io_dram_3_wdata_bits_wstrb_37(fringeCommon_io_dram_3_wdata_bits_wstrb_37),
    .io_dram_3_wdata_bits_wstrb_38(fringeCommon_io_dram_3_wdata_bits_wstrb_38),
    .io_dram_3_wdata_bits_wstrb_39(fringeCommon_io_dram_3_wdata_bits_wstrb_39),
    .io_dram_3_wdata_bits_wstrb_40(fringeCommon_io_dram_3_wdata_bits_wstrb_40),
    .io_dram_3_wdata_bits_wstrb_41(fringeCommon_io_dram_3_wdata_bits_wstrb_41),
    .io_dram_3_wdata_bits_wstrb_42(fringeCommon_io_dram_3_wdata_bits_wstrb_42),
    .io_dram_3_wdata_bits_wstrb_43(fringeCommon_io_dram_3_wdata_bits_wstrb_43),
    .io_dram_3_wdata_bits_wstrb_44(fringeCommon_io_dram_3_wdata_bits_wstrb_44),
    .io_dram_3_wdata_bits_wstrb_45(fringeCommon_io_dram_3_wdata_bits_wstrb_45),
    .io_dram_3_wdata_bits_wstrb_46(fringeCommon_io_dram_3_wdata_bits_wstrb_46),
    .io_dram_3_wdata_bits_wstrb_47(fringeCommon_io_dram_3_wdata_bits_wstrb_47),
    .io_dram_3_wdata_bits_wstrb_48(fringeCommon_io_dram_3_wdata_bits_wstrb_48),
    .io_dram_3_wdata_bits_wstrb_49(fringeCommon_io_dram_3_wdata_bits_wstrb_49),
    .io_dram_3_wdata_bits_wstrb_50(fringeCommon_io_dram_3_wdata_bits_wstrb_50),
    .io_dram_3_wdata_bits_wstrb_51(fringeCommon_io_dram_3_wdata_bits_wstrb_51),
    .io_dram_3_wdata_bits_wstrb_52(fringeCommon_io_dram_3_wdata_bits_wstrb_52),
    .io_dram_3_wdata_bits_wstrb_53(fringeCommon_io_dram_3_wdata_bits_wstrb_53),
    .io_dram_3_wdata_bits_wstrb_54(fringeCommon_io_dram_3_wdata_bits_wstrb_54),
    .io_dram_3_wdata_bits_wstrb_55(fringeCommon_io_dram_3_wdata_bits_wstrb_55),
    .io_dram_3_wdata_bits_wstrb_56(fringeCommon_io_dram_3_wdata_bits_wstrb_56),
    .io_dram_3_wdata_bits_wstrb_57(fringeCommon_io_dram_3_wdata_bits_wstrb_57),
    .io_dram_3_wdata_bits_wstrb_58(fringeCommon_io_dram_3_wdata_bits_wstrb_58),
    .io_dram_3_wdata_bits_wstrb_59(fringeCommon_io_dram_3_wdata_bits_wstrb_59),
    .io_dram_3_wdata_bits_wstrb_60(fringeCommon_io_dram_3_wdata_bits_wstrb_60),
    .io_dram_3_wdata_bits_wstrb_61(fringeCommon_io_dram_3_wdata_bits_wstrb_61),
    .io_dram_3_wdata_bits_wstrb_62(fringeCommon_io_dram_3_wdata_bits_wstrb_62),
    .io_dram_3_wdata_bits_wstrb_63(fringeCommon_io_dram_3_wdata_bits_wstrb_63),
    .io_dram_3_wdata_bits_wlast(fringeCommon_io_dram_3_wdata_bits_wlast),
    .io_dram_3_rresp_ready(fringeCommon_io_dram_3_rresp_ready),
    .io_dram_3_wresp_ready(fringeCommon_io_dram_3_wresp_ready),
    .io_dram_3_wresp_valid(fringeCommon_io_dram_3_wresp_valid),
    .io_dram_3_wresp_bits_tag(fringeCommon_io_dram_3_wresp_bits_tag),
    .io_heap_0_req_valid(fringeCommon_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(fringeCommon_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(fringeCommon_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(fringeCommon_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(fringeCommon_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(fringeCommon_io_heap_0_resp_bits_sizeAddr)
  );
  AXI4LiteToRFBridge AXI4LiteToRFBridge ( // @[FringeZynq.scala 90:31:@145532.4]
    .clock(AXI4LiteToRFBridge_clock),
    .reset(AXI4LiteToRFBridge_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridge_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridge_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridge_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridge_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridge_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridge_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridge_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridge_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridge_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridge_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridge_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridge_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridge_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridge_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridge_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridge_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridge_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridge_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridge_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridge_io_raddr),
    .io_wen(AXI4LiteToRFBridge_io_wen),
    .io_waddr(AXI4LiteToRFBridge_io_waddr),
    .io_wdata(AXI4LiteToRFBridge_io_wdata),
    .io_rdata(AXI4LiteToRFBridge_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 131:27:@145682.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_1 ( // @[FringeZynq.scala 131:27:@145838.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_1_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_1_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_1_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_1_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_1_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_1_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_1_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_1_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_1_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_1_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_1_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_1_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_1_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_1_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_1_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_1_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_1_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_1_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_1_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_1_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_1_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_1_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_1_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_1_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_1_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_1_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_1_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_1_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_1_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_1_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_1_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_1_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_2 ( // @[FringeZynq.scala 131:27:@145994.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_2_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_2_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_2_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_2_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_2_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_2_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_2_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_2_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_2_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_2_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_2_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_2_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_2_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_2_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_2_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_2_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_2_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_2_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_2_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_2_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_2_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_2_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_2_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_2_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_2_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_2_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_2_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_2_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_2_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_2_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_2_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_2_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_3 ( // @[FringeZynq.scala 131:27:@146150.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_3_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_3_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_3_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_3_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_3_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_3_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_3_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_3_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_3_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_3_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_3_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_3_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_3_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_3_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_3_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_3_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_3_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_3_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_3_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_3_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_3_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_3_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_3_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_3_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_3_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_3_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_3_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_3_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_3_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_3_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_3_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_3_io_M_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 91:28:@145550.4]
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 91:28:@145546.4]
  assign io_S_AXI_WREADY = AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 91:28:@145542.4]
  assign io_S_AXI_RDATA = AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 91:28:@145541.4]
  assign io_S_AXI_RRESP = AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 91:28:@145540.4]
  assign io_S_AXI_RVALID = AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 91:28:@145539.4]
  assign io_S_AXI_BRESP = AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 91:28:@145537.4]
  assign io_S_AXI_BVALID = AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 91:28:@145536.4]
  assign io_M_AXI_0_AWID = MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@145837.4]
  assign io_M_AXI_0_AWADDR = MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@145835.4]
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@145834.4]
  assign io_M_AXI_0_AWVALID = MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@145827.4]
  assign io_M_AXI_0_ARID = MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@145825.4]
  assign io_M_AXI_0_ARADDR = MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@145823.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@145822.4]
  assign io_M_AXI_0_ARVALID = MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@145815.4]
  assign io_M_AXI_0_WDATA = MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@145813.4]
  assign io_M_AXI_0_WSTRB = MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@145812.4]
  assign io_M_AXI_0_WLAST = MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@145811.4]
  assign io_M_AXI_0_WVALID = MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@145810.4]
  assign io_M_AXI_0_RREADY = MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@145802.4]
  assign io_M_AXI_0_BREADY = MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@145797.4]
  assign io_M_AXI_1_AWID = MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@145993.4]
  assign io_M_AXI_1_AWADDR = MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@145991.4]
  assign io_M_AXI_1_AWLEN = MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@145990.4]
  assign io_M_AXI_1_AWVALID = MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@145983.4]
  assign io_M_AXI_1_ARID = MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@145981.4]
  assign io_M_AXI_1_ARADDR = MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@145979.4]
  assign io_M_AXI_1_ARLEN = MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@145978.4]
  assign io_M_AXI_1_ARVALID = MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@145971.4]
  assign io_M_AXI_1_WDATA = MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@145969.4]
  assign io_M_AXI_1_WSTRB = MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@145968.4]
  assign io_M_AXI_1_WLAST = MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@145967.4]
  assign io_M_AXI_1_WVALID = MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@145966.4]
  assign io_M_AXI_1_RREADY = MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@145958.4]
  assign io_M_AXI_1_BREADY = MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@145953.4]
  assign io_M_AXI_2_AWID = MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@146149.4]
  assign io_M_AXI_2_AWADDR = MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@146147.4]
  assign io_M_AXI_2_AWLEN = MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@146146.4]
  assign io_M_AXI_2_AWVALID = MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@146139.4]
  assign io_M_AXI_2_ARID = MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@146137.4]
  assign io_M_AXI_2_ARADDR = MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@146135.4]
  assign io_M_AXI_2_ARLEN = MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@146134.4]
  assign io_M_AXI_2_ARVALID = MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@146127.4]
  assign io_M_AXI_2_WDATA = MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@146125.4]
  assign io_M_AXI_2_WSTRB = MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@146124.4]
  assign io_M_AXI_2_WLAST = MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@146123.4]
  assign io_M_AXI_2_WVALID = MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@146122.4]
  assign io_M_AXI_2_RREADY = MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@146114.4]
  assign io_M_AXI_2_BREADY = MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@146109.4]
  assign io_M_AXI_3_AWID = MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@146305.4]
  assign io_M_AXI_3_AWADDR = MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@146303.4]
  assign io_M_AXI_3_AWLEN = MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@146302.4]
  assign io_M_AXI_3_AWVALID = MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@146295.4]
  assign io_M_AXI_3_ARID = MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@146293.4]
  assign io_M_AXI_3_ARADDR = MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@146291.4]
  assign io_M_AXI_3_ARLEN = MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@146290.4]
  assign io_M_AXI_3_ARVALID = MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@146283.4]
  assign io_M_AXI_3_WDATA = MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@146281.4]
  assign io_M_AXI_3_WSTRB = MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@146280.4]
  assign io_M_AXI_3_WLAST = MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@146279.4]
  assign io_M_AXI_3_WVALID = MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@146278.4]
  assign io_M_AXI_3_RREADY = MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@146270.4]
  assign io_M_AXI_3_BREADY = MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@146265.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 115:13:@145560.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 119:12:@145564.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 121:13:@145565.4]
  assign io_argIns_1 = fringeCommon_io_argIns_1; // @[FringeZynq.scala 121:13:@145566.4]
  assign io_memStreams_stores_0_cmd_ready = fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 126:17:@145653.4]
  assign io_memStreams_stores_0_data_ready = fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 126:17:@145649.4]
  assign io_memStreams_stores_0_wresp_valid = fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 126:17:@145644.4]
  assign io_memStreams_stores_0_wresp_bits = fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 126:17:@145643.4]
  assign io_heap_0_resp_valid = fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 127:11:@145678.4]
  assign io_heap_0_resp_bits_allocDealloc = fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 127:11:@145677.4]
  assign io_heap_0_resp_bits_sizeAddr = fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 127:11:@145676.4]
  assign fringeCommon_clock = clock; // @[:@144627.4]
  assign fringeCommon_reset = reset; // @[:@144628.4 FringeZynq.scala 117:22:@145563.4]
  assign fringeCommon_io_raddr = AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 94:27:@145554.4]
  assign fringeCommon_io_wen = AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 95:27:@145555.4]
  assign fringeCommon_io_waddr = AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 96:27:@145556.4]
  assign fringeCommon_io_wdata = {{32'd0}, AXI4LiteToRFBridge_io_wdata}; // @[FringeZynq.scala 97:27:@145557.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 116:24:@145561.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 122:27:@145568.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 122:27:@145567.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 126:17:@145652.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 126:17:@145651.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 126:17:@145650.4]
  assign fringeCommon_io_memStreams_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 126:17:@145648.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 126:17:@145647.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 126:17:@145646.4]
  assign fringeCommon_io_memStreams_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 126:17:@145645.4]
  assign fringeCommon_io_dram_0_cmd_ready = MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@145796.4]
  assign fringeCommon_io_dram_0_wdata_ready = MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@145789.4]
  assign fringeCommon_io_dram_0_wresp_valid = MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@145686.4]
  assign fringeCommon_io_dram_0_wresp_bits_tag = MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@145685.4]
  assign fringeCommon_io_dram_1_cmd_ready = MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@145952.4]
  assign fringeCommon_io_dram_1_wdata_ready = MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@145945.4]
  assign fringeCommon_io_dram_1_wresp_valid = MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@145842.4]
  assign fringeCommon_io_dram_1_wresp_bits_tag = MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@145841.4]
  assign fringeCommon_io_dram_2_cmd_ready = MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@146108.4]
  assign fringeCommon_io_dram_2_wdata_ready = MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@146101.4]
  assign fringeCommon_io_dram_2_wresp_valid = MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@145998.4]
  assign fringeCommon_io_dram_2_wresp_bits_tag = MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@145997.4]
  assign fringeCommon_io_dram_3_cmd_ready = MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@146264.4]
  assign fringeCommon_io_dram_3_wdata_ready = MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@146257.4]
  assign fringeCommon_io_dram_3_wresp_valid = MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@146154.4]
  assign fringeCommon_io_dram_3_wresp_bits_tag = MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@146153.4]
  assign fringeCommon_io_heap_0_req_valid = io_heap_0_req_valid; // @[FringeZynq.scala 127:11:@145681.4]
  assign fringeCommon_io_heap_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 127:11:@145680.4]
  assign fringeCommon_io_heap_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 127:11:@145679.4]
  assign AXI4LiteToRFBridge_clock = clock; // @[:@145533.4]
  assign AXI4LiteToRFBridge_reset = reset; // @[:@145534.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[FringeZynq.scala 91:28:@145553.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[FringeZynq.scala 91:28:@145552.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[FringeZynq.scala 91:28:@145551.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[FringeZynq.scala 91:28:@145549.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[FringeZynq.scala 91:28:@145548.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[FringeZynq.scala 91:28:@145547.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[FringeZynq.scala 91:28:@145545.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[FringeZynq.scala 91:28:@145544.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[FringeZynq.scala 91:28:@145543.4]
  assign AXI4LiteToRFBridge_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[FringeZynq.scala 91:28:@145538.4]
  assign AXI4LiteToRFBridge_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[FringeZynq.scala 91:28:@145535.4]
  assign AXI4LiteToRFBridge_io_rdata = fringeCommon_io_rdata[31:0]; // @[FringeZynq.scala 98:28:@145558.4]
  assign MAGToAXI4Bridge_io_in_cmd_valid = fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 132:21:@145795.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_addr = fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 132:21:@145794.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_size = fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 132:21:@145793.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_isWr = fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@145791.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_tag = fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 132:21:@145790.4]
  assign MAGToAXI4Bridge_io_in_wdata_valid = fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 132:21:@145788.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@145772.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@145773.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@145774.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@145775.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@145776.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@145777.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@145778.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@145779.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@145780.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@145781.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@145782.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@145783.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@145784.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@145785.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@145786.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@145787.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@145708.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@145709.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@145710.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@145711.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@145712.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@145713.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@145714.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@145715.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@145716.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@145717.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@145718.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@145719.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@145720.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@145721.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@145722.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@145723.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@145724.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@145725.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@145726.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@145727.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@145728.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@145729.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@145730.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@145731.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@145732.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@145733.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@145734.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@145735.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@145736.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@145737.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@145738.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@145739.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@145740.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@145741.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@145742.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@145743.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@145744.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@145745.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@145746.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@145747.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@145748.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@145749.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@145750.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@145751.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@145752.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@145753.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@145754.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@145755.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@145756.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@145757.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@145758.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@145759.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@145760.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@145761.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@145762.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@145763.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@145764.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@145765.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@145766.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@145767.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@145768.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@145769.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@145770.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@145771.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wlast = fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@145707.4]
  assign MAGToAXI4Bridge_io_in_rresp_ready = fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 132:21:@145706.4]
  assign MAGToAXI4Bridge_io_in_wresp_ready = fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 132:21:@145687.4]
  assign MAGToAXI4Bridge_io_M_AXI_AWREADY = io_M_AXI_0_AWREADY; // @[FringeZynq.scala 133:10:@145826.4]
  assign MAGToAXI4Bridge_io_M_AXI_ARREADY = io_M_AXI_0_ARREADY; // @[FringeZynq.scala 133:10:@145814.4]
  assign MAGToAXI4Bridge_io_M_AXI_WREADY = io_M_AXI_0_WREADY; // @[FringeZynq.scala 133:10:@145809.4]
  assign MAGToAXI4Bridge_io_M_AXI_BID = io_M_AXI_0_BID; // @[FringeZynq.scala 133:10:@145801.4]
  assign MAGToAXI4Bridge_io_M_AXI_BVALID = io_M_AXI_0_BVALID; // @[FringeZynq.scala 133:10:@145798.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_valid = fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 132:21:@145951.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_addr = fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 132:21:@145950.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_size = fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 132:21:@145949.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_isWr = fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@145947.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_tag = fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 132:21:@145946.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_valid = fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 132:21:@145944.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@145928.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@145929.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@145930.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@145931.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@145932.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@145933.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@145934.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@145935.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@145936.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@145937.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@145938.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@145939.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@145940.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@145941.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@145942.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@145943.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@145864.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@145865.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@145866.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@145867.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@145868.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@145869.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@145870.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@145871.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@145872.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@145873.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@145874.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@145875.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@145876.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@145877.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@145878.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@145879.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@145880.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@145881.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@145882.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@145883.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@145884.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@145885.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@145886.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@145887.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@145888.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@145889.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@145890.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@145891.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@145892.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@145893.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@145894.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@145895.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@145896.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@145897.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@145898.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@145899.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@145900.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@145901.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@145902.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@145903.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@145904.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@145905.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@145906.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@145907.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@145908.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@145909.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@145910.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@145911.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@145912.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@145913.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@145914.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@145915.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@145916.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@145917.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@145918.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@145919.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@145920.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@145921.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@145922.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@145923.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@145924.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@145925.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@145926.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@145927.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wlast = fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@145863.4]
  assign MAGToAXI4Bridge_1_io_in_rresp_ready = fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 132:21:@145862.4]
  assign MAGToAXI4Bridge_1_io_in_wresp_ready = fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 132:21:@145843.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_AWREADY = io_M_AXI_1_AWREADY; // @[FringeZynq.scala 133:10:@145982.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_ARREADY = io_M_AXI_1_ARREADY; // @[FringeZynq.scala 133:10:@145970.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_WREADY = io_M_AXI_1_WREADY; // @[FringeZynq.scala 133:10:@145965.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BID = io_M_AXI_1_BID; // @[FringeZynq.scala 133:10:@145957.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BVALID = io_M_AXI_1_BVALID; // @[FringeZynq.scala 133:10:@145954.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_valid = fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 132:21:@146107.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_addr = fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 132:21:@146106.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_size = fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 132:21:@146105.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_isWr = fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@146103.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_tag = fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 132:21:@146102.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_valid = fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 132:21:@146100.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@146084.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@146085.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@146086.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@146087.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@146088.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@146089.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@146090.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@146091.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@146092.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@146093.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@146094.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@146095.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@146096.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@146097.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@146098.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@146099.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@146020.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@146021.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@146022.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@146023.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@146024.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@146025.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@146026.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@146027.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@146028.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@146029.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@146030.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@146031.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@146032.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@146033.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@146034.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@146035.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@146036.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@146037.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@146038.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@146039.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@146040.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@146041.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@146042.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@146043.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@146044.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@146045.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@146046.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@146047.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@146048.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@146049.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@146050.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@146051.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@146052.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@146053.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@146054.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@146055.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@146056.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@146057.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@146058.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@146059.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@146060.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@146061.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@146062.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@146063.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@146064.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@146065.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@146066.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@146067.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@146068.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@146069.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@146070.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@146071.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@146072.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@146073.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@146074.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@146075.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@146076.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@146077.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@146078.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@146079.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@146080.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@146081.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@146082.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@146083.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wlast = fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@146019.4]
  assign MAGToAXI4Bridge_2_io_in_rresp_ready = fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 132:21:@146018.4]
  assign MAGToAXI4Bridge_2_io_in_wresp_ready = fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 132:21:@145999.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_AWREADY = io_M_AXI_2_AWREADY; // @[FringeZynq.scala 133:10:@146138.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_ARREADY = io_M_AXI_2_ARREADY; // @[FringeZynq.scala 133:10:@146126.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_WREADY = io_M_AXI_2_WREADY; // @[FringeZynq.scala 133:10:@146121.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BID = io_M_AXI_2_BID; // @[FringeZynq.scala 133:10:@146113.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BVALID = io_M_AXI_2_BVALID; // @[FringeZynq.scala 133:10:@146110.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_valid = fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 132:21:@146263.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_addr = fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 132:21:@146262.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_size = fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 132:21:@146261.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_isWr = fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@146259.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_tag = fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 132:21:@146258.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_valid = fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 132:21:@146256.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@146240.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@146241.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@146242.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@146243.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@146244.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@146245.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@146246.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@146247.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@146248.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@146249.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@146250.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@146251.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@146252.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@146253.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@146254.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@146255.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@146176.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@146177.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@146178.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@146179.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@146180.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@146181.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@146182.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@146183.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@146184.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@146185.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@146186.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@146187.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@146188.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@146189.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@146190.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@146191.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@146192.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@146193.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@146194.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@146195.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@146196.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@146197.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@146198.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@146199.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@146200.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@146201.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@146202.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@146203.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@146204.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@146205.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@146206.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@146207.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@146208.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@146209.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@146210.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@146211.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@146212.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@146213.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@146214.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@146215.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@146216.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@146217.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@146218.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@146219.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@146220.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@146221.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@146222.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@146223.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@146224.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@146225.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@146226.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@146227.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@146228.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@146229.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@146230.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@146231.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@146232.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@146233.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@146234.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@146235.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@146236.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@146237.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@146238.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@146239.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wlast = fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@146175.4]
  assign MAGToAXI4Bridge_3_io_in_rresp_ready = fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 132:21:@146174.4]
  assign MAGToAXI4Bridge_3_io_in_wresp_ready = fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 132:21:@146155.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_AWREADY = io_M_AXI_3_AWREADY; // @[FringeZynq.scala 133:10:@146294.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_ARREADY = io_M_AXI_3_ARREADY; // @[FringeZynq.scala 133:10:@146282.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_WREADY = io_M_AXI_3_WREADY; // @[FringeZynq.scala 133:10:@146277.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BID = io_M_AXI_3_BID; // @[FringeZynq.scala 133:10:@146269.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BVALID = io_M_AXI_3_BVALID; // @[FringeZynq.scala 133:10:@146266.4]
endmodule
module SpatialIP( // @[:@146307.2]
  input          clock, // @[:@146308.4]
  input          reset, // @[:@146309.4]
  input          io_raddr, // @[:@146310.4]
  input          io_wen, // @[:@146310.4]
  input          io_waddr, // @[:@146310.4]
  input          io_wdata, // @[:@146310.4]
  output         io_rdata, // @[:@146310.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@146310.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@146310.4]
  input          io_S_AXI_AWVALID, // @[:@146310.4]
  output         io_S_AXI_AWREADY, // @[:@146310.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@146310.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@146310.4]
  input          io_S_AXI_ARVALID, // @[:@146310.4]
  output         io_S_AXI_ARREADY, // @[:@146310.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@146310.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@146310.4]
  input          io_S_AXI_WVALID, // @[:@146310.4]
  output         io_S_AXI_WREADY, // @[:@146310.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@146310.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@146310.4]
  output         io_S_AXI_RVALID, // @[:@146310.4]
  input          io_S_AXI_RREADY, // @[:@146310.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@146310.4]
  output         io_S_AXI_BVALID, // @[:@146310.4]
  input          io_S_AXI_BREADY, // @[:@146310.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@146310.4]
  output [31:0]  io_M_AXI_0_AWUSER, // @[:@146310.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@146310.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@146310.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@146310.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@146310.4]
  output         io_M_AXI_0_AWLOCK, // @[:@146310.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@146310.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@146310.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@146310.4]
  output         io_M_AXI_0_AWVALID, // @[:@146310.4]
  input          io_M_AXI_0_AWREADY, // @[:@146310.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@146310.4]
  output [31:0]  io_M_AXI_0_ARUSER, // @[:@146310.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@146310.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@146310.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@146310.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@146310.4]
  output         io_M_AXI_0_ARLOCK, // @[:@146310.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@146310.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@146310.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@146310.4]
  output         io_M_AXI_0_ARVALID, // @[:@146310.4]
  input          io_M_AXI_0_ARREADY, // @[:@146310.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@146310.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@146310.4]
  output         io_M_AXI_0_WLAST, // @[:@146310.4]
  output         io_M_AXI_0_WVALID, // @[:@146310.4]
  input          io_M_AXI_0_WREADY, // @[:@146310.4]
  input  [31:0]  io_M_AXI_0_RID, // @[:@146310.4]
  input  [31:0]  io_M_AXI_0_RUSER, // @[:@146310.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@146310.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@146310.4]
  input          io_M_AXI_0_RLAST, // @[:@146310.4]
  input          io_M_AXI_0_RVALID, // @[:@146310.4]
  output         io_M_AXI_0_RREADY, // @[:@146310.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@146310.4]
  input  [31:0]  io_M_AXI_0_BUSER, // @[:@146310.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@146310.4]
  input          io_M_AXI_0_BVALID, // @[:@146310.4]
  output         io_M_AXI_0_BREADY, // @[:@146310.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@146310.4]
  output [31:0]  io_M_AXI_1_AWUSER, // @[:@146310.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@146310.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@146310.4]
  output [2:0]   io_M_AXI_1_AWSIZE, // @[:@146310.4]
  output [1:0]   io_M_AXI_1_AWBURST, // @[:@146310.4]
  output         io_M_AXI_1_AWLOCK, // @[:@146310.4]
  output [3:0]   io_M_AXI_1_AWCACHE, // @[:@146310.4]
  output [2:0]   io_M_AXI_1_AWPROT, // @[:@146310.4]
  output [3:0]   io_M_AXI_1_AWQOS, // @[:@146310.4]
  output         io_M_AXI_1_AWVALID, // @[:@146310.4]
  input          io_M_AXI_1_AWREADY, // @[:@146310.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@146310.4]
  output [31:0]  io_M_AXI_1_ARUSER, // @[:@146310.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@146310.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@146310.4]
  output [2:0]   io_M_AXI_1_ARSIZE, // @[:@146310.4]
  output [1:0]   io_M_AXI_1_ARBURST, // @[:@146310.4]
  output         io_M_AXI_1_ARLOCK, // @[:@146310.4]
  output [3:0]   io_M_AXI_1_ARCACHE, // @[:@146310.4]
  output [2:0]   io_M_AXI_1_ARPROT, // @[:@146310.4]
  output [3:0]   io_M_AXI_1_ARQOS, // @[:@146310.4]
  output         io_M_AXI_1_ARVALID, // @[:@146310.4]
  input          io_M_AXI_1_ARREADY, // @[:@146310.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@146310.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@146310.4]
  output         io_M_AXI_1_WLAST, // @[:@146310.4]
  output         io_M_AXI_1_WVALID, // @[:@146310.4]
  input          io_M_AXI_1_WREADY, // @[:@146310.4]
  input  [31:0]  io_M_AXI_1_RID, // @[:@146310.4]
  input  [31:0]  io_M_AXI_1_RUSER, // @[:@146310.4]
  input  [511:0] io_M_AXI_1_RDATA, // @[:@146310.4]
  input  [1:0]   io_M_AXI_1_RRESP, // @[:@146310.4]
  input          io_M_AXI_1_RLAST, // @[:@146310.4]
  input          io_M_AXI_1_RVALID, // @[:@146310.4]
  output         io_M_AXI_1_RREADY, // @[:@146310.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@146310.4]
  input  [31:0]  io_M_AXI_1_BUSER, // @[:@146310.4]
  input  [1:0]   io_M_AXI_1_BRESP, // @[:@146310.4]
  input          io_M_AXI_1_BVALID, // @[:@146310.4]
  output         io_M_AXI_1_BREADY, // @[:@146310.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@146310.4]
  output [31:0]  io_M_AXI_2_AWUSER, // @[:@146310.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@146310.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@146310.4]
  output [2:0]   io_M_AXI_2_AWSIZE, // @[:@146310.4]
  output [1:0]   io_M_AXI_2_AWBURST, // @[:@146310.4]
  output         io_M_AXI_2_AWLOCK, // @[:@146310.4]
  output [3:0]   io_M_AXI_2_AWCACHE, // @[:@146310.4]
  output [2:0]   io_M_AXI_2_AWPROT, // @[:@146310.4]
  output [3:0]   io_M_AXI_2_AWQOS, // @[:@146310.4]
  output         io_M_AXI_2_AWVALID, // @[:@146310.4]
  input          io_M_AXI_2_AWREADY, // @[:@146310.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@146310.4]
  output [31:0]  io_M_AXI_2_ARUSER, // @[:@146310.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@146310.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@146310.4]
  output [2:0]   io_M_AXI_2_ARSIZE, // @[:@146310.4]
  output [1:0]   io_M_AXI_2_ARBURST, // @[:@146310.4]
  output         io_M_AXI_2_ARLOCK, // @[:@146310.4]
  output [3:0]   io_M_AXI_2_ARCACHE, // @[:@146310.4]
  output [2:0]   io_M_AXI_2_ARPROT, // @[:@146310.4]
  output [3:0]   io_M_AXI_2_ARQOS, // @[:@146310.4]
  output         io_M_AXI_2_ARVALID, // @[:@146310.4]
  input          io_M_AXI_2_ARREADY, // @[:@146310.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@146310.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@146310.4]
  output         io_M_AXI_2_WLAST, // @[:@146310.4]
  output         io_M_AXI_2_WVALID, // @[:@146310.4]
  input          io_M_AXI_2_WREADY, // @[:@146310.4]
  input  [31:0]  io_M_AXI_2_RID, // @[:@146310.4]
  input  [31:0]  io_M_AXI_2_RUSER, // @[:@146310.4]
  input  [511:0] io_M_AXI_2_RDATA, // @[:@146310.4]
  input  [1:0]   io_M_AXI_2_RRESP, // @[:@146310.4]
  input          io_M_AXI_2_RLAST, // @[:@146310.4]
  input          io_M_AXI_2_RVALID, // @[:@146310.4]
  output         io_M_AXI_2_RREADY, // @[:@146310.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@146310.4]
  input  [31:0]  io_M_AXI_2_BUSER, // @[:@146310.4]
  input  [1:0]   io_M_AXI_2_BRESP, // @[:@146310.4]
  input          io_M_AXI_2_BVALID, // @[:@146310.4]
  output         io_M_AXI_2_BREADY, // @[:@146310.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@146310.4]
  output [31:0]  io_M_AXI_3_AWUSER, // @[:@146310.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@146310.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@146310.4]
  output [2:0]   io_M_AXI_3_AWSIZE, // @[:@146310.4]
  output [1:0]   io_M_AXI_3_AWBURST, // @[:@146310.4]
  output         io_M_AXI_3_AWLOCK, // @[:@146310.4]
  output [3:0]   io_M_AXI_3_AWCACHE, // @[:@146310.4]
  output [2:0]   io_M_AXI_3_AWPROT, // @[:@146310.4]
  output [3:0]   io_M_AXI_3_AWQOS, // @[:@146310.4]
  output         io_M_AXI_3_AWVALID, // @[:@146310.4]
  input          io_M_AXI_3_AWREADY, // @[:@146310.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@146310.4]
  output [31:0]  io_M_AXI_3_ARUSER, // @[:@146310.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@146310.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@146310.4]
  output [2:0]   io_M_AXI_3_ARSIZE, // @[:@146310.4]
  output [1:0]   io_M_AXI_3_ARBURST, // @[:@146310.4]
  output         io_M_AXI_3_ARLOCK, // @[:@146310.4]
  output [3:0]   io_M_AXI_3_ARCACHE, // @[:@146310.4]
  output [2:0]   io_M_AXI_3_ARPROT, // @[:@146310.4]
  output [3:0]   io_M_AXI_3_ARQOS, // @[:@146310.4]
  output         io_M_AXI_3_ARVALID, // @[:@146310.4]
  input          io_M_AXI_3_ARREADY, // @[:@146310.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@146310.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@146310.4]
  output         io_M_AXI_3_WLAST, // @[:@146310.4]
  output         io_M_AXI_3_WVALID, // @[:@146310.4]
  input          io_M_AXI_3_WREADY, // @[:@146310.4]
  input  [31:0]  io_M_AXI_3_RID, // @[:@146310.4]
  input  [31:0]  io_M_AXI_3_RUSER, // @[:@146310.4]
  input  [511:0] io_M_AXI_3_RDATA, // @[:@146310.4]
  input  [1:0]   io_M_AXI_3_RRESP, // @[:@146310.4]
  input          io_M_AXI_3_RLAST, // @[:@146310.4]
  input          io_M_AXI_3_RVALID, // @[:@146310.4]
  output         io_M_AXI_3_RREADY, // @[:@146310.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@146310.4]
  input  [31:0]  io_M_AXI_3_BUSER, // @[:@146310.4]
  input  [1:0]   io_M_AXI_3_BRESP, // @[:@146310.4]
  input          io_M_AXI_3_BVALID, // @[:@146310.4]
  output         io_M_AXI_3_BREADY, // @[:@146310.4]
  input          io_TOP_AXI_AWID, // @[:@146310.4]
  input          io_TOP_AXI_AWUSER, // @[:@146310.4]
  input  [31:0]  io_TOP_AXI_AWADDR, // @[:@146310.4]
  input  [7:0]   io_TOP_AXI_AWLEN, // @[:@146310.4]
  input  [2:0]   io_TOP_AXI_AWSIZE, // @[:@146310.4]
  input  [1:0]   io_TOP_AXI_AWBURST, // @[:@146310.4]
  input          io_TOP_AXI_AWLOCK, // @[:@146310.4]
  input  [3:0]   io_TOP_AXI_AWCACHE, // @[:@146310.4]
  input  [2:0]   io_TOP_AXI_AWPROT, // @[:@146310.4]
  input  [3:0]   io_TOP_AXI_AWQOS, // @[:@146310.4]
  input          io_TOP_AXI_AWVALID, // @[:@146310.4]
  input          io_TOP_AXI_AWREADY, // @[:@146310.4]
  input          io_TOP_AXI_ARID, // @[:@146310.4]
  input          io_TOP_AXI_ARUSER, // @[:@146310.4]
  input  [31:0]  io_TOP_AXI_ARADDR, // @[:@146310.4]
  input  [7:0]   io_TOP_AXI_ARLEN, // @[:@146310.4]
  input  [2:0]   io_TOP_AXI_ARSIZE, // @[:@146310.4]
  input  [1:0]   io_TOP_AXI_ARBURST, // @[:@146310.4]
  input          io_TOP_AXI_ARLOCK, // @[:@146310.4]
  input  [3:0]   io_TOP_AXI_ARCACHE, // @[:@146310.4]
  input  [2:0]   io_TOP_AXI_ARPROT, // @[:@146310.4]
  input  [3:0]   io_TOP_AXI_ARQOS, // @[:@146310.4]
  input          io_TOP_AXI_ARVALID, // @[:@146310.4]
  input          io_TOP_AXI_ARREADY, // @[:@146310.4]
  input  [31:0]  io_TOP_AXI_WDATA, // @[:@146310.4]
  input  [63:0]  io_TOP_AXI_WSTRB, // @[:@146310.4]
  input          io_TOP_AXI_WLAST, // @[:@146310.4]
  input          io_TOP_AXI_WVALID, // @[:@146310.4]
  input          io_TOP_AXI_WREADY, // @[:@146310.4]
  input          io_TOP_AXI_RID, // @[:@146310.4]
  input          io_TOP_AXI_RUSER, // @[:@146310.4]
  input  [31:0]  io_TOP_AXI_RDATA, // @[:@146310.4]
  input  [1:0]   io_TOP_AXI_RRESP, // @[:@146310.4]
  input          io_TOP_AXI_RLAST, // @[:@146310.4]
  input          io_TOP_AXI_RVALID, // @[:@146310.4]
  input          io_TOP_AXI_RREADY, // @[:@146310.4]
  input          io_TOP_AXI_BID, // @[:@146310.4]
  input          io_TOP_AXI_BUSER, // @[:@146310.4]
  input  [1:0]   io_TOP_AXI_BRESP, // @[:@146310.4]
  input          io_TOP_AXI_BVALID, // @[:@146310.4]
  input          io_TOP_AXI_BREADY, // @[:@146310.4]
  input          io_DWIDTH_AXI_AWID, // @[:@146310.4]
  input          io_DWIDTH_AXI_AWUSER, // @[:@146310.4]
  input  [31:0]  io_DWIDTH_AXI_AWADDR, // @[:@146310.4]
  input  [7:0]   io_DWIDTH_AXI_AWLEN, // @[:@146310.4]
  input  [2:0]   io_DWIDTH_AXI_AWSIZE, // @[:@146310.4]
  input  [1:0]   io_DWIDTH_AXI_AWBURST, // @[:@146310.4]
  input          io_DWIDTH_AXI_AWLOCK, // @[:@146310.4]
  input  [3:0]   io_DWIDTH_AXI_AWCACHE, // @[:@146310.4]
  input  [2:0]   io_DWIDTH_AXI_AWPROT, // @[:@146310.4]
  input  [3:0]   io_DWIDTH_AXI_AWQOS, // @[:@146310.4]
  input          io_DWIDTH_AXI_AWVALID, // @[:@146310.4]
  input          io_DWIDTH_AXI_AWREADY, // @[:@146310.4]
  input          io_DWIDTH_AXI_ARID, // @[:@146310.4]
  input          io_DWIDTH_AXI_ARUSER, // @[:@146310.4]
  input  [31:0]  io_DWIDTH_AXI_ARADDR, // @[:@146310.4]
  input  [7:0]   io_DWIDTH_AXI_ARLEN, // @[:@146310.4]
  input  [2:0]   io_DWIDTH_AXI_ARSIZE, // @[:@146310.4]
  input  [1:0]   io_DWIDTH_AXI_ARBURST, // @[:@146310.4]
  input          io_DWIDTH_AXI_ARLOCK, // @[:@146310.4]
  input  [3:0]   io_DWIDTH_AXI_ARCACHE, // @[:@146310.4]
  input  [2:0]   io_DWIDTH_AXI_ARPROT, // @[:@146310.4]
  input  [3:0]   io_DWIDTH_AXI_ARQOS, // @[:@146310.4]
  input          io_DWIDTH_AXI_ARVALID, // @[:@146310.4]
  input          io_DWIDTH_AXI_ARREADY, // @[:@146310.4]
  input  [31:0]  io_DWIDTH_AXI_WDATA, // @[:@146310.4]
  input  [63:0]  io_DWIDTH_AXI_WSTRB, // @[:@146310.4]
  input          io_DWIDTH_AXI_WLAST, // @[:@146310.4]
  input          io_DWIDTH_AXI_WVALID, // @[:@146310.4]
  input          io_DWIDTH_AXI_WREADY, // @[:@146310.4]
  input          io_DWIDTH_AXI_RID, // @[:@146310.4]
  input          io_DWIDTH_AXI_RUSER, // @[:@146310.4]
  input  [31:0]  io_DWIDTH_AXI_RDATA, // @[:@146310.4]
  input  [1:0]   io_DWIDTH_AXI_RRESP, // @[:@146310.4]
  input          io_DWIDTH_AXI_RLAST, // @[:@146310.4]
  input          io_DWIDTH_AXI_RVALID, // @[:@146310.4]
  input          io_DWIDTH_AXI_RREADY, // @[:@146310.4]
  input          io_DWIDTH_AXI_BID, // @[:@146310.4]
  input          io_DWIDTH_AXI_BUSER, // @[:@146310.4]
  input  [1:0]   io_DWIDTH_AXI_BRESP, // @[:@146310.4]
  input          io_DWIDTH_AXI_BVALID, // @[:@146310.4]
  input          io_DWIDTH_AXI_BREADY, // @[:@146310.4]
  input          io_PROTOCOL_AXI_AWID, // @[:@146310.4]
  input          io_PROTOCOL_AXI_AWUSER, // @[:@146310.4]
  input  [31:0]  io_PROTOCOL_AXI_AWADDR, // @[:@146310.4]
  input  [7:0]   io_PROTOCOL_AXI_AWLEN, // @[:@146310.4]
  input  [2:0]   io_PROTOCOL_AXI_AWSIZE, // @[:@146310.4]
  input  [1:0]   io_PROTOCOL_AXI_AWBURST, // @[:@146310.4]
  input          io_PROTOCOL_AXI_AWLOCK, // @[:@146310.4]
  input  [3:0]   io_PROTOCOL_AXI_AWCACHE, // @[:@146310.4]
  input  [2:0]   io_PROTOCOL_AXI_AWPROT, // @[:@146310.4]
  input  [3:0]   io_PROTOCOL_AXI_AWQOS, // @[:@146310.4]
  input          io_PROTOCOL_AXI_AWVALID, // @[:@146310.4]
  input          io_PROTOCOL_AXI_AWREADY, // @[:@146310.4]
  input          io_PROTOCOL_AXI_ARID, // @[:@146310.4]
  input          io_PROTOCOL_AXI_ARUSER, // @[:@146310.4]
  input  [31:0]  io_PROTOCOL_AXI_ARADDR, // @[:@146310.4]
  input  [7:0]   io_PROTOCOL_AXI_ARLEN, // @[:@146310.4]
  input  [2:0]   io_PROTOCOL_AXI_ARSIZE, // @[:@146310.4]
  input  [1:0]   io_PROTOCOL_AXI_ARBURST, // @[:@146310.4]
  input          io_PROTOCOL_AXI_ARLOCK, // @[:@146310.4]
  input  [3:0]   io_PROTOCOL_AXI_ARCACHE, // @[:@146310.4]
  input  [2:0]   io_PROTOCOL_AXI_ARPROT, // @[:@146310.4]
  input  [3:0]   io_PROTOCOL_AXI_ARQOS, // @[:@146310.4]
  input          io_PROTOCOL_AXI_ARVALID, // @[:@146310.4]
  input          io_PROTOCOL_AXI_ARREADY, // @[:@146310.4]
  input  [31:0]  io_PROTOCOL_AXI_WDATA, // @[:@146310.4]
  input  [63:0]  io_PROTOCOL_AXI_WSTRB, // @[:@146310.4]
  input          io_PROTOCOL_AXI_WLAST, // @[:@146310.4]
  input          io_PROTOCOL_AXI_WVALID, // @[:@146310.4]
  input          io_PROTOCOL_AXI_WREADY, // @[:@146310.4]
  input          io_PROTOCOL_AXI_RID, // @[:@146310.4]
  input          io_PROTOCOL_AXI_RUSER, // @[:@146310.4]
  input  [31:0]  io_PROTOCOL_AXI_RDATA, // @[:@146310.4]
  input  [1:0]   io_PROTOCOL_AXI_RRESP, // @[:@146310.4]
  input          io_PROTOCOL_AXI_RLAST, // @[:@146310.4]
  input          io_PROTOCOL_AXI_RVALID, // @[:@146310.4]
  input          io_PROTOCOL_AXI_RREADY, // @[:@146310.4]
  input          io_PROTOCOL_AXI_BID, // @[:@146310.4]
  input          io_PROTOCOL_AXI_BUSER, // @[:@146310.4]
  input  [1:0]   io_PROTOCOL_AXI_BRESP, // @[:@146310.4]
  input          io_PROTOCOL_AXI_BVALID, // @[:@146310.4]
  input          io_PROTOCOL_AXI_BREADY, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_AWID, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_AWUSER, // @[:@146310.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_AWADDR, // @[:@146310.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_AWLEN, // @[:@146310.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWSIZE, // @[:@146310.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_AWBURST, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_AWLOCK, // @[:@146310.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWCACHE, // @[:@146310.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWPROT, // @[:@146310.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWQOS, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_AWVALID, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_AWREADY, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_ARID, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_ARUSER, // @[:@146310.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_ARADDR, // @[:@146310.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_ARLEN, // @[:@146310.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARSIZE, // @[:@146310.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_ARBURST, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_ARLOCK, // @[:@146310.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARCACHE, // @[:@146310.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARPROT, // @[:@146310.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARQOS, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_ARVALID, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_ARREADY, // @[:@146310.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_WDATA, // @[:@146310.4]
  input  [63:0]  io_CLOCKCONVERT_AXI_WSTRB, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_WLAST, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_WVALID, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_WREADY, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_RID, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_RUSER, // @[:@146310.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_RDATA, // @[:@146310.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_RRESP, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_RLAST, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_RVALID, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_RREADY, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_BID, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_BUSER, // @[:@146310.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_BRESP, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_BVALID, // @[:@146310.4]
  input          io_CLOCKCONVERT_AXI_BREADY // @[:@146310.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@146312.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@146312.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@146312.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@146312.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@146312.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@146312.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@146312.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@146312.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@146312.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@146312.4]
  wire  FringeZynq_clock; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_reset; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_S_AXI_AWADDR; // @[Zynq.scala 18:24:@146454.4]
  wire [2:0] FringeZynq_io_S_AXI_AWPROT; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_S_AXI_AWVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_S_AXI_ARADDR; // @[Zynq.scala 18:24:@146454.4]
  wire [2:0] FringeZynq_io_S_AXI_ARPROT; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_S_AXI_ARVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_S_AXI_WDATA; // @[Zynq.scala 18:24:@146454.4]
  wire [3:0] FringeZynq_io_S_AXI_WSTRB; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_S_AXI_WVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 18:24:@146454.4]
  wire [1:0] FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_S_AXI_RREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [1:0] FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_S_AXI_BREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 18:24:@146454.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_0_AWREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 18:24:@146454.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_0_ARREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [511:0] FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 18:24:@146454.4]
  wire [63:0] FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_0_WREADY; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_0_BID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_0_BVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 18:24:@146454.4]
  wire [7:0] FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_1_AWREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 18:24:@146454.4]
  wire [7:0] FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_1_ARREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [511:0] FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 18:24:@146454.4]
  wire [63:0] FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_1_WREADY; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_1_BID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_1_BVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 18:24:@146454.4]
  wire [7:0] FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_2_AWREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 18:24:@146454.4]
  wire [7:0] FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_2_ARREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [511:0] FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 18:24:@146454.4]
  wire [63:0] FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_2_WREADY; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_2_BID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_2_BVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 18:24:@146454.4]
  wire [7:0] FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_3_AWREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 18:24:@146454.4]
  wire [7:0] FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_3_ARREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [511:0] FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 18:24:@146454.4]
  wire [63:0] FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_3_WREADY; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_M_AXI_3_BID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_3_BVALID; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_enable; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_done; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_reset; // @[Zynq.scala 18:24:@146454.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[Zynq.scala 18:24:@146454.4]
  wire [63:0] FringeZynq_io_argIns_1; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[Zynq.scala 18:24:@146454.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 18:24:@146454.4]
  wire [63:0] FringeZynq_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_memStreams_stores_0_data_valid; // @[Zynq.scala 18:24:@146454.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_heap_0_req_valid; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 18:24:@146454.4]
  wire [63:0] FringeZynq_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 18:24:@146454.4]
  wire  FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 18:24:@146454.4]
  wire [63:0] FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 18:24:@146454.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@146312.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  FringeZynq FringeZynq ( // @[Zynq.scala 18:24:@146454.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWID(FringeZynq_io_M_AXI_0_AWID),
    .io_M_AXI_0_AWADDR(FringeZynq_io_M_AXI_0_AWADDR),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_AWVALID(FringeZynq_io_M_AXI_0_AWVALID),
    .io_M_AXI_0_AWREADY(FringeZynq_io_M_AXI_0_AWREADY),
    .io_M_AXI_0_ARID(FringeZynq_io_M_AXI_0_ARID),
    .io_M_AXI_0_ARADDR(FringeZynq_io_M_AXI_0_ARADDR),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_M_AXI_0_ARVALID(FringeZynq_io_M_AXI_0_ARVALID),
    .io_M_AXI_0_ARREADY(FringeZynq_io_M_AXI_0_ARREADY),
    .io_M_AXI_0_WDATA(FringeZynq_io_M_AXI_0_WDATA),
    .io_M_AXI_0_WSTRB(FringeZynq_io_M_AXI_0_WSTRB),
    .io_M_AXI_0_WLAST(FringeZynq_io_M_AXI_0_WLAST),
    .io_M_AXI_0_WVALID(FringeZynq_io_M_AXI_0_WVALID),
    .io_M_AXI_0_WREADY(FringeZynq_io_M_AXI_0_WREADY),
    .io_M_AXI_0_RREADY(FringeZynq_io_M_AXI_0_RREADY),
    .io_M_AXI_0_BID(FringeZynq_io_M_AXI_0_BID),
    .io_M_AXI_0_BVALID(FringeZynq_io_M_AXI_0_BVALID),
    .io_M_AXI_0_BREADY(FringeZynq_io_M_AXI_0_BREADY),
    .io_M_AXI_1_AWID(FringeZynq_io_M_AXI_1_AWID),
    .io_M_AXI_1_AWADDR(FringeZynq_io_M_AXI_1_AWADDR),
    .io_M_AXI_1_AWLEN(FringeZynq_io_M_AXI_1_AWLEN),
    .io_M_AXI_1_AWVALID(FringeZynq_io_M_AXI_1_AWVALID),
    .io_M_AXI_1_AWREADY(FringeZynq_io_M_AXI_1_AWREADY),
    .io_M_AXI_1_ARID(FringeZynq_io_M_AXI_1_ARID),
    .io_M_AXI_1_ARADDR(FringeZynq_io_M_AXI_1_ARADDR),
    .io_M_AXI_1_ARLEN(FringeZynq_io_M_AXI_1_ARLEN),
    .io_M_AXI_1_ARVALID(FringeZynq_io_M_AXI_1_ARVALID),
    .io_M_AXI_1_ARREADY(FringeZynq_io_M_AXI_1_ARREADY),
    .io_M_AXI_1_WDATA(FringeZynq_io_M_AXI_1_WDATA),
    .io_M_AXI_1_WSTRB(FringeZynq_io_M_AXI_1_WSTRB),
    .io_M_AXI_1_WLAST(FringeZynq_io_M_AXI_1_WLAST),
    .io_M_AXI_1_WVALID(FringeZynq_io_M_AXI_1_WVALID),
    .io_M_AXI_1_WREADY(FringeZynq_io_M_AXI_1_WREADY),
    .io_M_AXI_1_RREADY(FringeZynq_io_M_AXI_1_RREADY),
    .io_M_AXI_1_BID(FringeZynq_io_M_AXI_1_BID),
    .io_M_AXI_1_BVALID(FringeZynq_io_M_AXI_1_BVALID),
    .io_M_AXI_1_BREADY(FringeZynq_io_M_AXI_1_BREADY),
    .io_M_AXI_2_AWID(FringeZynq_io_M_AXI_2_AWID),
    .io_M_AXI_2_AWADDR(FringeZynq_io_M_AXI_2_AWADDR),
    .io_M_AXI_2_AWLEN(FringeZynq_io_M_AXI_2_AWLEN),
    .io_M_AXI_2_AWVALID(FringeZynq_io_M_AXI_2_AWVALID),
    .io_M_AXI_2_AWREADY(FringeZynq_io_M_AXI_2_AWREADY),
    .io_M_AXI_2_ARID(FringeZynq_io_M_AXI_2_ARID),
    .io_M_AXI_2_ARADDR(FringeZynq_io_M_AXI_2_ARADDR),
    .io_M_AXI_2_ARLEN(FringeZynq_io_M_AXI_2_ARLEN),
    .io_M_AXI_2_ARVALID(FringeZynq_io_M_AXI_2_ARVALID),
    .io_M_AXI_2_ARREADY(FringeZynq_io_M_AXI_2_ARREADY),
    .io_M_AXI_2_WDATA(FringeZynq_io_M_AXI_2_WDATA),
    .io_M_AXI_2_WSTRB(FringeZynq_io_M_AXI_2_WSTRB),
    .io_M_AXI_2_WLAST(FringeZynq_io_M_AXI_2_WLAST),
    .io_M_AXI_2_WVALID(FringeZynq_io_M_AXI_2_WVALID),
    .io_M_AXI_2_WREADY(FringeZynq_io_M_AXI_2_WREADY),
    .io_M_AXI_2_RREADY(FringeZynq_io_M_AXI_2_RREADY),
    .io_M_AXI_2_BID(FringeZynq_io_M_AXI_2_BID),
    .io_M_AXI_2_BVALID(FringeZynq_io_M_AXI_2_BVALID),
    .io_M_AXI_2_BREADY(FringeZynq_io_M_AXI_2_BREADY),
    .io_M_AXI_3_AWID(FringeZynq_io_M_AXI_3_AWID),
    .io_M_AXI_3_AWADDR(FringeZynq_io_M_AXI_3_AWADDR),
    .io_M_AXI_3_AWLEN(FringeZynq_io_M_AXI_3_AWLEN),
    .io_M_AXI_3_AWVALID(FringeZynq_io_M_AXI_3_AWVALID),
    .io_M_AXI_3_AWREADY(FringeZynq_io_M_AXI_3_AWREADY),
    .io_M_AXI_3_ARID(FringeZynq_io_M_AXI_3_ARID),
    .io_M_AXI_3_ARADDR(FringeZynq_io_M_AXI_3_ARADDR),
    .io_M_AXI_3_ARLEN(FringeZynq_io_M_AXI_3_ARLEN),
    .io_M_AXI_3_ARVALID(FringeZynq_io_M_AXI_3_ARVALID),
    .io_M_AXI_3_ARREADY(FringeZynq_io_M_AXI_3_ARREADY),
    .io_M_AXI_3_WDATA(FringeZynq_io_M_AXI_3_WDATA),
    .io_M_AXI_3_WSTRB(FringeZynq_io_M_AXI_3_WSTRB),
    .io_M_AXI_3_WLAST(FringeZynq_io_M_AXI_3_WLAST),
    .io_M_AXI_3_WVALID(FringeZynq_io_M_AXI_3_WVALID),
    .io_M_AXI_3_WREADY(FringeZynq_io_M_AXI_3_WREADY),
    .io_M_AXI_3_RREADY(FringeZynq_io_M_AXI_3_RREADY),
    .io_M_AXI_3_BID(FringeZynq_io_M_AXI_3_BID),
    .io_M_AXI_3_BVALID(FringeZynq_io_M_AXI_3_BVALID),
    .io_M_AXI_3_BREADY(FringeZynq_io_M_AXI_3_BREADY),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argIns_1(FringeZynq_io_argIns_1),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(FringeZynq_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(FringeZynq_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(FringeZynq_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(FringeZynq_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(FringeZynq_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(FringeZynq_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(FringeZynq_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(FringeZynq_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(FringeZynq_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(FringeZynq_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(FringeZynq_io_memStreams_stores_0_wresp_bits),
    .io_heap_0_req_valid(FringeZynq_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(FringeZynq_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(FringeZynq_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(FringeZynq_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(FringeZynq_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(FringeZynq_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 21:21:@146472.4]
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 21:21:@146468.4]
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 21:21:@146464.4]
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 21:21:@146463.4]
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 21:21:@146462.4]
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 21:21:@146461.4]
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 21:21:@146459.4]
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 21:21:@146458.4]
  assign io_M_AXI_0_AWID = FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 24:14:@146516.4]
  assign io_M_AXI_0_AWUSER = 32'h0; // @[Zynq.scala 24:14:@146515.4]
  assign io_M_AXI_0_AWADDR = FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 24:14:@146514.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 24:14:@146513.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@146512.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[Zynq.scala 24:14:@146511.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@146510.4]
  assign io_M_AXI_0_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@146509.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[Zynq.scala 24:14:@146508.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[Zynq.scala 24:14:@146507.4]
  assign io_M_AXI_0_AWVALID = FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 24:14:@146506.4]
  assign io_M_AXI_0_ARID = FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 24:14:@146504.4]
  assign io_M_AXI_0_ARUSER = 32'h0; // @[Zynq.scala 24:14:@146503.4]
  assign io_M_AXI_0_ARADDR = FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 24:14:@146502.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 24:14:@146501.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@146500.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[Zynq.scala 24:14:@146499.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@146498.4]
  assign io_M_AXI_0_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@146497.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[Zynq.scala 24:14:@146496.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[Zynq.scala 24:14:@146495.4]
  assign io_M_AXI_0_ARVALID = FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 24:14:@146494.4]
  assign io_M_AXI_0_WDATA = FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 24:14:@146492.4]
  assign io_M_AXI_0_WSTRB = FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 24:14:@146491.4]
  assign io_M_AXI_0_WLAST = FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 24:14:@146490.4]
  assign io_M_AXI_0_WVALID = FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 24:14:@146489.4]
  assign io_M_AXI_0_RREADY = FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 24:14:@146481.4]
  assign io_M_AXI_0_BREADY = FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 24:14:@146476.4]
  assign io_M_AXI_1_AWID = FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 24:14:@146557.4]
  assign io_M_AXI_1_AWUSER = 32'h0; // @[Zynq.scala 24:14:@146556.4]
  assign io_M_AXI_1_AWADDR = FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 24:14:@146555.4]
  assign io_M_AXI_1_AWLEN = FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 24:14:@146554.4]
  assign io_M_AXI_1_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@146553.4]
  assign io_M_AXI_1_AWBURST = 2'h1; // @[Zynq.scala 24:14:@146552.4]
  assign io_M_AXI_1_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@146551.4]
  assign io_M_AXI_1_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@146550.4]
  assign io_M_AXI_1_AWPROT = 3'h0; // @[Zynq.scala 24:14:@146549.4]
  assign io_M_AXI_1_AWQOS = 4'h0; // @[Zynq.scala 24:14:@146548.4]
  assign io_M_AXI_1_AWVALID = FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 24:14:@146547.4]
  assign io_M_AXI_1_ARID = FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 24:14:@146545.4]
  assign io_M_AXI_1_ARUSER = 32'h0; // @[Zynq.scala 24:14:@146544.4]
  assign io_M_AXI_1_ARADDR = FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 24:14:@146543.4]
  assign io_M_AXI_1_ARLEN = FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 24:14:@146542.4]
  assign io_M_AXI_1_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@146541.4]
  assign io_M_AXI_1_ARBURST = 2'h1; // @[Zynq.scala 24:14:@146540.4]
  assign io_M_AXI_1_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@146539.4]
  assign io_M_AXI_1_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@146538.4]
  assign io_M_AXI_1_ARPROT = 3'h0; // @[Zynq.scala 24:14:@146537.4]
  assign io_M_AXI_1_ARQOS = 4'h0; // @[Zynq.scala 24:14:@146536.4]
  assign io_M_AXI_1_ARVALID = FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 24:14:@146535.4]
  assign io_M_AXI_1_WDATA = FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 24:14:@146533.4]
  assign io_M_AXI_1_WSTRB = FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 24:14:@146532.4]
  assign io_M_AXI_1_WLAST = FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 24:14:@146531.4]
  assign io_M_AXI_1_WVALID = FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 24:14:@146530.4]
  assign io_M_AXI_1_RREADY = FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 24:14:@146522.4]
  assign io_M_AXI_1_BREADY = FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 24:14:@146517.4]
  assign io_M_AXI_2_AWID = FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 24:14:@146598.4]
  assign io_M_AXI_2_AWUSER = 32'h0; // @[Zynq.scala 24:14:@146597.4]
  assign io_M_AXI_2_AWADDR = FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 24:14:@146596.4]
  assign io_M_AXI_2_AWLEN = FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 24:14:@146595.4]
  assign io_M_AXI_2_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@146594.4]
  assign io_M_AXI_2_AWBURST = 2'h1; // @[Zynq.scala 24:14:@146593.4]
  assign io_M_AXI_2_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@146592.4]
  assign io_M_AXI_2_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@146591.4]
  assign io_M_AXI_2_AWPROT = 3'h0; // @[Zynq.scala 24:14:@146590.4]
  assign io_M_AXI_2_AWQOS = 4'h0; // @[Zynq.scala 24:14:@146589.4]
  assign io_M_AXI_2_AWVALID = FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 24:14:@146588.4]
  assign io_M_AXI_2_ARID = FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 24:14:@146586.4]
  assign io_M_AXI_2_ARUSER = 32'h0; // @[Zynq.scala 24:14:@146585.4]
  assign io_M_AXI_2_ARADDR = FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 24:14:@146584.4]
  assign io_M_AXI_2_ARLEN = FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 24:14:@146583.4]
  assign io_M_AXI_2_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@146582.4]
  assign io_M_AXI_2_ARBURST = 2'h1; // @[Zynq.scala 24:14:@146581.4]
  assign io_M_AXI_2_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@146580.4]
  assign io_M_AXI_2_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@146579.4]
  assign io_M_AXI_2_ARPROT = 3'h0; // @[Zynq.scala 24:14:@146578.4]
  assign io_M_AXI_2_ARQOS = 4'h0; // @[Zynq.scala 24:14:@146577.4]
  assign io_M_AXI_2_ARVALID = FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 24:14:@146576.4]
  assign io_M_AXI_2_WDATA = FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 24:14:@146574.4]
  assign io_M_AXI_2_WSTRB = FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 24:14:@146573.4]
  assign io_M_AXI_2_WLAST = FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 24:14:@146572.4]
  assign io_M_AXI_2_WVALID = FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 24:14:@146571.4]
  assign io_M_AXI_2_RREADY = FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 24:14:@146563.4]
  assign io_M_AXI_2_BREADY = FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 24:14:@146558.4]
  assign io_M_AXI_3_AWID = FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 24:14:@146639.4]
  assign io_M_AXI_3_AWUSER = 32'h0; // @[Zynq.scala 24:14:@146638.4]
  assign io_M_AXI_3_AWADDR = FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 24:14:@146637.4]
  assign io_M_AXI_3_AWLEN = FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 24:14:@146636.4]
  assign io_M_AXI_3_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@146635.4]
  assign io_M_AXI_3_AWBURST = 2'h1; // @[Zynq.scala 24:14:@146634.4]
  assign io_M_AXI_3_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@146633.4]
  assign io_M_AXI_3_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@146632.4]
  assign io_M_AXI_3_AWPROT = 3'h0; // @[Zynq.scala 24:14:@146631.4]
  assign io_M_AXI_3_AWQOS = 4'h0; // @[Zynq.scala 24:14:@146630.4]
  assign io_M_AXI_3_AWVALID = FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 24:14:@146629.4]
  assign io_M_AXI_3_ARID = FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 24:14:@146627.4]
  assign io_M_AXI_3_ARUSER = 32'h0; // @[Zynq.scala 24:14:@146626.4]
  assign io_M_AXI_3_ARADDR = FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 24:14:@146625.4]
  assign io_M_AXI_3_ARLEN = FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 24:14:@146624.4]
  assign io_M_AXI_3_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@146623.4]
  assign io_M_AXI_3_ARBURST = 2'h1; // @[Zynq.scala 24:14:@146622.4]
  assign io_M_AXI_3_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@146621.4]
  assign io_M_AXI_3_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@146620.4]
  assign io_M_AXI_3_ARPROT = 3'h0; // @[Zynq.scala 24:14:@146619.4]
  assign io_M_AXI_3_ARQOS = 4'h0; // @[Zynq.scala 24:14:@146618.4]
  assign io_M_AXI_3_ARVALID = FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 24:14:@146617.4]
  assign io_M_AXI_3_WDATA = FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 24:14:@146615.4]
  assign io_M_AXI_3_WSTRB = FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 24:14:@146614.4]
  assign io_M_AXI_3_WLAST = FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 24:14:@146613.4]
  assign io_M_AXI_3_WVALID = FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 24:14:@146612.4]
  assign io_M_AXI_3_RREADY = FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 24:14:@146604.4]
  assign io_M_AXI_3_BREADY = FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 24:14:@146599.4]
  assign accel_clock = clock; // @[:@146313.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@146314.4 Zynq.scala 54:17:@146928.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[Zynq.scala 51:21:@146923.4]
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@146916.4]
  assign accel_io_memStreams_loads_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@146911.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0; // @[Zynq.scala 49:26:@146895.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0; // @[Zynq.scala 49:26:@146896.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0; // @[Zynq.scala 49:26:@146897.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0; // @[Zynq.scala 49:26:@146898.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0; // @[Zynq.scala 49:26:@146899.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0; // @[Zynq.scala 49:26:@146900.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0; // @[Zynq.scala 49:26:@146901.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0; // @[Zynq.scala 49:26:@146902.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0; // @[Zynq.scala 49:26:@146903.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0; // @[Zynq.scala 49:26:@146904.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0; // @[Zynq.scala 49:26:@146905.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0; // @[Zynq.scala 49:26:@146906.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0; // @[Zynq.scala 49:26:@146907.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0; // @[Zynq.scala 49:26:@146908.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0; // @[Zynq.scala 49:26:@146909.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0; // @[Zynq.scala 49:26:@146910.4]
  assign accel_io_memStreams_stores_0_cmd_ready = FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 49:26:@146894.4]
  assign accel_io_memStreams_stores_0_data_ready = FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 49:26:@146890.4]
  assign accel_io_memStreams_stores_0_wresp_valid = FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 49:26:@146885.4]
  assign accel_io_memStreams_stores_0_wresp_bits = FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 49:26:@146884.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@146883.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@146864.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0; // @[Zynq.scala 49:26:@146848.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0; // @[Zynq.scala 49:26:@146849.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0; // @[Zynq.scala 49:26:@146850.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0; // @[Zynq.scala 49:26:@146851.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0; // @[Zynq.scala 49:26:@146852.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0; // @[Zynq.scala 49:26:@146853.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0; // @[Zynq.scala 49:26:@146854.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0; // @[Zynq.scala 49:26:@146855.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0; // @[Zynq.scala 49:26:@146856.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0; // @[Zynq.scala 49:26:@146857.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0; // @[Zynq.scala 49:26:@146858.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0; // @[Zynq.scala 49:26:@146859.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0; // @[Zynq.scala 49:26:@146860.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0; // @[Zynq.scala 49:26:@146861.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0; // @[Zynq.scala 49:26:@146862.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0; // @[Zynq.scala 49:26:@146863.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@146847.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[Zynq.scala 49:26:@146812.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[Zynq.scala 49:26:@146811.4]
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 50:20:@146919.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 50:20:@146918.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 50:20:@146917.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[Zynq.scala 34:21:@146805.4]
  assign accel_io_argIns_1 = FringeZynq_io_argIns_1; // @[Zynq.scala 34:21:@146806.4]
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0; // @[Zynq.scala 40:24:@146809.4]
  assign FringeZynq_clock = clock; // @[:@146455.4]
  assign FringeZynq_reset = reset == 1'h0; // @[:@146456.4 Zynq.scala 53:18:@146927.4]
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[Zynq.scala 21:21:@146475.4]
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[Zynq.scala 21:21:@146474.4]
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[Zynq.scala 21:21:@146473.4]
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[Zynq.scala 21:21:@146471.4]
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[Zynq.scala 21:21:@146470.4]
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[Zynq.scala 21:21:@146469.4]
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[Zynq.scala 21:21:@146467.4]
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[Zynq.scala 21:21:@146466.4]
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[Zynq.scala 21:21:@146465.4]
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[Zynq.scala 21:21:@146460.4]
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[Zynq.scala 21:21:@146457.4]
  assign FringeZynq_io_M_AXI_0_AWREADY = io_M_AXI_0_AWREADY; // @[Zynq.scala 24:14:@146505.4]
  assign FringeZynq_io_M_AXI_0_ARREADY = io_M_AXI_0_ARREADY; // @[Zynq.scala 24:14:@146493.4]
  assign FringeZynq_io_M_AXI_0_WREADY = io_M_AXI_0_WREADY; // @[Zynq.scala 24:14:@146488.4]
  assign FringeZynq_io_M_AXI_0_BID = io_M_AXI_0_BID; // @[Zynq.scala 24:14:@146480.4]
  assign FringeZynq_io_M_AXI_0_BVALID = io_M_AXI_0_BVALID; // @[Zynq.scala 24:14:@146477.4]
  assign FringeZynq_io_M_AXI_1_AWREADY = io_M_AXI_1_AWREADY; // @[Zynq.scala 24:14:@146546.4]
  assign FringeZynq_io_M_AXI_1_ARREADY = io_M_AXI_1_ARREADY; // @[Zynq.scala 24:14:@146534.4]
  assign FringeZynq_io_M_AXI_1_WREADY = io_M_AXI_1_WREADY; // @[Zynq.scala 24:14:@146529.4]
  assign FringeZynq_io_M_AXI_1_BID = io_M_AXI_1_BID; // @[Zynq.scala 24:14:@146521.4]
  assign FringeZynq_io_M_AXI_1_BVALID = io_M_AXI_1_BVALID; // @[Zynq.scala 24:14:@146518.4]
  assign FringeZynq_io_M_AXI_2_AWREADY = io_M_AXI_2_AWREADY; // @[Zynq.scala 24:14:@146587.4]
  assign FringeZynq_io_M_AXI_2_ARREADY = io_M_AXI_2_ARREADY; // @[Zynq.scala 24:14:@146575.4]
  assign FringeZynq_io_M_AXI_2_WREADY = io_M_AXI_2_WREADY; // @[Zynq.scala 24:14:@146570.4]
  assign FringeZynq_io_M_AXI_2_BID = io_M_AXI_2_BID; // @[Zynq.scala 24:14:@146562.4]
  assign FringeZynq_io_M_AXI_2_BVALID = io_M_AXI_2_BVALID; // @[Zynq.scala 24:14:@146559.4]
  assign FringeZynq_io_M_AXI_3_AWREADY = io_M_AXI_3_AWREADY; // @[Zynq.scala 24:14:@146628.4]
  assign FringeZynq_io_M_AXI_3_ARREADY = io_M_AXI_3_ARREADY; // @[Zynq.scala 24:14:@146616.4]
  assign FringeZynq_io_M_AXI_3_WREADY = io_M_AXI_3_WREADY; // @[Zynq.scala 24:14:@146611.4]
  assign FringeZynq_io_M_AXI_3_BID = io_M_AXI_3_BID; // @[Zynq.scala 24:14:@146603.4]
  assign FringeZynq_io_M_AXI_3_BVALID = io_M_AXI_3_BVALID; // @[Zynq.scala 24:14:@146600.4]
  assign FringeZynq_io_done = accel_io_done; // @[Zynq.scala 52:20:@146924.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[Zynq.scala 37:26:@146808.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[Zynq.scala 36:25:@146807.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_valid = accel_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 49:26:@146893.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_addr = accel_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 49:26:@146892.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_size = accel_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 49:26:@146891.4]
  assign FringeZynq_io_memStreams_stores_0_data_valid = accel_io_memStreams_stores_0_data_valid; // @[Zynq.scala 49:26:@146889.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wdata_0 = accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 49:26:@146888.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wstrb = accel_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 49:26:@146887.4]
  assign FringeZynq_io_memStreams_stores_0_wresp_ready = accel_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 49:26:@146886.4]
  assign FringeZynq_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[Zynq.scala 50:20:@146922.4]
  assign FringeZynq_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 50:20:@146921.4]
  assign FringeZynq_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 50:20:@146920.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
module SRAMVerilogDualRead
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr0,
    input [AWIDTH-1:0] raddr1,
    input [AWIDTH-1:0] waddr,
    input raddrEn0,
    input raddrEn1,
    input waddrEn,
    input wen,
    input backpressure0,
    input backpressure1,
    input [DWIDTH-1:0] wdata,
    output reg [DWIDTH-1:0] rdata0,
    output reg [DWIDTH-1:0] rdata1
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk)
    begin
            if (wen)
            begin
                mem[waddr] <= wdata;
            end
            if (backpressure0) rdata0 <= mem[raddr0];
    end


    always @(posedge clk)
    begin
        if (backpressure1) rdata1 <= mem[raddr1];
    end
endmodule




