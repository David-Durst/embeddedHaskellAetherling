module FIFO(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  input  [7:0] I_4,
  input  [7:0] I_5,
  input  [7:0] I_6,
  input  [7:0] I_7,
  input  [7:0] I_8,
  input  [7:0] I_9,
  input  [7:0] I_10,
  input  [7:0] I_11,
  input  [7:0] I_12,
  input  [7:0] I_13,
  input  [7:0] I_14,
  input  [7:0] I_15,
  input  [7:0] I_16,
  input  [7:0] I_17,
  input  [7:0] I_18,
  input  [7:0] I_19,
  input  [7:0] I_20,
  input  [7:0] I_21,
  input  [7:0] I_22,
  input  [7:0] I_23,
  input  [7:0] I_24,
  input  [7:0] I_25,
  input  [7:0] I_26,
  input  [7:0] I_27,
  input  [7:0] I_28,
  input  [7:0] I_29,
  input  [7:0] I_30,
  input  [7:0] I_31,
  input  [7:0] I_32,
  input  [7:0] I_33,
  input  [7:0] I_34,
  input  [7:0] I_35,
  input  [7:0] I_36,
  input  [7:0] I_37,
  input  [7:0] I_38,
  input  [7:0] I_39,
  input  [7:0] I_40,
  input  [7:0] I_41,
  input  [7:0] I_42,
  input  [7:0] I_43,
  input  [7:0] I_44,
  input  [7:0] I_45,
  input  [7:0] I_46,
  input  [7:0] I_47,
  input  [7:0] I_48,
  input  [7:0] I_49,
  input  [7:0] I_50,
  input  [7:0] I_51,
  input  [7:0] I_52,
  input  [7:0] I_53,
  input  [7:0] I_54,
  input  [7:0] I_55,
  input  [7:0] I_56,
  input  [7:0] I_57,
  input  [7:0] I_58,
  input  [7:0] I_59,
  input  [7:0] I_60,
  input  [7:0] I_61,
  input  [7:0] I_62,
  input  [7:0] I_63,
  input  [7:0] I_64,
  input  [7:0] I_65,
  input  [7:0] I_66,
  input  [7:0] I_67,
  input  [7:0] I_68,
  input  [7:0] I_69,
  input  [7:0] I_70,
  input  [7:0] I_71,
  input  [7:0] I_72,
  input  [7:0] I_73,
  input  [7:0] I_74,
  input  [7:0] I_75,
  input  [7:0] I_76,
  input  [7:0] I_77,
  input  [7:0] I_78,
  input  [7:0] I_79,
  input  [7:0] I_80,
  input  [7:0] I_81,
  input  [7:0] I_82,
  input  [7:0] I_83,
  input  [7:0] I_84,
  input  [7:0] I_85,
  input  [7:0] I_86,
  input  [7:0] I_87,
  input  [7:0] I_88,
  input  [7:0] I_89,
  input  [7:0] I_90,
  input  [7:0] I_91,
  input  [7:0] I_92,
  input  [7:0] I_93,
  input  [7:0] I_94,
  input  [7:0] I_95,
  input  [7:0] I_96,
  input  [7:0] I_97,
  input  [7:0] I_98,
  input  [7:0] I_99,
  input  [7:0] I_100,
  input  [7:0] I_101,
  input  [7:0] I_102,
  input  [7:0] I_103,
  input  [7:0] I_104,
  input  [7:0] I_105,
  input  [7:0] I_106,
  input  [7:0] I_107,
  input  [7:0] I_108,
  input  [7:0] I_109,
  input  [7:0] I_110,
  input  [7:0] I_111,
  input  [7:0] I_112,
  input  [7:0] I_113,
  input  [7:0] I_114,
  input  [7:0] I_115,
  input  [7:0] I_116,
  input  [7:0] I_117,
  input  [7:0] I_118,
  input  [7:0] I_119,
  input  [7:0] I_120,
  input  [7:0] I_121,
  input  [7:0] I_122,
  input  [7:0] I_123,
  input  [7:0] I_124,
  input  [7:0] I_125,
  input  [7:0] I_126,
  input  [7:0] I_127,
  input  [7:0] I_128,
  input  [7:0] I_129,
  input  [7:0] I_130,
  input  [7:0] I_131,
  input  [7:0] I_132,
  input  [7:0] I_133,
  input  [7:0] I_134,
  input  [7:0] I_135,
  input  [7:0] I_136,
  input  [7:0] I_137,
  input  [7:0] I_138,
  input  [7:0] I_139,
  input  [7:0] I_140,
  input  [7:0] I_141,
  input  [7:0] I_142,
  input  [7:0] I_143,
  input  [7:0] I_144,
  input  [7:0] I_145,
  input  [7:0] I_146,
  input  [7:0] I_147,
  input  [7:0] I_148,
  input  [7:0] I_149,
  input  [7:0] I_150,
  input  [7:0] I_151,
  input  [7:0] I_152,
  input  [7:0] I_153,
  input  [7:0] I_154,
  input  [7:0] I_155,
  input  [7:0] I_156,
  input  [7:0] I_157,
  input  [7:0] I_158,
  input  [7:0] I_159,
  input  [7:0] I_160,
  input  [7:0] I_161,
  input  [7:0] I_162,
  input  [7:0] I_163,
  input  [7:0] I_164,
  input  [7:0] I_165,
  input  [7:0] I_166,
  input  [7:0] I_167,
  input  [7:0] I_168,
  input  [7:0] I_169,
  input  [7:0] I_170,
  input  [7:0] I_171,
  input  [7:0] I_172,
  input  [7:0] I_173,
  input  [7:0] I_174,
  input  [7:0] I_175,
  input  [7:0] I_176,
  input  [7:0] I_177,
  input  [7:0] I_178,
  input  [7:0] I_179,
  input  [7:0] I_180,
  input  [7:0] I_181,
  input  [7:0] I_182,
  input  [7:0] I_183,
  input  [7:0] I_184,
  input  [7:0] I_185,
  input  [7:0] I_186,
  input  [7:0] I_187,
  input  [7:0] I_188,
  input  [7:0] I_189,
  input  [7:0] I_190,
  input  [7:0] I_191,
  input  [7:0] I_192,
  input  [7:0] I_193,
  input  [7:0] I_194,
  input  [7:0] I_195,
  input  [7:0] I_196,
  input  [7:0] I_197,
  input  [7:0] I_198,
  input  [7:0] I_199,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15,
  output [7:0] O_16,
  output [7:0] O_17,
  output [7:0] O_18,
  output [7:0] O_19,
  output [7:0] O_20,
  output [7:0] O_21,
  output [7:0] O_22,
  output [7:0] O_23,
  output [7:0] O_24,
  output [7:0] O_25,
  output [7:0] O_26,
  output [7:0] O_27,
  output [7:0] O_28,
  output [7:0] O_29,
  output [7:0] O_30,
  output [7:0] O_31,
  output [7:0] O_32,
  output [7:0] O_33,
  output [7:0] O_34,
  output [7:0] O_35,
  output [7:0] O_36,
  output [7:0] O_37,
  output [7:0] O_38,
  output [7:0] O_39,
  output [7:0] O_40,
  output [7:0] O_41,
  output [7:0] O_42,
  output [7:0] O_43,
  output [7:0] O_44,
  output [7:0] O_45,
  output [7:0] O_46,
  output [7:0] O_47,
  output [7:0] O_48,
  output [7:0] O_49,
  output [7:0] O_50,
  output [7:0] O_51,
  output [7:0] O_52,
  output [7:0] O_53,
  output [7:0] O_54,
  output [7:0] O_55,
  output [7:0] O_56,
  output [7:0] O_57,
  output [7:0] O_58,
  output [7:0] O_59,
  output [7:0] O_60,
  output [7:0] O_61,
  output [7:0] O_62,
  output [7:0] O_63,
  output [7:0] O_64,
  output [7:0] O_65,
  output [7:0] O_66,
  output [7:0] O_67,
  output [7:0] O_68,
  output [7:0] O_69,
  output [7:0] O_70,
  output [7:0] O_71,
  output [7:0] O_72,
  output [7:0] O_73,
  output [7:0] O_74,
  output [7:0] O_75,
  output [7:0] O_76,
  output [7:0] O_77,
  output [7:0] O_78,
  output [7:0] O_79,
  output [7:0] O_80,
  output [7:0] O_81,
  output [7:0] O_82,
  output [7:0] O_83,
  output [7:0] O_84,
  output [7:0] O_85,
  output [7:0] O_86,
  output [7:0] O_87,
  output [7:0] O_88,
  output [7:0] O_89,
  output [7:0] O_90,
  output [7:0] O_91,
  output [7:0] O_92,
  output [7:0] O_93,
  output [7:0] O_94,
  output [7:0] O_95,
  output [7:0] O_96,
  output [7:0] O_97,
  output [7:0] O_98,
  output [7:0] O_99,
  output [7:0] O_100,
  output [7:0] O_101,
  output [7:0] O_102,
  output [7:0] O_103,
  output [7:0] O_104,
  output [7:0] O_105,
  output [7:0] O_106,
  output [7:0] O_107,
  output [7:0] O_108,
  output [7:0] O_109,
  output [7:0] O_110,
  output [7:0] O_111,
  output [7:0] O_112,
  output [7:0] O_113,
  output [7:0] O_114,
  output [7:0] O_115,
  output [7:0] O_116,
  output [7:0] O_117,
  output [7:0] O_118,
  output [7:0] O_119,
  output [7:0] O_120,
  output [7:0] O_121,
  output [7:0] O_122,
  output [7:0] O_123,
  output [7:0] O_124,
  output [7:0] O_125,
  output [7:0] O_126,
  output [7:0] O_127,
  output [7:0] O_128,
  output [7:0] O_129,
  output [7:0] O_130,
  output [7:0] O_131,
  output [7:0] O_132,
  output [7:0] O_133,
  output [7:0] O_134,
  output [7:0] O_135,
  output [7:0] O_136,
  output [7:0] O_137,
  output [7:0] O_138,
  output [7:0] O_139,
  output [7:0] O_140,
  output [7:0] O_141,
  output [7:0] O_142,
  output [7:0] O_143,
  output [7:0] O_144,
  output [7:0] O_145,
  output [7:0] O_146,
  output [7:0] O_147,
  output [7:0] O_148,
  output [7:0] O_149,
  output [7:0] O_150,
  output [7:0] O_151,
  output [7:0] O_152,
  output [7:0] O_153,
  output [7:0] O_154,
  output [7:0] O_155,
  output [7:0] O_156,
  output [7:0] O_157,
  output [7:0] O_158,
  output [7:0] O_159,
  output [7:0] O_160,
  output [7:0] O_161,
  output [7:0] O_162,
  output [7:0] O_163,
  output [7:0] O_164,
  output [7:0] O_165,
  output [7:0] O_166,
  output [7:0] O_167,
  output [7:0] O_168,
  output [7:0] O_169,
  output [7:0] O_170,
  output [7:0] O_171,
  output [7:0] O_172,
  output [7:0] O_173,
  output [7:0] O_174,
  output [7:0] O_175,
  output [7:0] O_176,
  output [7:0] O_177,
  output [7:0] O_178,
  output [7:0] O_179,
  output [7:0] O_180,
  output [7:0] O_181,
  output [7:0] O_182,
  output [7:0] O_183,
  output [7:0] O_184,
  output [7:0] O_185,
  output [7:0] O_186,
  output [7:0] O_187,
  output [7:0] O_188,
  output [7:0] O_189,
  output [7:0] O_190,
  output [7:0] O_191,
  output [7:0] O_192,
  output [7:0] O_193,
  output [7:0] O_194,
  output [7:0] O_195,
  output [7:0] O_196,
  output [7:0] O_197,
  output [7:0] O_198,
  output [7:0] O_199
);
  reg [7:0] _T__0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg [7:0] _T__1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_1;
  reg [7:0] _T__2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_2;
  reg [7:0] _T__3; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_3;
  reg [7:0] _T__4; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_4;
  reg [7:0] _T__5; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_5;
  reg [7:0] _T__6; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_6;
  reg [7:0] _T__7; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_7;
  reg [7:0] _T__8; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_8;
  reg [7:0] _T__9; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_9;
  reg [7:0] _T__10; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_10;
  reg [7:0] _T__11; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_11;
  reg [7:0] _T__12; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_12;
  reg [7:0] _T__13; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_13;
  reg [7:0] _T__14; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_14;
  reg [7:0] _T__15; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_15;
  reg [7:0] _T__16; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_16;
  reg [7:0] _T__17; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_17;
  reg [7:0] _T__18; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_18;
  reg [7:0] _T__19; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_19;
  reg [7:0] _T__20; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_20;
  reg [7:0] _T__21; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_21;
  reg [7:0] _T__22; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_22;
  reg [7:0] _T__23; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_23;
  reg [7:0] _T__24; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_24;
  reg [7:0] _T__25; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_25;
  reg [7:0] _T__26; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_26;
  reg [7:0] _T__27; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_27;
  reg [7:0] _T__28; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_28;
  reg [7:0] _T__29; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_29;
  reg [7:0] _T__30; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_30;
  reg [7:0] _T__31; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_31;
  reg [7:0] _T__32; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_32;
  reg [7:0] _T__33; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_33;
  reg [7:0] _T__34; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_34;
  reg [7:0] _T__35; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_35;
  reg [7:0] _T__36; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_36;
  reg [7:0] _T__37; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_37;
  reg [7:0] _T__38; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_38;
  reg [7:0] _T__39; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_39;
  reg [7:0] _T__40; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_40;
  reg [7:0] _T__41; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_41;
  reg [7:0] _T__42; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_42;
  reg [7:0] _T__43; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_43;
  reg [7:0] _T__44; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_44;
  reg [7:0] _T__45; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_45;
  reg [7:0] _T__46; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_46;
  reg [7:0] _T__47; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_47;
  reg [7:0] _T__48; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_48;
  reg [7:0] _T__49; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_49;
  reg [7:0] _T__50; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_50;
  reg [7:0] _T__51; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_51;
  reg [7:0] _T__52; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_52;
  reg [7:0] _T__53; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_53;
  reg [7:0] _T__54; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_54;
  reg [7:0] _T__55; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_55;
  reg [7:0] _T__56; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_56;
  reg [7:0] _T__57; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_57;
  reg [7:0] _T__58; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_58;
  reg [7:0] _T__59; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_59;
  reg [7:0] _T__60; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_60;
  reg [7:0] _T__61; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_61;
  reg [7:0] _T__62; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_62;
  reg [7:0] _T__63; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_63;
  reg [7:0] _T__64; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_64;
  reg [7:0] _T__65; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_65;
  reg [7:0] _T__66; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_66;
  reg [7:0] _T__67; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_67;
  reg [7:0] _T__68; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_68;
  reg [7:0] _T__69; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_69;
  reg [7:0] _T__70; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_70;
  reg [7:0] _T__71; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_71;
  reg [7:0] _T__72; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_72;
  reg [7:0] _T__73; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_73;
  reg [7:0] _T__74; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_74;
  reg [7:0] _T__75; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_75;
  reg [7:0] _T__76; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_76;
  reg [7:0] _T__77; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_77;
  reg [7:0] _T__78; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_78;
  reg [7:0] _T__79; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_79;
  reg [7:0] _T__80; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_80;
  reg [7:0] _T__81; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_81;
  reg [7:0] _T__82; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_82;
  reg [7:0] _T__83; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_83;
  reg [7:0] _T__84; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_84;
  reg [7:0] _T__85; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_85;
  reg [7:0] _T__86; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_86;
  reg [7:0] _T__87; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_87;
  reg [7:0] _T__88; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_88;
  reg [7:0] _T__89; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_89;
  reg [7:0] _T__90; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_90;
  reg [7:0] _T__91; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_91;
  reg [7:0] _T__92; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_92;
  reg [7:0] _T__93; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_93;
  reg [7:0] _T__94; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_94;
  reg [7:0] _T__95; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_95;
  reg [7:0] _T__96; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_96;
  reg [7:0] _T__97; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_97;
  reg [7:0] _T__98; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_98;
  reg [7:0] _T__99; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_99;
  reg [7:0] _T__100; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_100;
  reg [7:0] _T__101; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_101;
  reg [7:0] _T__102; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_102;
  reg [7:0] _T__103; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_103;
  reg [7:0] _T__104; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_104;
  reg [7:0] _T__105; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_105;
  reg [7:0] _T__106; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_106;
  reg [7:0] _T__107; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_107;
  reg [7:0] _T__108; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_108;
  reg [7:0] _T__109; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_109;
  reg [7:0] _T__110; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_110;
  reg [7:0] _T__111; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_111;
  reg [7:0] _T__112; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_112;
  reg [7:0] _T__113; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_113;
  reg [7:0] _T__114; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_114;
  reg [7:0] _T__115; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_115;
  reg [7:0] _T__116; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_116;
  reg [7:0] _T__117; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_117;
  reg [7:0] _T__118; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_118;
  reg [7:0] _T__119; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_119;
  reg [7:0] _T__120; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_120;
  reg [7:0] _T__121; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_121;
  reg [7:0] _T__122; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_122;
  reg [7:0] _T__123; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_123;
  reg [7:0] _T__124; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_124;
  reg [7:0] _T__125; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_125;
  reg [7:0] _T__126; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_126;
  reg [7:0] _T__127; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_127;
  reg [7:0] _T__128; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_128;
  reg [7:0] _T__129; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_129;
  reg [7:0] _T__130; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_130;
  reg [7:0] _T__131; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_131;
  reg [7:0] _T__132; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_132;
  reg [7:0] _T__133; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_133;
  reg [7:0] _T__134; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_134;
  reg [7:0] _T__135; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_135;
  reg [7:0] _T__136; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_136;
  reg [7:0] _T__137; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_137;
  reg [7:0] _T__138; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_138;
  reg [7:0] _T__139; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_139;
  reg [7:0] _T__140; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_140;
  reg [7:0] _T__141; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_141;
  reg [7:0] _T__142; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_142;
  reg [7:0] _T__143; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_143;
  reg [7:0] _T__144; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_144;
  reg [7:0] _T__145; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_145;
  reg [7:0] _T__146; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_146;
  reg [7:0] _T__147; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_147;
  reg [7:0] _T__148; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_148;
  reg [7:0] _T__149; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_149;
  reg [7:0] _T__150; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_150;
  reg [7:0] _T__151; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_151;
  reg [7:0] _T__152; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_152;
  reg [7:0] _T__153; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_153;
  reg [7:0] _T__154; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_154;
  reg [7:0] _T__155; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_155;
  reg [7:0] _T__156; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_156;
  reg [7:0] _T__157; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_157;
  reg [7:0] _T__158; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_158;
  reg [7:0] _T__159; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_159;
  reg [7:0] _T__160; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_160;
  reg [7:0] _T__161; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_161;
  reg [7:0] _T__162; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_162;
  reg [7:0] _T__163; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_163;
  reg [7:0] _T__164; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_164;
  reg [7:0] _T__165; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_165;
  reg [7:0] _T__166; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_166;
  reg [7:0] _T__167; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_167;
  reg [7:0] _T__168; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_168;
  reg [7:0] _T__169; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_169;
  reg [7:0] _T__170; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_170;
  reg [7:0] _T__171; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_171;
  reg [7:0] _T__172; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_172;
  reg [7:0] _T__173; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_173;
  reg [7:0] _T__174; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_174;
  reg [7:0] _T__175; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_175;
  reg [7:0] _T__176; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_176;
  reg [7:0] _T__177; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_177;
  reg [7:0] _T__178; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_178;
  reg [7:0] _T__179; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_179;
  reg [7:0] _T__180; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_180;
  reg [7:0] _T__181; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_181;
  reg [7:0] _T__182; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_182;
  reg [7:0] _T__183; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_183;
  reg [7:0] _T__184; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_184;
  reg [7:0] _T__185; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_185;
  reg [7:0] _T__186; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_186;
  reg [7:0] _T__187; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_187;
  reg [7:0] _T__188; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_188;
  reg [7:0] _T__189; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_189;
  reg [7:0] _T__190; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_190;
  reg [7:0] _T__191; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_191;
  reg [7:0] _T__192; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_192;
  reg [7:0] _T__193; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_193;
  reg [7:0] _T__194; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_194;
  reg [7:0] _T__195; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_195;
  reg [7:0] _T__196; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_196;
  reg [7:0] _T__197; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_197;
  reg [7:0] _T__198; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_198;
  reg [7:0] _T__199; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_199;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_200;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O_0 = _T__0; // @[FIFO.scala 14:7]
  assign O_1 = _T__1; // @[FIFO.scala 14:7]
  assign O_2 = _T__2; // @[FIFO.scala 14:7]
  assign O_3 = _T__3; // @[FIFO.scala 14:7]
  assign O_4 = _T__4; // @[FIFO.scala 14:7]
  assign O_5 = _T__5; // @[FIFO.scala 14:7]
  assign O_6 = _T__6; // @[FIFO.scala 14:7]
  assign O_7 = _T__7; // @[FIFO.scala 14:7]
  assign O_8 = _T__8; // @[FIFO.scala 14:7]
  assign O_9 = _T__9; // @[FIFO.scala 14:7]
  assign O_10 = _T__10; // @[FIFO.scala 14:7]
  assign O_11 = _T__11; // @[FIFO.scala 14:7]
  assign O_12 = _T__12; // @[FIFO.scala 14:7]
  assign O_13 = _T__13; // @[FIFO.scala 14:7]
  assign O_14 = _T__14; // @[FIFO.scala 14:7]
  assign O_15 = _T__15; // @[FIFO.scala 14:7]
  assign O_16 = _T__16; // @[FIFO.scala 14:7]
  assign O_17 = _T__17; // @[FIFO.scala 14:7]
  assign O_18 = _T__18; // @[FIFO.scala 14:7]
  assign O_19 = _T__19; // @[FIFO.scala 14:7]
  assign O_20 = _T__20; // @[FIFO.scala 14:7]
  assign O_21 = _T__21; // @[FIFO.scala 14:7]
  assign O_22 = _T__22; // @[FIFO.scala 14:7]
  assign O_23 = _T__23; // @[FIFO.scala 14:7]
  assign O_24 = _T__24; // @[FIFO.scala 14:7]
  assign O_25 = _T__25; // @[FIFO.scala 14:7]
  assign O_26 = _T__26; // @[FIFO.scala 14:7]
  assign O_27 = _T__27; // @[FIFO.scala 14:7]
  assign O_28 = _T__28; // @[FIFO.scala 14:7]
  assign O_29 = _T__29; // @[FIFO.scala 14:7]
  assign O_30 = _T__30; // @[FIFO.scala 14:7]
  assign O_31 = _T__31; // @[FIFO.scala 14:7]
  assign O_32 = _T__32; // @[FIFO.scala 14:7]
  assign O_33 = _T__33; // @[FIFO.scala 14:7]
  assign O_34 = _T__34; // @[FIFO.scala 14:7]
  assign O_35 = _T__35; // @[FIFO.scala 14:7]
  assign O_36 = _T__36; // @[FIFO.scala 14:7]
  assign O_37 = _T__37; // @[FIFO.scala 14:7]
  assign O_38 = _T__38; // @[FIFO.scala 14:7]
  assign O_39 = _T__39; // @[FIFO.scala 14:7]
  assign O_40 = _T__40; // @[FIFO.scala 14:7]
  assign O_41 = _T__41; // @[FIFO.scala 14:7]
  assign O_42 = _T__42; // @[FIFO.scala 14:7]
  assign O_43 = _T__43; // @[FIFO.scala 14:7]
  assign O_44 = _T__44; // @[FIFO.scala 14:7]
  assign O_45 = _T__45; // @[FIFO.scala 14:7]
  assign O_46 = _T__46; // @[FIFO.scala 14:7]
  assign O_47 = _T__47; // @[FIFO.scala 14:7]
  assign O_48 = _T__48; // @[FIFO.scala 14:7]
  assign O_49 = _T__49; // @[FIFO.scala 14:7]
  assign O_50 = _T__50; // @[FIFO.scala 14:7]
  assign O_51 = _T__51; // @[FIFO.scala 14:7]
  assign O_52 = _T__52; // @[FIFO.scala 14:7]
  assign O_53 = _T__53; // @[FIFO.scala 14:7]
  assign O_54 = _T__54; // @[FIFO.scala 14:7]
  assign O_55 = _T__55; // @[FIFO.scala 14:7]
  assign O_56 = _T__56; // @[FIFO.scala 14:7]
  assign O_57 = _T__57; // @[FIFO.scala 14:7]
  assign O_58 = _T__58; // @[FIFO.scala 14:7]
  assign O_59 = _T__59; // @[FIFO.scala 14:7]
  assign O_60 = _T__60; // @[FIFO.scala 14:7]
  assign O_61 = _T__61; // @[FIFO.scala 14:7]
  assign O_62 = _T__62; // @[FIFO.scala 14:7]
  assign O_63 = _T__63; // @[FIFO.scala 14:7]
  assign O_64 = _T__64; // @[FIFO.scala 14:7]
  assign O_65 = _T__65; // @[FIFO.scala 14:7]
  assign O_66 = _T__66; // @[FIFO.scala 14:7]
  assign O_67 = _T__67; // @[FIFO.scala 14:7]
  assign O_68 = _T__68; // @[FIFO.scala 14:7]
  assign O_69 = _T__69; // @[FIFO.scala 14:7]
  assign O_70 = _T__70; // @[FIFO.scala 14:7]
  assign O_71 = _T__71; // @[FIFO.scala 14:7]
  assign O_72 = _T__72; // @[FIFO.scala 14:7]
  assign O_73 = _T__73; // @[FIFO.scala 14:7]
  assign O_74 = _T__74; // @[FIFO.scala 14:7]
  assign O_75 = _T__75; // @[FIFO.scala 14:7]
  assign O_76 = _T__76; // @[FIFO.scala 14:7]
  assign O_77 = _T__77; // @[FIFO.scala 14:7]
  assign O_78 = _T__78; // @[FIFO.scala 14:7]
  assign O_79 = _T__79; // @[FIFO.scala 14:7]
  assign O_80 = _T__80; // @[FIFO.scala 14:7]
  assign O_81 = _T__81; // @[FIFO.scala 14:7]
  assign O_82 = _T__82; // @[FIFO.scala 14:7]
  assign O_83 = _T__83; // @[FIFO.scala 14:7]
  assign O_84 = _T__84; // @[FIFO.scala 14:7]
  assign O_85 = _T__85; // @[FIFO.scala 14:7]
  assign O_86 = _T__86; // @[FIFO.scala 14:7]
  assign O_87 = _T__87; // @[FIFO.scala 14:7]
  assign O_88 = _T__88; // @[FIFO.scala 14:7]
  assign O_89 = _T__89; // @[FIFO.scala 14:7]
  assign O_90 = _T__90; // @[FIFO.scala 14:7]
  assign O_91 = _T__91; // @[FIFO.scala 14:7]
  assign O_92 = _T__92; // @[FIFO.scala 14:7]
  assign O_93 = _T__93; // @[FIFO.scala 14:7]
  assign O_94 = _T__94; // @[FIFO.scala 14:7]
  assign O_95 = _T__95; // @[FIFO.scala 14:7]
  assign O_96 = _T__96; // @[FIFO.scala 14:7]
  assign O_97 = _T__97; // @[FIFO.scala 14:7]
  assign O_98 = _T__98; // @[FIFO.scala 14:7]
  assign O_99 = _T__99; // @[FIFO.scala 14:7]
  assign O_100 = _T__100; // @[FIFO.scala 14:7]
  assign O_101 = _T__101; // @[FIFO.scala 14:7]
  assign O_102 = _T__102; // @[FIFO.scala 14:7]
  assign O_103 = _T__103; // @[FIFO.scala 14:7]
  assign O_104 = _T__104; // @[FIFO.scala 14:7]
  assign O_105 = _T__105; // @[FIFO.scala 14:7]
  assign O_106 = _T__106; // @[FIFO.scala 14:7]
  assign O_107 = _T__107; // @[FIFO.scala 14:7]
  assign O_108 = _T__108; // @[FIFO.scala 14:7]
  assign O_109 = _T__109; // @[FIFO.scala 14:7]
  assign O_110 = _T__110; // @[FIFO.scala 14:7]
  assign O_111 = _T__111; // @[FIFO.scala 14:7]
  assign O_112 = _T__112; // @[FIFO.scala 14:7]
  assign O_113 = _T__113; // @[FIFO.scala 14:7]
  assign O_114 = _T__114; // @[FIFO.scala 14:7]
  assign O_115 = _T__115; // @[FIFO.scala 14:7]
  assign O_116 = _T__116; // @[FIFO.scala 14:7]
  assign O_117 = _T__117; // @[FIFO.scala 14:7]
  assign O_118 = _T__118; // @[FIFO.scala 14:7]
  assign O_119 = _T__119; // @[FIFO.scala 14:7]
  assign O_120 = _T__120; // @[FIFO.scala 14:7]
  assign O_121 = _T__121; // @[FIFO.scala 14:7]
  assign O_122 = _T__122; // @[FIFO.scala 14:7]
  assign O_123 = _T__123; // @[FIFO.scala 14:7]
  assign O_124 = _T__124; // @[FIFO.scala 14:7]
  assign O_125 = _T__125; // @[FIFO.scala 14:7]
  assign O_126 = _T__126; // @[FIFO.scala 14:7]
  assign O_127 = _T__127; // @[FIFO.scala 14:7]
  assign O_128 = _T__128; // @[FIFO.scala 14:7]
  assign O_129 = _T__129; // @[FIFO.scala 14:7]
  assign O_130 = _T__130; // @[FIFO.scala 14:7]
  assign O_131 = _T__131; // @[FIFO.scala 14:7]
  assign O_132 = _T__132; // @[FIFO.scala 14:7]
  assign O_133 = _T__133; // @[FIFO.scala 14:7]
  assign O_134 = _T__134; // @[FIFO.scala 14:7]
  assign O_135 = _T__135; // @[FIFO.scala 14:7]
  assign O_136 = _T__136; // @[FIFO.scala 14:7]
  assign O_137 = _T__137; // @[FIFO.scala 14:7]
  assign O_138 = _T__138; // @[FIFO.scala 14:7]
  assign O_139 = _T__139; // @[FIFO.scala 14:7]
  assign O_140 = _T__140; // @[FIFO.scala 14:7]
  assign O_141 = _T__141; // @[FIFO.scala 14:7]
  assign O_142 = _T__142; // @[FIFO.scala 14:7]
  assign O_143 = _T__143; // @[FIFO.scala 14:7]
  assign O_144 = _T__144; // @[FIFO.scala 14:7]
  assign O_145 = _T__145; // @[FIFO.scala 14:7]
  assign O_146 = _T__146; // @[FIFO.scala 14:7]
  assign O_147 = _T__147; // @[FIFO.scala 14:7]
  assign O_148 = _T__148; // @[FIFO.scala 14:7]
  assign O_149 = _T__149; // @[FIFO.scala 14:7]
  assign O_150 = _T__150; // @[FIFO.scala 14:7]
  assign O_151 = _T__151; // @[FIFO.scala 14:7]
  assign O_152 = _T__152; // @[FIFO.scala 14:7]
  assign O_153 = _T__153; // @[FIFO.scala 14:7]
  assign O_154 = _T__154; // @[FIFO.scala 14:7]
  assign O_155 = _T__155; // @[FIFO.scala 14:7]
  assign O_156 = _T__156; // @[FIFO.scala 14:7]
  assign O_157 = _T__157; // @[FIFO.scala 14:7]
  assign O_158 = _T__158; // @[FIFO.scala 14:7]
  assign O_159 = _T__159; // @[FIFO.scala 14:7]
  assign O_160 = _T__160; // @[FIFO.scala 14:7]
  assign O_161 = _T__161; // @[FIFO.scala 14:7]
  assign O_162 = _T__162; // @[FIFO.scala 14:7]
  assign O_163 = _T__163; // @[FIFO.scala 14:7]
  assign O_164 = _T__164; // @[FIFO.scala 14:7]
  assign O_165 = _T__165; // @[FIFO.scala 14:7]
  assign O_166 = _T__166; // @[FIFO.scala 14:7]
  assign O_167 = _T__167; // @[FIFO.scala 14:7]
  assign O_168 = _T__168; // @[FIFO.scala 14:7]
  assign O_169 = _T__169; // @[FIFO.scala 14:7]
  assign O_170 = _T__170; // @[FIFO.scala 14:7]
  assign O_171 = _T__171; // @[FIFO.scala 14:7]
  assign O_172 = _T__172; // @[FIFO.scala 14:7]
  assign O_173 = _T__173; // @[FIFO.scala 14:7]
  assign O_174 = _T__174; // @[FIFO.scala 14:7]
  assign O_175 = _T__175; // @[FIFO.scala 14:7]
  assign O_176 = _T__176; // @[FIFO.scala 14:7]
  assign O_177 = _T__177; // @[FIFO.scala 14:7]
  assign O_178 = _T__178; // @[FIFO.scala 14:7]
  assign O_179 = _T__179; // @[FIFO.scala 14:7]
  assign O_180 = _T__180; // @[FIFO.scala 14:7]
  assign O_181 = _T__181; // @[FIFO.scala 14:7]
  assign O_182 = _T__182; // @[FIFO.scala 14:7]
  assign O_183 = _T__183; // @[FIFO.scala 14:7]
  assign O_184 = _T__184; // @[FIFO.scala 14:7]
  assign O_185 = _T__185; // @[FIFO.scala 14:7]
  assign O_186 = _T__186; // @[FIFO.scala 14:7]
  assign O_187 = _T__187; // @[FIFO.scala 14:7]
  assign O_188 = _T__188; // @[FIFO.scala 14:7]
  assign O_189 = _T__189; // @[FIFO.scala 14:7]
  assign O_190 = _T__190; // @[FIFO.scala 14:7]
  assign O_191 = _T__191; // @[FIFO.scala 14:7]
  assign O_192 = _T__192; // @[FIFO.scala 14:7]
  assign O_193 = _T__193; // @[FIFO.scala 14:7]
  assign O_194 = _T__194; // @[FIFO.scala 14:7]
  assign O_195 = _T__195; // @[FIFO.scala 14:7]
  assign O_196 = _T__196; // @[FIFO.scala 14:7]
  assign O_197 = _T__197; // @[FIFO.scala 14:7]
  assign O_198 = _T__198; // @[FIFO.scala 14:7]
  assign O_199 = _T__199; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T__0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T__1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__3 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T__4 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T__5 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__6 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__7 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T__8 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T__9 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T__10 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T__11 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T__12 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T__13 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T__14 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T__15 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T__16 = _RAND_16[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T__17 = _RAND_17[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T__18 = _RAND_18[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T__19 = _RAND_19[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T__20 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T__21 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T__22 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T__23 = _RAND_23[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T__24 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T__25 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T__26 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T__27 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T__28 = _RAND_28[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T__29 = _RAND_29[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T__30 = _RAND_30[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T__31 = _RAND_31[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T__32 = _RAND_32[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T__33 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T__34 = _RAND_34[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T__35 = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T__36 = _RAND_36[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T__37 = _RAND_37[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T__38 = _RAND_38[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T__39 = _RAND_39[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T__40 = _RAND_40[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T__41 = _RAND_41[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T__42 = _RAND_42[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T__43 = _RAND_43[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T__44 = _RAND_44[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T__45 = _RAND_45[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T__46 = _RAND_46[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T__47 = _RAND_47[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T__48 = _RAND_48[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T__49 = _RAND_49[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T__50 = _RAND_50[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T__51 = _RAND_51[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T__52 = _RAND_52[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T__53 = _RAND_53[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T__54 = _RAND_54[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T__55 = _RAND_55[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T__56 = _RAND_56[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T__57 = _RAND_57[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T__58 = _RAND_58[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T__59 = _RAND_59[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T__60 = _RAND_60[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T__61 = _RAND_61[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T__62 = _RAND_62[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T__63 = _RAND_63[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T__64 = _RAND_64[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T__65 = _RAND_65[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T__66 = _RAND_66[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T__67 = _RAND_67[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T__68 = _RAND_68[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T__69 = _RAND_69[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T__70 = _RAND_70[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T__71 = _RAND_71[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T__72 = _RAND_72[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T__73 = _RAND_73[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T__74 = _RAND_74[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T__75 = _RAND_75[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T__76 = _RAND_76[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T__77 = _RAND_77[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T__78 = _RAND_78[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T__79 = _RAND_79[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T__80 = _RAND_80[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T__81 = _RAND_81[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T__82 = _RAND_82[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T__83 = _RAND_83[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T__84 = _RAND_84[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T__85 = _RAND_85[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T__86 = _RAND_86[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T__87 = _RAND_87[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T__88 = _RAND_88[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T__89 = _RAND_89[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T__90 = _RAND_90[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T__91 = _RAND_91[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T__92 = _RAND_92[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T__93 = _RAND_93[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T__94 = _RAND_94[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T__95 = _RAND_95[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T__96 = _RAND_96[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T__97 = _RAND_97[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T__98 = _RAND_98[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T__99 = _RAND_99[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T__100 = _RAND_100[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T__101 = _RAND_101[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T__102 = _RAND_102[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T__103 = _RAND_103[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T__104 = _RAND_104[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T__105 = _RAND_105[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T__106 = _RAND_106[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T__107 = _RAND_107[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T__108 = _RAND_108[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T__109 = _RAND_109[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T__110 = _RAND_110[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T__111 = _RAND_111[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T__112 = _RAND_112[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T__113 = _RAND_113[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T__114 = _RAND_114[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T__115 = _RAND_115[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T__116 = _RAND_116[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T__117 = _RAND_117[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T__118 = _RAND_118[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T__119 = _RAND_119[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T__120 = _RAND_120[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T__121 = _RAND_121[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T__122 = _RAND_122[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T__123 = _RAND_123[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T__124 = _RAND_124[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T__125 = _RAND_125[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T__126 = _RAND_126[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T__127 = _RAND_127[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T__128 = _RAND_128[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T__129 = _RAND_129[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T__130 = _RAND_130[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T__131 = _RAND_131[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T__132 = _RAND_132[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T__133 = _RAND_133[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T__134 = _RAND_134[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T__135 = _RAND_135[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T__136 = _RAND_136[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T__137 = _RAND_137[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T__138 = _RAND_138[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T__139 = _RAND_139[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T__140 = _RAND_140[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T__141 = _RAND_141[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T__142 = _RAND_142[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T__143 = _RAND_143[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T__144 = _RAND_144[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T__145 = _RAND_145[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T__146 = _RAND_146[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T__147 = _RAND_147[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T__148 = _RAND_148[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T__149 = _RAND_149[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T__150 = _RAND_150[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T__151 = _RAND_151[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T__152 = _RAND_152[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T__153 = _RAND_153[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T__154 = _RAND_154[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T__155 = _RAND_155[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T__156 = _RAND_156[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T__157 = _RAND_157[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T__158 = _RAND_158[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T__159 = _RAND_159[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T__160 = _RAND_160[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T__161 = _RAND_161[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T__162 = _RAND_162[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T__163 = _RAND_163[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T__164 = _RAND_164[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T__165 = _RAND_165[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T__166 = _RAND_166[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T__167 = _RAND_167[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T__168 = _RAND_168[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T__169 = _RAND_169[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T__170 = _RAND_170[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T__171 = _RAND_171[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T__172 = _RAND_172[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T__173 = _RAND_173[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T__174 = _RAND_174[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T__175 = _RAND_175[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T__176 = _RAND_176[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T__177 = _RAND_177[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T__178 = _RAND_178[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T__179 = _RAND_179[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T__180 = _RAND_180[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T__181 = _RAND_181[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T__182 = _RAND_182[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T__183 = _RAND_183[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T__184 = _RAND_184[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T__185 = _RAND_185[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T__186 = _RAND_186[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T__187 = _RAND_187[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T__188 = _RAND_188[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T__189 = _RAND_189[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T__190 = _RAND_190[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T__191 = _RAND_191[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T__192 = _RAND_192[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T__193 = _RAND_193[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T__194 = _RAND_194[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T__195 = _RAND_195[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T__196 = _RAND_196[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T__197 = _RAND_197[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T__198 = _RAND_198[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T__199 = _RAND_199[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_1 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T__0 <= I_0;
    _T__1 <= I_1;
    _T__2 <= I_2;
    _T__3 <= I_3;
    _T__4 <= I_4;
    _T__5 <= I_5;
    _T__6 <= I_6;
    _T__7 <= I_7;
    _T__8 <= I_8;
    _T__9 <= I_9;
    _T__10 <= I_10;
    _T__11 <= I_11;
    _T__12 <= I_12;
    _T__13 <= I_13;
    _T__14 <= I_14;
    _T__15 <= I_15;
    _T__16 <= I_16;
    _T__17 <= I_17;
    _T__18 <= I_18;
    _T__19 <= I_19;
    _T__20 <= I_20;
    _T__21 <= I_21;
    _T__22 <= I_22;
    _T__23 <= I_23;
    _T__24 <= I_24;
    _T__25 <= I_25;
    _T__26 <= I_26;
    _T__27 <= I_27;
    _T__28 <= I_28;
    _T__29 <= I_29;
    _T__30 <= I_30;
    _T__31 <= I_31;
    _T__32 <= I_32;
    _T__33 <= I_33;
    _T__34 <= I_34;
    _T__35 <= I_35;
    _T__36 <= I_36;
    _T__37 <= I_37;
    _T__38 <= I_38;
    _T__39 <= I_39;
    _T__40 <= I_40;
    _T__41 <= I_41;
    _T__42 <= I_42;
    _T__43 <= I_43;
    _T__44 <= I_44;
    _T__45 <= I_45;
    _T__46 <= I_46;
    _T__47 <= I_47;
    _T__48 <= I_48;
    _T__49 <= I_49;
    _T__50 <= I_50;
    _T__51 <= I_51;
    _T__52 <= I_52;
    _T__53 <= I_53;
    _T__54 <= I_54;
    _T__55 <= I_55;
    _T__56 <= I_56;
    _T__57 <= I_57;
    _T__58 <= I_58;
    _T__59 <= I_59;
    _T__60 <= I_60;
    _T__61 <= I_61;
    _T__62 <= I_62;
    _T__63 <= I_63;
    _T__64 <= I_64;
    _T__65 <= I_65;
    _T__66 <= I_66;
    _T__67 <= I_67;
    _T__68 <= I_68;
    _T__69 <= I_69;
    _T__70 <= I_70;
    _T__71 <= I_71;
    _T__72 <= I_72;
    _T__73 <= I_73;
    _T__74 <= I_74;
    _T__75 <= I_75;
    _T__76 <= I_76;
    _T__77 <= I_77;
    _T__78 <= I_78;
    _T__79 <= I_79;
    _T__80 <= I_80;
    _T__81 <= I_81;
    _T__82 <= I_82;
    _T__83 <= I_83;
    _T__84 <= I_84;
    _T__85 <= I_85;
    _T__86 <= I_86;
    _T__87 <= I_87;
    _T__88 <= I_88;
    _T__89 <= I_89;
    _T__90 <= I_90;
    _T__91 <= I_91;
    _T__92 <= I_92;
    _T__93 <= I_93;
    _T__94 <= I_94;
    _T__95 <= I_95;
    _T__96 <= I_96;
    _T__97 <= I_97;
    _T__98 <= I_98;
    _T__99 <= I_99;
    _T__100 <= I_100;
    _T__101 <= I_101;
    _T__102 <= I_102;
    _T__103 <= I_103;
    _T__104 <= I_104;
    _T__105 <= I_105;
    _T__106 <= I_106;
    _T__107 <= I_107;
    _T__108 <= I_108;
    _T__109 <= I_109;
    _T__110 <= I_110;
    _T__111 <= I_111;
    _T__112 <= I_112;
    _T__113 <= I_113;
    _T__114 <= I_114;
    _T__115 <= I_115;
    _T__116 <= I_116;
    _T__117 <= I_117;
    _T__118 <= I_118;
    _T__119 <= I_119;
    _T__120 <= I_120;
    _T__121 <= I_121;
    _T__122 <= I_122;
    _T__123 <= I_123;
    _T__124 <= I_124;
    _T__125 <= I_125;
    _T__126 <= I_126;
    _T__127 <= I_127;
    _T__128 <= I_128;
    _T__129 <= I_129;
    _T__130 <= I_130;
    _T__131 <= I_131;
    _T__132 <= I_132;
    _T__133 <= I_133;
    _T__134 <= I_134;
    _T__135 <= I_135;
    _T__136 <= I_136;
    _T__137 <= I_137;
    _T__138 <= I_138;
    _T__139 <= I_139;
    _T__140 <= I_140;
    _T__141 <= I_141;
    _T__142 <= I_142;
    _T__143 <= I_143;
    _T__144 <= I_144;
    _T__145 <= I_145;
    _T__146 <= I_146;
    _T__147 <= I_147;
    _T__148 <= I_148;
    _T__149 <= I_149;
    _T__150 <= I_150;
    _T__151 <= I_151;
    _T__152 <= I_152;
    _T__153 <= I_153;
    _T__154 <= I_154;
    _T__155 <= I_155;
    _T__156 <= I_156;
    _T__157 <= I_157;
    _T__158 <= I_158;
    _T__159 <= I_159;
    _T__160 <= I_160;
    _T__161 <= I_161;
    _T__162 <= I_162;
    _T__163 <= I_163;
    _T__164 <= I_164;
    _T__165 <= I_165;
    _T__166 <= I_166;
    _T__167 <= I_167;
    _T__168 <= I_168;
    _T__169 <= I_169;
    _T__170 <= I_170;
    _T__171 <= I_171;
    _T__172 <= I_172;
    _T__173 <= I_173;
    _T__174 <= I_174;
    _T__175 <= I_175;
    _T__176 <= I_176;
    _T__177 <= I_177;
    _T__178 <= I_178;
    _T__179 <= I_179;
    _T__180 <= I_180;
    _T__181 <= I_181;
    _T__182 <= I_182;
    _T__183 <= I_183;
    _T__184 <= I_184;
    _T__185 <= I_185;
    _T__186 <= I_186;
    _T__187 <= I_187;
    _T__188 <= I_188;
    _T__189 <= I_189;
    _T__190 <= I_190;
    _T__191 <= I_191;
    _T__192 <= I_192;
    _T__193 <= I_193;
    _T__194 <= I_194;
    _T__195 <= I_195;
    _T__196 <= I_196;
    _T__197 <= I_197;
    _T__198 <= I_198;
    _T__199 <= I_199;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module InitialDelayCounter(
  input   clock,
  input   reset,
  output  valid_down
);
  reg  value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire  _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 1'h1; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 1'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 1'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module AtomTuple(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  output [7:0] O_t0b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
endmodule
module Add(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  output [7:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 108:14]
  assign O = I_t0b + 8'h5; // @[Arithmetic.scala 106:7]
endmodule
module Module_0(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I,
  output [7:0] O
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n5_valid_up; // @[Top.scala 18:20]
  wire  n5_valid_down; // @[Top.scala 18:20]
  wire [7:0] n5_I0; // @[Top.scala 18:20]
  wire [7:0] n5_O_t0b; // @[Top.scala 18:20]
  wire  n6_valid_up; // @[Top.scala 22:20]
  wire  n6_valid_down; // @[Top.scala 22:20]
  wire [7:0] n6_I_t0b; // @[Top.scala 22:20]
  wire [7:0] n6_O; // @[Top.scala 22:20]
  InitialDelayCounter InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  AtomTuple n5 ( // @[Top.scala 18:20]
    .valid_up(n5_valid_up),
    .valid_down(n5_valid_down),
    .I0(n5_I0),
    .O_t0b(n5_O_t0b)
  );
  Add n6 ( // @[Top.scala 22:20]
    .valid_up(n6_valid_up),
    .valid_down(n6_valid_down),
    .I_t0b(n6_I_t0b),
    .O(n6_O)
  );
  assign valid_down = n6_valid_down; // @[Top.scala 26:16]
  assign O = n6_O; // @[Top.scala 25:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n5_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 21:17]
  assign n5_I0 = I; // @[Top.scala 19:11]
  assign n6_valid_up = n5_valid_down; // @[Top.scala 24:17]
  assign n6_I_t0b = n5_O_t0b; // @[Top.scala 23:10]
endmodule
module MapS(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  input  [7:0] I_4,
  input  [7:0] I_5,
  input  [7:0] I_6,
  input  [7:0] I_7,
  input  [7:0] I_8,
  input  [7:0] I_9,
  input  [7:0] I_10,
  input  [7:0] I_11,
  input  [7:0] I_12,
  input  [7:0] I_13,
  input  [7:0] I_14,
  input  [7:0] I_15,
  input  [7:0] I_16,
  input  [7:0] I_17,
  input  [7:0] I_18,
  input  [7:0] I_19,
  input  [7:0] I_20,
  input  [7:0] I_21,
  input  [7:0] I_22,
  input  [7:0] I_23,
  input  [7:0] I_24,
  input  [7:0] I_25,
  input  [7:0] I_26,
  input  [7:0] I_27,
  input  [7:0] I_28,
  input  [7:0] I_29,
  input  [7:0] I_30,
  input  [7:0] I_31,
  input  [7:0] I_32,
  input  [7:0] I_33,
  input  [7:0] I_34,
  input  [7:0] I_35,
  input  [7:0] I_36,
  input  [7:0] I_37,
  input  [7:0] I_38,
  input  [7:0] I_39,
  input  [7:0] I_40,
  input  [7:0] I_41,
  input  [7:0] I_42,
  input  [7:0] I_43,
  input  [7:0] I_44,
  input  [7:0] I_45,
  input  [7:0] I_46,
  input  [7:0] I_47,
  input  [7:0] I_48,
  input  [7:0] I_49,
  input  [7:0] I_50,
  input  [7:0] I_51,
  input  [7:0] I_52,
  input  [7:0] I_53,
  input  [7:0] I_54,
  input  [7:0] I_55,
  input  [7:0] I_56,
  input  [7:0] I_57,
  input  [7:0] I_58,
  input  [7:0] I_59,
  input  [7:0] I_60,
  input  [7:0] I_61,
  input  [7:0] I_62,
  input  [7:0] I_63,
  input  [7:0] I_64,
  input  [7:0] I_65,
  input  [7:0] I_66,
  input  [7:0] I_67,
  input  [7:0] I_68,
  input  [7:0] I_69,
  input  [7:0] I_70,
  input  [7:0] I_71,
  input  [7:0] I_72,
  input  [7:0] I_73,
  input  [7:0] I_74,
  input  [7:0] I_75,
  input  [7:0] I_76,
  input  [7:0] I_77,
  input  [7:0] I_78,
  input  [7:0] I_79,
  input  [7:0] I_80,
  input  [7:0] I_81,
  input  [7:0] I_82,
  input  [7:0] I_83,
  input  [7:0] I_84,
  input  [7:0] I_85,
  input  [7:0] I_86,
  input  [7:0] I_87,
  input  [7:0] I_88,
  input  [7:0] I_89,
  input  [7:0] I_90,
  input  [7:0] I_91,
  input  [7:0] I_92,
  input  [7:0] I_93,
  input  [7:0] I_94,
  input  [7:0] I_95,
  input  [7:0] I_96,
  input  [7:0] I_97,
  input  [7:0] I_98,
  input  [7:0] I_99,
  input  [7:0] I_100,
  input  [7:0] I_101,
  input  [7:0] I_102,
  input  [7:0] I_103,
  input  [7:0] I_104,
  input  [7:0] I_105,
  input  [7:0] I_106,
  input  [7:0] I_107,
  input  [7:0] I_108,
  input  [7:0] I_109,
  input  [7:0] I_110,
  input  [7:0] I_111,
  input  [7:0] I_112,
  input  [7:0] I_113,
  input  [7:0] I_114,
  input  [7:0] I_115,
  input  [7:0] I_116,
  input  [7:0] I_117,
  input  [7:0] I_118,
  input  [7:0] I_119,
  input  [7:0] I_120,
  input  [7:0] I_121,
  input  [7:0] I_122,
  input  [7:0] I_123,
  input  [7:0] I_124,
  input  [7:0] I_125,
  input  [7:0] I_126,
  input  [7:0] I_127,
  input  [7:0] I_128,
  input  [7:0] I_129,
  input  [7:0] I_130,
  input  [7:0] I_131,
  input  [7:0] I_132,
  input  [7:0] I_133,
  input  [7:0] I_134,
  input  [7:0] I_135,
  input  [7:0] I_136,
  input  [7:0] I_137,
  input  [7:0] I_138,
  input  [7:0] I_139,
  input  [7:0] I_140,
  input  [7:0] I_141,
  input  [7:0] I_142,
  input  [7:0] I_143,
  input  [7:0] I_144,
  input  [7:0] I_145,
  input  [7:0] I_146,
  input  [7:0] I_147,
  input  [7:0] I_148,
  input  [7:0] I_149,
  input  [7:0] I_150,
  input  [7:0] I_151,
  input  [7:0] I_152,
  input  [7:0] I_153,
  input  [7:0] I_154,
  input  [7:0] I_155,
  input  [7:0] I_156,
  input  [7:0] I_157,
  input  [7:0] I_158,
  input  [7:0] I_159,
  input  [7:0] I_160,
  input  [7:0] I_161,
  input  [7:0] I_162,
  input  [7:0] I_163,
  input  [7:0] I_164,
  input  [7:0] I_165,
  input  [7:0] I_166,
  input  [7:0] I_167,
  input  [7:0] I_168,
  input  [7:0] I_169,
  input  [7:0] I_170,
  input  [7:0] I_171,
  input  [7:0] I_172,
  input  [7:0] I_173,
  input  [7:0] I_174,
  input  [7:0] I_175,
  input  [7:0] I_176,
  input  [7:0] I_177,
  input  [7:0] I_178,
  input  [7:0] I_179,
  input  [7:0] I_180,
  input  [7:0] I_181,
  input  [7:0] I_182,
  input  [7:0] I_183,
  input  [7:0] I_184,
  input  [7:0] I_185,
  input  [7:0] I_186,
  input  [7:0] I_187,
  input  [7:0] I_188,
  input  [7:0] I_189,
  input  [7:0] I_190,
  input  [7:0] I_191,
  input  [7:0] I_192,
  input  [7:0] I_193,
  input  [7:0] I_194,
  input  [7:0] I_195,
  input  [7:0] I_196,
  input  [7:0] I_197,
  input  [7:0] I_198,
  input  [7:0] I_199,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15,
  output [7:0] O_16,
  output [7:0] O_17,
  output [7:0] O_18,
  output [7:0] O_19,
  output [7:0] O_20,
  output [7:0] O_21,
  output [7:0] O_22,
  output [7:0] O_23,
  output [7:0] O_24,
  output [7:0] O_25,
  output [7:0] O_26,
  output [7:0] O_27,
  output [7:0] O_28,
  output [7:0] O_29,
  output [7:0] O_30,
  output [7:0] O_31,
  output [7:0] O_32,
  output [7:0] O_33,
  output [7:0] O_34,
  output [7:0] O_35,
  output [7:0] O_36,
  output [7:0] O_37,
  output [7:0] O_38,
  output [7:0] O_39,
  output [7:0] O_40,
  output [7:0] O_41,
  output [7:0] O_42,
  output [7:0] O_43,
  output [7:0] O_44,
  output [7:0] O_45,
  output [7:0] O_46,
  output [7:0] O_47,
  output [7:0] O_48,
  output [7:0] O_49,
  output [7:0] O_50,
  output [7:0] O_51,
  output [7:0] O_52,
  output [7:0] O_53,
  output [7:0] O_54,
  output [7:0] O_55,
  output [7:0] O_56,
  output [7:0] O_57,
  output [7:0] O_58,
  output [7:0] O_59,
  output [7:0] O_60,
  output [7:0] O_61,
  output [7:0] O_62,
  output [7:0] O_63,
  output [7:0] O_64,
  output [7:0] O_65,
  output [7:0] O_66,
  output [7:0] O_67,
  output [7:0] O_68,
  output [7:0] O_69,
  output [7:0] O_70,
  output [7:0] O_71,
  output [7:0] O_72,
  output [7:0] O_73,
  output [7:0] O_74,
  output [7:0] O_75,
  output [7:0] O_76,
  output [7:0] O_77,
  output [7:0] O_78,
  output [7:0] O_79,
  output [7:0] O_80,
  output [7:0] O_81,
  output [7:0] O_82,
  output [7:0] O_83,
  output [7:0] O_84,
  output [7:0] O_85,
  output [7:0] O_86,
  output [7:0] O_87,
  output [7:0] O_88,
  output [7:0] O_89,
  output [7:0] O_90,
  output [7:0] O_91,
  output [7:0] O_92,
  output [7:0] O_93,
  output [7:0] O_94,
  output [7:0] O_95,
  output [7:0] O_96,
  output [7:0] O_97,
  output [7:0] O_98,
  output [7:0] O_99,
  output [7:0] O_100,
  output [7:0] O_101,
  output [7:0] O_102,
  output [7:0] O_103,
  output [7:0] O_104,
  output [7:0] O_105,
  output [7:0] O_106,
  output [7:0] O_107,
  output [7:0] O_108,
  output [7:0] O_109,
  output [7:0] O_110,
  output [7:0] O_111,
  output [7:0] O_112,
  output [7:0] O_113,
  output [7:0] O_114,
  output [7:0] O_115,
  output [7:0] O_116,
  output [7:0] O_117,
  output [7:0] O_118,
  output [7:0] O_119,
  output [7:0] O_120,
  output [7:0] O_121,
  output [7:0] O_122,
  output [7:0] O_123,
  output [7:0] O_124,
  output [7:0] O_125,
  output [7:0] O_126,
  output [7:0] O_127,
  output [7:0] O_128,
  output [7:0] O_129,
  output [7:0] O_130,
  output [7:0] O_131,
  output [7:0] O_132,
  output [7:0] O_133,
  output [7:0] O_134,
  output [7:0] O_135,
  output [7:0] O_136,
  output [7:0] O_137,
  output [7:0] O_138,
  output [7:0] O_139,
  output [7:0] O_140,
  output [7:0] O_141,
  output [7:0] O_142,
  output [7:0] O_143,
  output [7:0] O_144,
  output [7:0] O_145,
  output [7:0] O_146,
  output [7:0] O_147,
  output [7:0] O_148,
  output [7:0] O_149,
  output [7:0] O_150,
  output [7:0] O_151,
  output [7:0] O_152,
  output [7:0] O_153,
  output [7:0] O_154,
  output [7:0] O_155,
  output [7:0] O_156,
  output [7:0] O_157,
  output [7:0] O_158,
  output [7:0] O_159,
  output [7:0] O_160,
  output [7:0] O_161,
  output [7:0] O_162,
  output [7:0] O_163,
  output [7:0] O_164,
  output [7:0] O_165,
  output [7:0] O_166,
  output [7:0] O_167,
  output [7:0] O_168,
  output [7:0] O_169,
  output [7:0] O_170,
  output [7:0] O_171,
  output [7:0] O_172,
  output [7:0] O_173,
  output [7:0] O_174,
  output [7:0] O_175,
  output [7:0] O_176,
  output [7:0] O_177,
  output [7:0] O_178,
  output [7:0] O_179,
  output [7:0] O_180,
  output [7:0] O_181,
  output [7:0] O_182,
  output [7:0] O_183,
  output [7:0] O_184,
  output [7:0] O_185,
  output [7:0] O_186,
  output [7:0] O_187,
  output [7:0] O_188,
  output [7:0] O_189,
  output [7:0] O_190,
  output [7:0] O_191,
  output [7:0] O_192,
  output [7:0] O_193,
  output [7:0] O_194,
  output [7:0] O_195,
  output [7:0] O_196,
  output [7:0] O_197,
  output [7:0] O_198,
  output [7:0] O_199
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O; // @[MapS.scala 10:86]
  wire  other_ops_2_clock; // @[MapS.scala 10:86]
  wire  other_ops_2_reset; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O; // @[MapS.scala 10:86]
  wire  other_ops_3_clock; // @[MapS.scala 10:86]
  wire  other_ops_3_reset; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O; // @[MapS.scala 10:86]
  wire  other_ops_4_clock; // @[MapS.scala 10:86]
  wire  other_ops_4_reset; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O; // @[MapS.scala 10:86]
  wire  other_ops_5_clock; // @[MapS.scala 10:86]
  wire  other_ops_5_reset; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O; // @[MapS.scala 10:86]
  wire  other_ops_6_clock; // @[MapS.scala 10:86]
  wire  other_ops_6_reset; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O; // @[MapS.scala 10:86]
  wire  other_ops_7_clock; // @[MapS.scala 10:86]
  wire  other_ops_7_reset; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O; // @[MapS.scala 10:86]
  wire  other_ops_8_clock; // @[MapS.scala 10:86]
  wire  other_ops_8_reset; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O; // @[MapS.scala 10:86]
  wire  other_ops_9_clock; // @[MapS.scala 10:86]
  wire  other_ops_9_reset; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O; // @[MapS.scala 10:86]
  wire  other_ops_10_clock; // @[MapS.scala 10:86]
  wire  other_ops_10_reset; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O; // @[MapS.scala 10:86]
  wire  other_ops_11_clock; // @[MapS.scala 10:86]
  wire  other_ops_11_reset; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O; // @[MapS.scala 10:86]
  wire  other_ops_12_clock; // @[MapS.scala 10:86]
  wire  other_ops_12_reset; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O; // @[MapS.scala 10:86]
  wire  other_ops_13_clock; // @[MapS.scala 10:86]
  wire  other_ops_13_reset; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O; // @[MapS.scala 10:86]
  wire  other_ops_14_clock; // @[MapS.scala 10:86]
  wire  other_ops_14_reset; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O; // @[MapS.scala 10:86]
  wire  other_ops_15_clock; // @[MapS.scala 10:86]
  wire  other_ops_15_reset; // @[MapS.scala 10:86]
  wire  other_ops_15_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_15_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_15_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_15_O; // @[MapS.scala 10:86]
  wire  other_ops_16_clock; // @[MapS.scala 10:86]
  wire  other_ops_16_reset; // @[MapS.scala 10:86]
  wire  other_ops_16_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_16_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_16_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_16_O; // @[MapS.scala 10:86]
  wire  other_ops_17_clock; // @[MapS.scala 10:86]
  wire  other_ops_17_reset; // @[MapS.scala 10:86]
  wire  other_ops_17_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_17_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_17_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_17_O; // @[MapS.scala 10:86]
  wire  other_ops_18_clock; // @[MapS.scala 10:86]
  wire  other_ops_18_reset; // @[MapS.scala 10:86]
  wire  other_ops_18_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_18_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_18_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_18_O; // @[MapS.scala 10:86]
  wire  other_ops_19_clock; // @[MapS.scala 10:86]
  wire  other_ops_19_reset; // @[MapS.scala 10:86]
  wire  other_ops_19_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_19_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_19_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_19_O; // @[MapS.scala 10:86]
  wire  other_ops_20_clock; // @[MapS.scala 10:86]
  wire  other_ops_20_reset; // @[MapS.scala 10:86]
  wire  other_ops_20_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_20_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_20_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_20_O; // @[MapS.scala 10:86]
  wire  other_ops_21_clock; // @[MapS.scala 10:86]
  wire  other_ops_21_reset; // @[MapS.scala 10:86]
  wire  other_ops_21_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_21_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_21_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_21_O; // @[MapS.scala 10:86]
  wire  other_ops_22_clock; // @[MapS.scala 10:86]
  wire  other_ops_22_reset; // @[MapS.scala 10:86]
  wire  other_ops_22_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_22_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_22_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_22_O; // @[MapS.scala 10:86]
  wire  other_ops_23_clock; // @[MapS.scala 10:86]
  wire  other_ops_23_reset; // @[MapS.scala 10:86]
  wire  other_ops_23_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_23_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_23_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_23_O; // @[MapS.scala 10:86]
  wire  other_ops_24_clock; // @[MapS.scala 10:86]
  wire  other_ops_24_reset; // @[MapS.scala 10:86]
  wire  other_ops_24_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_24_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_24_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_24_O; // @[MapS.scala 10:86]
  wire  other_ops_25_clock; // @[MapS.scala 10:86]
  wire  other_ops_25_reset; // @[MapS.scala 10:86]
  wire  other_ops_25_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_25_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_25_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_25_O; // @[MapS.scala 10:86]
  wire  other_ops_26_clock; // @[MapS.scala 10:86]
  wire  other_ops_26_reset; // @[MapS.scala 10:86]
  wire  other_ops_26_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_26_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_26_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_26_O; // @[MapS.scala 10:86]
  wire  other_ops_27_clock; // @[MapS.scala 10:86]
  wire  other_ops_27_reset; // @[MapS.scala 10:86]
  wire  other_ops_27_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_27_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_27_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_27_O; // @[MapS.scala 10:86]
  wire  other_ops_28_clock; // @[MapS.scala 10:86]
  wire  other_ops_28_reset; // @[MapS.scala 10:86]
  wire  other_ops_28_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_28_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_28_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_28_O; // @[MapS.scala 10:86]
  wire  other_ops_29_clock; // @[MapS.scala 10:86]
  wire  other_ops_29_reset; // @[MapS.scala 10:86]
  wire  other_ops_29_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_29_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_29_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_29_O; // @[MapS.scala 10:86]
  wire  other_ops_30_clock; // @[MapS.scala 10:86]
  wire  other_ops_30_reset; // @[MapS.scala 10:86]
  wire  other_ops_30_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_30_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_30_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_30_O; // @[MapS.scala 10:86]
  wire  other_ops_31_clock; // @[MapS.scala 10:86]
  wire  other_ops_31_reset; // @[MapS.scala 10:86]
  wire  other_ops_31_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_31_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_31_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_31_O; // @[MapS.scala 10:86]
  wire  other_ops_32_clock; // @[MapS.scala 10:86]
  wire  other_ops_32_reset; // @[MapS.scala 10:86]
  wire  other_ops_32_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_32_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_32_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_32_O; // @[MapS.scala 10:86]
  wire  other_ops_33_clock; // @[MapS.scala 10:86]
  wire  other_ops_33_reset; // @[MapS.scala 10:86]
  wire  other_ops_33_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_33_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_33_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_33_O; // @[MapS.scala 10:86]
  wire  other_ops_34_clock; // @[MapS.scala 10:86]
  wire  other_ops_34_reset; // @[MapS.scala 10:86]
  wire  other_ops_34_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_34_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_34_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_34_O; // @[MapS.scala 10:86]
  wire  other_ops_35_clock; // @[MapS.scala 10:86]
  wire  other_ops_35_reset; // @[MapS.scala 10:86]
  wire  other_ops_35_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_35_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_35_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_35_O; // @[MapS.scala 10:86]
  wire  other_ops_36_clock; // @[MapS.scala 10:86]
  wire  other_ops_36_reset; // @[MapS.scala 10:86]
  wire  other_ops_36_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_36_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_36_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_36_O; // @[MapS.scala 10:86]
  wire  other_ops_37_clock; // @[MapS.scala 10:86]
  wire  other_ops_37_reset; // @[MapS.scala 10:86]
  wire  other_ops_37_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_37_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_37_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_37_O; // @[MapS.scala 10:86]
  wire  other_ops_38_clock; // @[MapS.scala 10:86]
  wire  other_ops_38_reset; // @[MapS.scala 10:86]
  wire  other_ops_38_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_38_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_38_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_38_O; // @[MapS.scala 10:86]
  wire  other_ops_39_clock; // @[MapS.scala 10:86]
  wire  other_ops_39_reset; // @[MapS.scala 10:86]
  wire  other_ops_39_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_39_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_39_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_39_O; // @[MapS.scala 10:86]
  wire  other_ops_40_clock; // @[MapS.scala 10:86]
  wire  other_ops_40_reset; // @[MapS.scala 10:86]
  wire  other_ops_40_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_40_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_40_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_40_O; // @[MapS.scala 10:86]
  wire  other_ops_41_clock; // @[MapS.scala 10:86]
  wire  other_ops_41_reset; // @[MapS.scala 10:86]
  wire  other_ops_41_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_41_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_41_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_41_O; // @[MapS.scala 10:86]
  wire  other_ops_42_clock; // @[MapS.scala 10:86]
  wire  other_ops_42_reset; // @[MapS.scala 10:86]
  wire  other_ops_42_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_42_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_42_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_42_O; // @[MapS.scala 10:86]
  wire  other_ops_43_clock; // @[MapS.scala 10:86]
  wire  other_ops_43_reset; // @[MapS.scala 10:86]
  wire  other_ops_43_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_43_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_43_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_43_O; // @[MapS.scala 10:86]
  wire  other_ops_44_clock; // @[MapS.scala 10:86]
  wire  other_ops_44_reset; // @[MapS.scala 10:86]
  wire  other_ops_44_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_44_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_44_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_44_O; // @[MapS.scala 10:86]
  wire  other_ops_45_clock; // @[MapS.scala 10:86]
  wire  other_ops_45_reset; // @[MapS.scala 10:86]
  wire  other_ops_45_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_45_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_45_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_45_O; // @[MapS.scala 10:86]
  wire  other_ops_46_clock; // @[MapS.scala 10:86]
  wire  other_ops_46_reset; // @[MapS.scala 10:86]
  wire  other_ops_46_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_46_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_46_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_46_O; // @[MapS.scala 10:86]
  wire  other_ops_47_clock; // @[MapS.scala 10:86]
  wire  other_ops_47_reset; // @[MapS.scala 10:86]
  wire  other_ops_47_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_47_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_47_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_47_O; // @[MapS.scala 10:86]
  wire  other_ops_48_clock; // @[MapS.scala 10:86]
  wire  other_ops_48_reset; // @[MapS.scala 10:86]
  wire  other_ops_48_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_48_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_48_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_48_O; // @[MapS.scala 10:86]
  wire  other_ops_49_clock; // @[MapS.scala 10:86]
  wire  other_ops_49_reset; // @[MapS.scala 10:86]
  wire  other_ops_49_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_49_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_49_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_49_O; // @[MapS.scala 10:86]
  wire  other_ops_50_clock; // @[MapS.scala 10:86]
  wire  other_ops_50_reset; // @[MapS.scala 10:86]
  wire  other_ops_50_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_50_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_50_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_50_O; // @[MapS.scala 10:86]
  wire  other_ops_51_clock; // @[MapS.scala 10:86]
  wire  other_ops_51_reset; // @[MapS.scala 10:86]
  wire  other_ops_51_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_51_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_51_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_51_O; // @[MapS.scala 10:86]
  wire  other_ops_52_clock; // @[MapS.scala 10:86]
  wire  other_ops_52_reset; // @[MapS.scala 10:86]
  wire  other_ops_52_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_52_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_52_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_52_O; // @[MapS.scala 10:86]
  wire  other_ops_53_clock; // @[MapS.scala 10:86]
  wire  other_ops_53_reset; // @[MapS.scala 10:86]
  wire  other_ops_53_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_53_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_53_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_53_O; // @[MapS.scala 10:86]
  wire  other_ops_54_clock; // @[MapS.scala 10:86]
  wire  other_ops_54_reset; // @[MapS.scala 10:86]
  wire  other_ops_54_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_54_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_54_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_54_O; // @[MapS.scala 10:86]
  wire  other_ops_55_clock; // @[MapS.scala 10:86]
  wire  other_ops_55_reset; // @[MapS.scala 10:86]
  wire  other_ops_55_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_55_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_55_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_55_O; // @[MapS.scala 10:86]
  wire  other_ops_56_clock; // @[MapS.scala 10:86]
  wire  other_ops_56_reset; // @[MapS.scala 10:86]
  wire  other_ops_56_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_56_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_56_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_56_O; // @[MapS.scala 10:86]
  wire  other_ops_57_clock; // @[MapS.scala 10:86]
  wire  other_ops_57_reset; // @[MapS.scala 10:86]
  wire  other_ops_57_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_57_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_57_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_57_O; // @[MapS.scala 10:86]
  wire  other_ops_58_clock; // @[MapS.scala 10:86]
  wire  other_ops_58_reset; // @[MapS.scala 10:86]
  wire  other_ops_58_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_58_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_58_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_58_O; // @[MapS.scala 10:86]
  wire  other_ops_59_clock; // @[MapS.scala 10:86]
  wire  other_ops_59_reset; // @[MapS.scala 10:86]
  wire  other_ops_59_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_59_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_59_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_59_O; // @[MapS.scala 10:86]
  wire  other_ops_60_clock; // @[MapS.scala 10:86]
  wire  other_ops_60_reset; // @[MapS.scala 10:86]
  wire  other_ops_60_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_60_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_60_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_60_O; // @[MapS.scala 10:86]
  wire  other_ops_61_clock; // @[MapS.scala 10:86]
  wire  other_ops_61_reset; // @[MapS.scala 10:86]
  wire  other_ops_61_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_61_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_61_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_61_O; // @[MapS.scala 10:86]
  wire  other_ops_62_clock; // @[MapS.scala 10:86]
  wire  other_ops_62_reset; // @[MapS.scala 10:86]
  wire  other_ops_62_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_62_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_62_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_62_O; // @[MapS.scala 10:86]
  wire  other_ops_63_clock; // @[MapS.scala 10:86]
  wire  other_ops_63_reset; // @[MapS.scala 10:86]
  wire  other_ops_63_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_63_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_63_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_63_O; // @[MapS.scala 10:86]
  wire  other_ops_64_clock; // @[MapS.scala 10:86]
  wire  other_ops_64_reset; // @[MapS.scala 10:86]
  wire  other_ops_64_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_64_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_64_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_64_O; // @[MapS.scala 10:86]
  wire  other_ops_65_clock; // @[MapS.scala 10:86]
  wire  other_ops_65_reset; // @[MapS.scala 10:86]
  wire  other_ops_65_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_65_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_65_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_65_O; // @[MapS.scala 10:86]
  wire  other_ops_66_clock; // @[MapS.scala 10:86]
  wire  other_ops_66_reset; // @[MapS.scala 10:86]
  wire  other_ops_66_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_66_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_66_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_66_O; // @[MapS.scala 10:86]
  wire  other_ops_67_clock; // @[MapS.scala 10:86]
  wire  other_ops_67_reset; // @[MapS.scala 10:86]
  wire  other_ops_67_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_67_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_67_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_67_O; // @[MapS.scala 10:86]
  wire  other_ops_68_clock; // @[MapS.scala 10:86]
  wire  other_ops_68_reset; // @[MapS.scala 10:86]
  wire  other_ops_68_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_68_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_68_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_68_O; // @[MapS.scala 10:86]
  wire  other_ops_69_clock; // @[MapS.scala 10:86]
  wire  other_ops_69_reset; // @[MapS.scala 10:86]
  wire  other_ops_69_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_69_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_69_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_69_O; // @[MapS.scala 10:86]
  wire  other_ops_70_clock; // @[MapS.scala 10:86]
  wire  other_ops_70_reset; // @[MapS.scala 10:86]
  wire  other_ops_70_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_70_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_70_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_70_O; // @[MapS.scala 10:86]
  wire  other_ops_71_clock; // @[MapS.scala 10:86]
  wire  other_ops_71_reset; // @[MapS.scala 10:86]
  wire  other_ops_71_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_71_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_71_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_71_O; // @[MapS.scala 10:86]
  wire  other_ops_72_clock; // @[MapS.scala 10:86]
  wire  other_ops_72_reset; // @[MapS.scala 10:86]
  wire  other_ops_72_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_72_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_72_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_72_O; // @[MapS.scala 10:86]
  wire  other_ops_73_clock; // @[MapS.scala 10:86]
  wire  other_ops_73_reset; // @[MapS.scala 10:86]
  wire  other_ops_73_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_73_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_73_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_73_O; // @[MapS.scala 10:86]
  wire  other_ops_74_clock; // @[MapS.scala 10:86]
  wire  other_ops_74_reset; // @[MapS.scala 10:86]
  wire  other_ops_74_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_74_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_74_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_74_O; // @[MapS.scala 10:86]
  wire  other_ops_75_clock; // @[MapS.scala 10:86]
  wire  other_ops_75_reset; // @[MapS.scala 10:86]
  wire  other_ops_75_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_75_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_75_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_75_O; // @[MapS.scala 10:86]
  wire  other_ops_76_clock; // @[MapS.scala 10:86]
  wire  other_ops_76_reset; // @[MapS.scala 10:86]
  wire  other_ops_76_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_76_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_76_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_76_O; // @[MapS.scala 10:86]
  wire  other_ops_77_clock; // @[MapS.scala 10:86]
  wire  other_ops_77_reset; // @[MapS.scala 10:86]
  wire  other_ops_77_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_77_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_77_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_77_O; // @[MapS.scala 10:86]
  wire  other_ops_78_clock; // @[MapS.scala 10:86]
  wire  other_ops_78_reset; // @[MapS.scala 10:86]
  wire  other_ops_78_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_78_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_78_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_78_O; // @[MapS.scala 10:86]
  wire  other_ops_79_clock; // @[MapS.scala 10:86]
  wire  other_ops_79_reset; // @[MapS.scala 10:86]
  wire  other_ops_79_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_79_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_79_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_79_O; // @[MapS.scala 10:86]
  wire  other_ops_80_clock; // @[MapS.scala 10:86]
  wire  other_ops_80_reset; // @[MapS.scala 10:86]
  wire  other_ops_80_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_80_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_80_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_80_O; // @[MapS.scala 10:86]
  wire  other_ops_81_clock; // @[MapS.scala 10:86]
  wire  other_ops_81_reset; // @[MapS.scala 10:86]
  wire  other_ops_81_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_81_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_81_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_81_O; // @[MapS.scala 10:86]
  wire  other_ops_82_clock; // @[MapS.scala 10:86]
  wire  other_ops_82_reset; // @[MapS.scala 10:86]
  wire  other_ops_82_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_82_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_82_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_82_O; // @[MapS.scala 10:86]
  wire  other_ops_83_clock; // @[MapS.scala 10:86]
  wire  other_ops_83_reset; // @[MapS.scala 10:86]
  wire  other_ops_83_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_83_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_83_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_83_O; // @[MapS.scala 10:86]
  wire  other_ops_84_clock; // @[MapS.scala 10:86]
  wire  other_ops_84_reset; // @[MapS.scala 10:86]
  wire  other_ops_84_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_84_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_84_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_84_O; // @[MapS.scala 10:86]
  wire  other_ops_85_clock; // @[MapS.scala 10:86]
  wire  other_ops_85_reset; // @[MapS.scala 10:86]
  wire  other_ops_85_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_85_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_85_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_85_O; // @[MapS.scala 10:86]
  wire  other_ops_86_clock; // @[MapS.scala 10:86]
  wire  other_ops_86_reset; // @[MapS.scala 10:86]
  wire  other_ops_86_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_86_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_86_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_86_O; // @[MapS.scala 10:86]
  wire  other_ops_87_clock; // @[MapS.scala 10:86]
  wire  other_ops_87_reset; // @[MapS.scala 10:86]
  wire  other_ops_87_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_87_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_87_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_87_O; // @[MapS.scala 10:86]
  wire  other_ops_88_clock; // @[MapS.scala 10:86]
  wire  other_ops_88_reset; // @[MapS.scala 10:86]
  wire  other_ops_88_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_88_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_88_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_88_O; // @[MapS.scala 10:86]
  wire  other_ops_89_clock; // @[MapS.scala 10:86]
  wire  other_ops_89_reset; // @[MapS.scala 10:86]
  wire  other_ops_89_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_89_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_89_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_89_O; // @[MapS.scala 10:86]
  wire  other_ops_90_clock; // @[MapS.scala 10:86]
  wire  other_ops_90_reset; // @[MapS.scala 10:86]
  wire  other_ops_90_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_90_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_90_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_90_O; // @[MapS.scala 10:86]
  wire  other_ops_91_clock; // @[MapS.scala 10:86]
  wire  other_ops_91_reset; // @[MapS.scala 10:86]
  wire  other_ops_91_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_91_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_91_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_91_O; // @[MapS.scala 10:86]
  wire  other_ops_92_clock; // @[MapS.scala 10:86]
  wire  other_ops_92_reset; // @[MapS.scala 10:86]
  wire  other_ops_92_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_92_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_92_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_92_O; // @[MapS.scala 10:86]
  wire  other_ops_93_clock; // @[MapS.scala 10:86]
  wire  other_ops_93_reset; // @[MapS.scala 10:86]
  wire  other_ops_93_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_93_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_93_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_93_O; // @[MapS.scala 10:86]
  wire  other_ops_94_clock; // @[MapS.scala 10:86]
  wire  other_ops_94_reset; // @[MapS.scala 10:86]
  wire  other_ops_94_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_94_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_94_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_94_O; // @[MapS.scala 10:86]
  wire  other_ops_95_clock; // @[MapS.scala 10:86]
  wire  other_ops_95_reset; // @[MapS.scala 10:86]
  wire  other_ops_95_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_95_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_95_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_95_O; // @[MapS.scala 10:86]
  wire  other_ops_96_clock; // @[MapS.scala 10:86]
  wire  other_ops_96_reset; // @[MapS.scala 10:86]
  wire  other_ops_96_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_96_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_96_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_96_O; // @[MapS.scala 10:86]
  wire  other_ops_97_clock; // @[MapS.scala 10:86]
  wire  other_ops_97_reset; // @[MapS.scala 10:86]
  wire  other_ops_97_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_97_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_97_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_97_O; // @[MapS.scala 10:86]
  wire  other_ops_98_clock; // @[MapS.scala 10:86]
  wire  other_ops_98_reset; // @[MapS.scala 10:86]
  wire  other_ops_98_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_98_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_98_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_98_O; // @[MapS.scala 10:86]
  wire  other_ops_99_clock; // @[MapS.scala 10:86]
  wire  other_ops_99_reset; // @[MapS.scala 10:86]
  wire  other_ops_99_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_99_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_99_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_99_O; // @[MapS.scala 10:86]
  wire  other_ops_100_clock; // @[MapS.scala 10:86]
  wire  other_ops_100_reset; // @[MapS.scala 10:86]
  wire  other_ops_100_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_100_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_100_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_100_O; // @[MapS.scala 10:86]
  wire  other_ops_101_clock; // @[MapS.scala 10:86]
  wire  other_ops_101_reset; // @[MapS.scala 10:86]
  wire  other_ops_101_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_101_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_101_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_101_O; // @[MapS.scala 10:86]
  wire  other_ops_102_clock; // @[MapS.scala 10:86]
  wire  other_ops_102_reset; // @[MapS.scala 10:86]
  wire  other_ops_102_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_102_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_102_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_102_O; // @[MapS.scala 10:86]
  wire  other_ops_103_clock; // @[MapS.scala 10:86]
  wire  other_ops_103_reset; // @[MapS.scala 10:86]
  wire  other_ops_103_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_103_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_103_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_103_O; // @[MapS.scala 10:86]
  wire  other_ops_104_clock; // @[MapS.scala 10:86]
  wire  other_ops_104_reset; // @[MapS.scala 10:86]
  wire  other_ops_104_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_104_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_104_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_104_O; // @[MapS.scala 10:86]
  wire  other_ops_105_clock; // @[MapS.scala 10:86]
  wire  other_ops_105_reset; // @[MapS.scala 10:86]
  wire  other_ops_105_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_105_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_105_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_105_O; // @[MapS.scala 10:86]
  wire  other_ops_106_clock; // @[MapS.scala 10:86]
  wire  other_ops_106_reset; // @[MapS.scala 10:86]
  wire  other_ops_106_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_106_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_106_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_106_O; // @[MapS.scala 10:86]
  wire  other_ops_107_clock; // @[MapS.scala 10:86]
  wire  other_ops_107_reset; // @[MapS.scala 10:86]
  wire  other_ops_107_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_107_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_107_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_107_O; // @[MapS.scala 10:86]
  wire  other_ops_108_clock; // @[MapS.scala 10:86]
  wire  other_ops_108_reset; // @[MapS.scala 10:86]
  wire  other_ops_108_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_108_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_108_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_108_O; // @[MapS.scala 10:86]
  wire  other_ops_109_clock; // @[MapS.scala 10:86]
  wire  other_ops_109_reset; // @[MapS.scala 10:86]
  wire  other_ops_109_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_109_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_109_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_109_O; // @[MapS.scala 10:86]
  wire  other_ops_110_clock; // @[MapS.scala 10:86]
  wire  other_ops_110_reset; // @[MapS.scala 10:86]
  wire  other_ops_110_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_110_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_110_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_110_O; // @[MapS.scala 10:86]
  wire  other_ops_111_clock; // @[MapS.scala 10:86]
  wire  other_ops_111_reset; // @[MapS.scala 10:86]
  wire  other_ops_111_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_111_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_111_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_111_O; // @[MapS.scala 10:86]
  wire  other_ops_112_clock; // @[MapS.scala 10:86]
  wire  other_ops_112_reset; // @[MapS.scala 10:86]
  wire  other_ops_112_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_112_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_112_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_112_O; // @[MapS.scala 10:86]
  wire  other_ops_113_clock; // @[MapS.scala 10:86]
  wire  other_ops_113_reset; // @[MapS.scala 10:86]
  wire  other_ops_113_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_113_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_113_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_113_O; // @[MapS.scala 10:86]
  wire  other_ops_114_clock; // @[MapS.scala 10:86]
  wire  other_ops_114_reset; // @[MapS.scala 10:86]
  wire  other_ops_114_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_114_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_114_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_114_O; // @[MapS.scala 10:86]
  wire  other_ops_115_clock; // @[MapS.scala 10:86]
  wire  other_ops_115_reset; // @[MapS.scala 10:86]
  wire  other_ops_115_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_115_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_115_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_115_O; // @[MapS.scala 10:86]
  wire  other_ops_116_clock; // @[MapS.scala 10:86]
  wire  other_ops_116_reset; // @[MapS.scala 10:86]
  wire  other_ops_116_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_116_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_116_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_116_O; // @[MapS.scala 10:86]
  wire  other_ops_117_clock; // @[MapS.scala 10:86]
  wire  other_ops_117_reset; // @[MapS.scala 10:86]
  wire  other_ops_117_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_117_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_117_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_117_O; // @[MapS.scala 10:86]
  wire  other_ops_118_clock; // @[MapS.scala 10:86]
  wire  other_ops_118_reset; // @[MapS.scala 10:86]
  wire  other_ops_118_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_118_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_118_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_118_O; // @[MapS.scala 10:86]
  wire  other_ops_119_clock; // @[MapS.scala 10:86]
  wire  other_ops_119_reset; // @[MapS.scala 10:86]
  wire  other_ops_119_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_119_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_119_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_119_O; // @[MapS.scala 10:86]
  wire  other_ops_120_clock; // @[MapS.scala 10:86]
  wire  other_ops_120_reset; // @[MapS.scala 10:86]
  wire  other_ops_120_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_120_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_120_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_120_O; // @[MapS.scala 10:86]
  wire  other_ops_121_clock; // @[MapS.scala 10:86]
  wire  other_ops_121_reset; // @[MapS.scala 10:86]
  wire  other_ops_121_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_121_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_121_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_121_O; // @[MapS.scala 10:86]
  wire  other_ops_122_clock; // @[MapS.scala 10:86]
  wire  other_ops_122_reset; // @[MapS.scala 10:86]
  wire  other_ops_122_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_122_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_122_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_122_O; // @[MapS.scala 10:86]
  wire  other_ops_123_clock; // @[MapS.scala 10:86]
  wire  other_ops_123_reset; // @[MapS.scala 10:86]
  wire  other_ops_123_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_123_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_123_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_123_O; // @[MapS.scala 10:86]
  wire  other_ops_124_clock; // @[MapS.scala 10:86]
  wire  other_ops_124_reset; // @[MapS.scala 10:86]
  wire  other_ops_124_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_124_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_124_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_124_O; // @[MapS.scala 10:86]
  wire  other_ops_125_clock; // @[MapS.scala 10:86]
  wire  other_ops_125_reset; // @[MapS.scala 10:86]
  wire  other_ops_125_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_125_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_125_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_125_O; // @[MapS.scala 10:86]
  wire  other_ops_126_clock; // @[MapS.scala 10:86]
  wire  other_ops_126_reset; // @[MapS.scala 10:86]
  wire  other_ops_126_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_126_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_126_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_126_O; // @[MapS.scala 10:86]
  wire  other_ops_127_clock; // @[MapS.scala 10:86]
  wire  other_ops_127_reset; // @[MapS.scala 10:86]
  wire  other_ops_127_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_127_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_127_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_127_O; // @[MapS.scala 10:86]
  wire  other_ops_128_clock; // @[MapS.scala 10:86]
  wire  other_ops_128_reset; // @[MapS.scala 10:86]
  wire  other_ops_128_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_128_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_128_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_128_O; // @[MapS.scala 10:86]
  wire  other_ops_129_clock; // @[MapS.scala 10:86]
  wire  other_ops_129_reset; // @[MapS.scala 10:86]
  wire  other_ops_129_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_129_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_129_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_129_O; // @[MapS.scala 10:86]
  wire  other_ops_130_clock; // @[MapS.scala 10:86]
  wire  other_ops_130_reset; // @[MapS.scala 10:86]
  wire  other_ops_130_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_130_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_130_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_130_O; // @[MapS.scala 10:86]
  wire  other_ops_131_clock; // @[MapS.scala 10:86]
  wire  other_ops_131_reset; // @[MapS.scala 10:86]
  wire  other_ops_131_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_131_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_131_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_131_O; // @[MapS.scala 10:86]
  wire  other_ops_132_clock; // @[MapS.scala 10:86]
  wire  other_ops_132_reset; // @[MapS.scala 10:86]
  wire  other_ops_132_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_132_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_132_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_132_O; // @[MapS.scala 10:86]
  wire  other_ops_133_clock; // @[MapS.scala 10:86]
  wire  other_ops_133_reset; // @[MapS.scala 10:86]
  wire  other_ops_133_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_133_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_133_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_133_O; // @[MapS.scala 10:86]
  wire  other_ops_134_clock; // @[MapS.scala 10:86]
  wire  other_ops_134_reset; // @[MapS.scala 10:86]
  wire  other_ops_134_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_134_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_134_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_134_O; // @[MapS.scala 10:86]
  wire  other_ops_135_clock; // @[MapS.scala 10:86]
  wire  other_ops_135_reset; // @[MapS.scala 10:86]
  wire  other_ops_135_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_135_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_135_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_135_O; // @[MapS.scala 10:86]
  wire  other_ops_136_clock; // @[MapS.scala 10:86]
  wire  other_ops_136_reset; // @[MapS.scala 10:86]
  wire  other_ops_136_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_136_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_136_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_136_O; // @[MapS.scala 10:86]
  wire  other_ops_137_clock; // @[MapS.scala 10:86]
  wire  other_ops_137_reset; // @[MapS.scala 10:86]
  wire  other_ops_137_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_137_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_137_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_137_O; // @[MapS.scala 10:86]
  wire  other_ops_138_clock; // @[MapS.scala 10:86]
  wire  other_ops_138_reset; // @[MapS.scala 10:86]
  wire  other_ops_138_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_138_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_138_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_138_O; // @[MapS.scala 10:86]
  wire  other_ops_139_clock; // @[MapS.scala 10:86]
  wire  other_ops_139_reset; // @[MapS.scala 10:86]
  wire  other_ops_139_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_139_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_139_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_139_O; // @[MapS.scala 10:86]
  wire  other_ops_140_clock; // @[MapS.scala 10:86]
  wire  other_ops_140_reset; // @[MapS.scala 10:86]
  wire  other_ops_140_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_140_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_140_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_140_O; // @[MapS.scala 10:86]
  wire  other_ops_141_clock; // @[MapS.scala 10:86]
  wire  other_ops_141_reset; // @[MapS.scala 10:86]
  wire  other_ops_141_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_141_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_141_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_141_O; // @[MapS.scala 10:86]
  wire  other_ops_142_clock; // @[MapS.scala 10:86]
  wire  other_ops_142_reset; // @[MapS.scala 10:86]
  wire  other_ops_142_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_142_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_142_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_142_O; // @[MapS.scala 10:86]
  wire  other_ops_143_clock; // @[MapS.scala 10:86]
  wire  other_ops_143_reset; // @[MapS.scala 10:86]
  wire  other_ops_143_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_143_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_143_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_143_O; // @[MapS.scala 10:86]
  wire  other_ops_144_clock; // @[MapS.scala 10:86]
  wire  other_ops_144_reset; // @[MapS.scala 10:86]
  wire  other_ops_144_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_144_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_144_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_144_O; // @[MapS.scala 10:86]
  wire  other_ops_145_clock; // @[MapS.scala 10:86]
  wire  other_ops_145_reset; // @[MapS.scala 10:86]
  wire  other_ops_145_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_145_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_145_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_145_O; // @[MapS.scala 10:86]
  wire  other_ops_146_clock; // @[MapS.scala 10:86]
  wire  other_ops_146_reset; // @[MapS.scala 10:86]
  wire  other_ops_146_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_146_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_146_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_146_O; // @[MapS.scala 10:86]
  wire  other_ops_147_clock; // @[MapS.scala 10:86]
  wire  other_ops_147_reset; // @[MapS.scala 10:86]
  wire  other_ops_147_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_147_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_147_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_147_O; // @[MapS.scala 10:86]
  wire  other_ops_148_clock; // @[MapS.scala 10:86]
  wire  other_ops_148_reset; // @[MapS.scala 10:86]
  wire  other_ops_148_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_148_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_148_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_148_O; // @[MapS.scala 10:86]
  wire  other_ops_149_clock; // @[MapS.scala 10:86]
  wire  other_ops_149_reset; // @[MapS.scala 10:86]
  wire  other_ops_149_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_149_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_149_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_149_O; // @[MapS.scala 10:86]
  wire  other_ops_150_clock; // @[MapS.scala 10:86]
  wire  other_ops_150_reset; // @[MapS.scala 10:86]
  wire  other_ops_150_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_150_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_150_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_150_O; // @[MapS.scala 10:86]
  wire  other_ops_151_clock; // @[MapS.scala 10:86]
  wire  other_ops_151_reset; // @[MapS.scala 10:86]
  wire  other_ops_151_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_151_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_151_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_151_O; // @[MapS.scala 10:86]
  wire  other_ops_152_clock; // @[MapS.scala 10:86]
  wire  other_ops_152_reset; // @[MapS.scala 10:86]
  wire  other_ops_152_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_152_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_152_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_152_O; // @[MapS.scala 10:86]
  wire  other_ops_153_clock; // @[MapS.scala 10:86]
  wire  other_ops_153_reset; // @[MapS.scala 10:86]
  wire  other_ops_153_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_153_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_153_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_153_O; // @[MapS.scala 10:86]
  wire  other_ops_154_clock; // @[MapS.scala 10:86]
  wire  other_ops_154_reset; // @[MapS.scala 10:86]
  wire  other_ops_154_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_154_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_154_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_154_O; // @[MapS.scala 10:86]
  wire  other_ops_155_clock; // @[MapS.scala 10:86]
  wire  other_ops_155_reset; // @[MapS.scala 10:86]
  wire  other_ops_155_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_155_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_155_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_155_O; // @[MapS.scala 10:86]
  wire  other_ops_156_clock; // @[MapS.scala 10:86]
  wire  other_ops_156_reset; // @[MapS.scala 10:86]
  wire  other_ops_156_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_156_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_156_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_156_O; // @[MapS.scala 10:86]
  wire  other_ops_157_clock; // @[MapS.scala 10:86]
  wire  other_ops_157_reset; // @[MapS.scala 10:86]
  wire  other_ops_157_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_157_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_157_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_157_O; // @[MapS.scala 10:86]
  wire  other_ops_158_clock; // @[MapS.scala 10:86]
  wire  other_ops_158_reset; // @[MapS.scala 10:86]
  wire  other_ops_158_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_158_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_158_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_158_O; // @[MapS.scala 10:86]
  wire  other_ops_159_clock; // @[MapS.scala 10:86]
  wire  other_ops_159_reset; // @[MapS.scala 10:86]
  wire  other_ops_159_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_159_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_159_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_159_O; // @[MapS.scala 10:86]
  wire  other_ops_160_clock; // @[MapS.scala 10:86]
  wire  other_ops_160_reset; // @[MapS.scala 10:86]
  wire  other_ops_160_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_160_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_160_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_160_O; // @[MapS.scala 10:86]
  wire  other_ops_161_clock; // @[MapS.scala 10:86]
  wire  other_ops_161_reset; // @[MapS.scala 10:86]
  wire  other_ops_161_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_161_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_161_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_161_O; // @[MapS.scala 10:86]
  wire  other_ops_162_clock; // @[MapS.scala 10:86]
  wire  other_ops_162_reset; // @[MapS.scala 10:86]
  wire  other_ops_162_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_162_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_162_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_162_O; // @[MapS.scala 10:86]
  wire  other_ops_163_clock; // @[MapS.scala 10:86]
  wire  other_ops_163_reset; // @[MapS.scala 10:86]
  wire  other_ops_163_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_163_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_163_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_163_O; // @[MapS.scala 10:86]
  wire  other_ops_164_clock; // @[MapS.scala 10:86]
  wire  other_ops_164_reset; // @[MapS.scala 10:86]
  wire  other_ops_164_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_164_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_164_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_164_O; // @[MapS.scala 10:86]
  wire  other_ops_165_clock; // @[MapS.scala 10:86]
  wire  other_ops_165_reset; // @[MapS.scala 10:86]
  wire  other_ops_165_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_165_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_165_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_165_O; // @[MapS.scala 10:86]
  wire  other_ops_166_clock; // @[MapS.scala 10:86]
  wire  other_ops_166_reset; // @[MapS.scala 10:86]
  wire  other_ops_166_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_166_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_166_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_166_O; // @[MapS.scala 10:86]
  wire  other_ops_167_clock; // @[MapS.scala 10:86]
  wire  other_ops_167_reset; // @[MapS.scala 10:86]
  wire  other_ops_167_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_167_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_167_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_167_O; // @[MapS.scala 10:86]
  wire  other_ops_168_clock; // @[MapS.scala 10:86]
  wire  other_ops_168_reset; // @[MapS.scala 10:86]
  wire  other_ops_168_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_168_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_168_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_168_O; // @[MapS.scala 10:86]
  wire  other_ops_169_clock; // @[MapS.scala 10:86]
  wire  other_ops_169_reset; // @[MapS.scala 10:86]
  wire  other_ops_169_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_169_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_169_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_169_O; // @[MapS.scala 10:86]
  wire  other_ops_170_clock; // @[MapS.scala 10:86]
  wire  other_ops_170_reset; // @[MapS.scala 10:86]
  wire  other_ops_170_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_170_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_170_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_170_O; // @[MapS.scala 10:86]
  wire  other_ops_171_clock; // @[MapS.scala 10:86]
  wire  other_ops_171_reset; // @[MapS.scala 10:86]
  wire  other_ops_171_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_171_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_171_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_171_O; // @[MapS.scala 10:86]
  wire  other_ops_172_clock; // @[MapS.scala 10:86]
  wire  other_ops_172_reset; // @[MapS.scala 10:86]
  wire  other_ops_172_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_172_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_172_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_172_O; // @[MapS.scala 10:86]
  wire  other_ops_173_clock; // @[MapS.scala 10:86]
  wire  other_ops_173_reset; // @[MapS.scala 10:86]
  wire  other_ops_173_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_173_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_173_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_173_O; // @[MapS.scala 10:86]
  wire  other_ops_174_clock; // @[MapS.scala 10:86]
  wire  other_ops_174_reset; // @[MapS.scala 10:86]
  wire  other_ops_174_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_174_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_174_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_174_O; // @[MapS.scala 10:86]
  wire  other_ops_175_clock; // @[MapS.scala 10:86]
  wire  other_ops_175_reset; // @[MapS.scala 10:86]
  wire  other_ops_175_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_175_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_175_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_175_O; // @[MapS.scala 10:86]
  wire  other_ops_176_clock; // @[MapS.scala 10:86]
  wire  other_ops_176_reset; // @[MapS.scala 10:86]
  wire  other_ops_176_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_176_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_176_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_176_O; // @[MapS.scala 10:86]
  wire  other_ops_177_clock; // @[MapS.scala 10:86]
  wire  other_ops_177_reset; // @[MapS.scala 10:86]
  wire  other_ops_177_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_177_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_177_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_177_O; // @[MapS.scala 10:86]
  wire  other_ops_178_clock; // @[MapS.scala 10:86]
  wire  other_ops_178_reset; // @[MapS.scala 10:86]
  wire  other_ops_178_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_178_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_178_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_178_O; // @[MapS.scala 10:86]
  wire  other_ops_179_clock; // @[MapS.scala 10:86]
  wire  other_ops_179_reset; // @[MapS.scala 10:86]
  wire  other_ops_179_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_179_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_179_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_179_O; // @[MapS.scala 10:86]
  wire  other_ops_180_clock; // @[MapS.scala 10:86]
  wire  other_ops_180_reset; // @[MapS.scala 10:86]
  wire  other_ops_180_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_180_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_180_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_180_O; // @[MapS.scala 10:86]
  wire  other_ops_181_clock; // @[MapS.scala 10:86]
  wire  other_ops_181_reset; // @[MapS.scala 10:86]
  wire  other_ops_181_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_181_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_181_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_181_O; // @[MapS.scala 10:86]
  wire  other_ops_182_clock; // @[MapS.scala 10:86]
  wire  other_ops_182_reset; // @[MapS.scala 10:86]
  wire  other_ops_182_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_182_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_182_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_182_O; // @[MapS.scala 10:86]
  wire  other_ops_183_clock; // @[MapS.scala 10:86]
  wire  other_ops_183_reset; // @[MapS.scala 10:86]
  wire  other_ops_183_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_183_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_183_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_183_O; // @[MapS.scala 10:86]
  wire  other_ops_184_clock; // @[MapS.scala 10:86]
  wire  other_ops_184_reset; // @[MapS.scala 10:86]
  wire  other_ops_184_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_184_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_184_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_184_O; // @[MapS.scala 10:86]
  wire  other_ops_185_clock; // @[MapS.scala 10:86]
  wire  other_ops_185_reset; // @[MapS.scala 10:86]
  wire  other_ops_185_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_185_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_185_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_185_O; // @[MapS.scala 10:86]
  wire  other_ops_186_clock; // @[MapS.scala 10:86]
  wire  other_ops_186_reset; // @[MapS.scala 10:86]
  wire  other_ops_186_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_186_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_186_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_186_O; // @[MapS.scala 10:86]
  wire  other_ops_187_clock; // @[MapS.scala 10:86]
  wire  other_ops_187_reset; // @[MapS.scala 10:86]
  wire  other_ops_187_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_187_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_187_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_187_O; // @[MapS.scala 10:86]
  wire  other_ops_188_clock; // @[MapS.scala 10:86]
  wire  other_ops_188_reset; // @[MapS.scala 10:86]
  wire  other_ops_188_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_188_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_188_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_188_O; // @[MapS.scala 10:86]
  wire  other_ops_189_clock; // @[MapS.scala 10:86]
  wire  other_ops_189_reset; // @[MapS.scala 10:86]
  wire  other_ops_189_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_189_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_189_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_189_O; // @[MapS.scala 10:86]
  wire  other_ops_190_clock; // @[MapS.scala 10:86]
  wire  other_ops_190_reset; // @[MapS.scala 10:86]
  wire  other_ops_190_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_190_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_190_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_190_O; // @[MapS.scala 10:86]
  wire  other_ops_191_clock; // @[MapS.scala 10:86]
  wire  other_ops_191_reset; // @[MapS.scala 10:86]
  wire  other_ops_191_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_191_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_191_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_191_O; // @[MapS.scala 10:86]
  wire  other_ops_192_clock; // @[MapS.scala 10:86]
  wire  other_ops_192_reset; // @[MapS.scala 10:86]
  wire  other_ops_192_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_192_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_192_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_192_O; // @[MapS.scala 10:86]
  wire  other_ops_193_clock; // @[MapS.scala 10:86]
  wire  other_ops_193_reset; // @[MapS.scala 10:86]
  wire  other_ops_193_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_193_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_193_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_193_O; // @[MapS.scala 10:86]
  wire  other_ops_194_clock; // @[MapS.scala 10:86]
  wire  other_ops_194_reset; // @[MapS.scala 10:86]
  wire  other_ops_194_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_194_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_194_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_194_O; // @[MapS.scala 10:86]
  wire  other_ops_195_clock; // @[MapS.scala 10:86]
  wire  other_ops_195_reset; // @[MapS.scala 10:86]
  wire  other_ops_195_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_195_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_195_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_195_O; // @[MapS.scala 10:86]
  wire  other_ops_196_clock; // @[MapS.scala 10:86]
  wire  other_ops_196_reset; // @[MapS.scala 10:86]
  wire  other_ops_196_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_196_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_196_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_196_O; // @[MapS.scala 10:86]
  wire  other_ops_197_clock; // @[MapS.scala 10:86]
  wire  other_ops_197_reset; // @[MapS.scala 10:86]
  wire  other_ops_197_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_197_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_197_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_197_O; // @[MapS.scala 10:86]
  wire  other_ops_198_clock; // @[MapS.scala 10:86]
  wire  other_ops_198_reset; // @[MapS.scala 10:86]
  wire  other_ops_198_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_198_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_198_I; // @[MapS.scala 10:86]
  wire [7:0] other_ops_198_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  wire  _T_14; // @[MapS.scala 23:83]
  wire  _T_15; // @[MapS.scala 23:83]
  wire  _T_16; // @[MapS.scala 23:83]
  wire  _T_17; // @[MapS.scala 23:83]
  wire  _T_18; // @[MapS.scala 23:83]
  wire  _T_19; // @[MapS.scala 23:83]
  wire  _T_20; // @[MapS.scala 23:83]
  wire  _T_21; // @[MapS.scala 23:83]
  wire  _T_22; // @[MapS.scala 23:83]
  wire  _T_23; // @[MapS.scala 23:83]
  wire  _T_24; // @[MapS.scala 23:83]
  wire  _T_25; // @[MapS.scala 23:83]
  wire  _T_26; // @[MapS.scala 23:83]
  wire  _T_27; // @[MapS.scala 23:83]
  wire  _T_28; // @[MapS.scala 23:83]
  wire  _T_29; // @[MapS.scala 23:83]
  wire  _T_30; // @[MapS.scala 23:83]
  wire  _T_31; // @[MapS.scala 23:83]
  wire  _T_32; // @[MapS.scala 23:83]
  wire  _T_33; // @[MapS.scala 23:83]
  wire  _T_34; // @[MapS.scala 23:83]
  wire  _T_35; // @[MapS.scala 23:83]
  wire  _T_36; // @[MapS.scala 23:83]
  wire  _T_37; // @[MapS.scala 23:83]
  wire  _T_38; // @[MapS.scala 23:83]
  wire  _T_39; // @[MapS.scala 23:83]
  wire  _T_40; // @[MapS.scala 23:83]
  wire  _T_41; // @[MapS.scala 23:83]
  wire  _T_42; // @[MapS.scala 23:83]
  wire  _T_43; // @[MapS.scala 23:83]
  wire  _T_44; // @[MapS.scala 23:83]
  wire  _T_45; // @[MapS.scala 23:83]
  wire  _T_46; // @[MapS.scala 23:83]
  wire  _T_47; // @[MapS.scala 23:83]
  wire  _T_48; // @[MapS.scala 23:83]
  wire  _T_49; // @[MapS.scala 23:83]
  wire  _T_50; // @[MapS.scala 23:83]
  wire  _T_51; // @[MapS.scala 23:83]
  wire  _T_52; // @[MapS.scala 23:83]
  wire  _T_53; // @[MapS.scala 23:83]
  wire  _T_54; // @[MapS.scala 23:83]
  wire  _T_55; // @[MapS.scala 23:83]
  wire  _T_56; // @[MapS.scala 23:83]
  wire  _T_57; // @[MapS.scala 23:83]
  wire  _T_58; // @[MapS.scala 23:83]
  wire  _T_59; // @[MapS.scala 23:83]
  wire  _T_60; // @[MapS.scala 23:83]
  wire  _T_61; // @[MapS.scala 23:83]
  wire  _T_62; // @[MapS.scala 23:83]
  wire  _T_63; // @[MapS.scala 23:83]
  wire  _T_64; // @[MapS.scala 23:83]
  wire  _T_65; // @[MapS.scala 23:83]
  wire  _T_66; // @[MapS.scala 23:83]
  wire  _T_67; // @[MapS.scala 23:83]
  wire  _T_68; // @[MapS.scala 23:83]
  wire  _T_69; // @[MapS.scala 23:83]
  wire  _T_70; // @[MapS.scala 23:83]
  wire  _T_71; // @[MapS.scala 23:83]
  wire  _T_72; // @[MapS.scala 23:83]
  wire  _T_73; // @[MapS.scala 23:83]
  wire  _T_74; // @[MapS.scala 23:83]
  wire  _T_75; // @[MapS.scala 23:83]
  wire  _T_76; // @[MapS.scala 23:83]
  wire  _T_77; // @[MapS.scala 23:83]
  wire  _T_78; // @[MapS.scala 23:83]
  wire  _T_79; // @[MapS.scala 23:83]
  wire  _T_80; // @[MapS.scala 23:83]
  wire  _T_81; // @[MapS.scala 23:83]
  wire  _T_82; // @[MapS.scala 23:83]
  wire  _T_83; // @[MapS.scala 23:83]
  wire  _T_84; // @[MapS.scala 23:83]
  wire  _T_85; // @[MapS.scala 23:83]
  wire  _T_86; // @[MapS.scala 23:83]
  wire  _T_87; // @[MapS.scala 23:83]
  wire  _T_88; // @[MapS.scala 23:83]
  wire  _T_89; // @[MapS.scala 23:83]
  wire  _T_90; // @[MapS.scala 23:83]
  wire  _T_91; // @[MapS.scala 23:83]
  wire  _T_92; // @[MapS.scala 23:83]
  wire  _T_93; // @[MapS.scala 23:83]
  wire  _T_94; // @[MapS.scala 23:83]
  wire  _T_95; // @[MapS.scala 23:83]
  wire  _T_96; // @[MapS.scala 23:83]
  wire  _T_97; // @[MapS.scala 23:83]
  wire  _T_98; // @[MapS.scala 23:83]
  wire  _T_99; // @[MapS.scala 23:83]
  wire  _T_100; // @[MapS.scala 23:83]
  wire  _T_101; // @[MapS.scala 23:83]
  wire  _T_102; // @[MapS.scala 23:83]
  wire  _T_103; // @[MapS.scala 23:83]
  wire  _T_104; // @[MapS.scala 23:83]
  wire  _T_105; // @[MapS.scala 23:83]
  wire  _T_106; // @[MapS.scala 23:83]
  wire  _T_107; // @[MapS.scala 23:83]
  wire  _T_108; // @[MapS.scala 23:83]
  wire  _T_109; // @[MapS.scala 23:83]
  wire  _T_110; // @[MapS.scala 23:83]
  wire  _T_111; // @[MapS.scala 23:83]
  wire  _T_112; // @[MapS.scala 23:83]
  wire  _T_113; // @[MapS.scala 23:83]
  wire  _T_114; // @[MapS.scala 23:83]
  wire  _T_115; // @[MapS.scala 23:83]
  wire  _T_116; // @[MapS.scala 23:83]
  wire  _T_117; // @[MapS.scala 23:83]
  wire  _T_118; // @[MapS.scala 23:83]
  wire  _T_119; // @[MapS.scala 23:83]
  wire  _T_120; // @[MapS.scala 23:83]
  wire  _T_121; // @[MapS.scala 23:83]
  wire  _T_122; // @[MapS.scala 23:83]
  wire  _T_123; // @[MapS.scala 23:83]
  wire  _T_124; // @[MapS.scala 23:83]
  wire  _T_125; // @[MapS.scala 23:83]
  wire  _T_126; // @[MapS.scala 23:83]
  wire  _T_127; // @[MapS.scala 23:83]
  wire  _T_128; // @[MapS.scala 23:83]
  wire  _T_129; // @[MapS.scala 23:83]
  wire  _T_130; // @[MapS.scala 23:83]
  wire  _T_131; // @[MapS.scala 23:83]
  wire  _T_132; // @[MapS.scala 23:83]
  wire  _T_133; // @[MapS.scala 23:83]
  wire  _T_134; // @[MapS.scala 23:83]
  wire  _T_135; // @[MapS.scala 23:83]
  wire  _T_136; // @[MapS.scala 23:83]
  wire  _T_137; // @[MapS.scala 23:83]
  wire  _T_138; // @[MapS.scala 23:83]
  wire  _T_139; // @[MapS.scala 23:83]
  wire  _T_140; // @[MapS.scala 23:83]
  wire  _T_141; // @[MapS.scala 23:83]
  wire  _T_142; // @[MapS.scala 23:83]
  wire  _T_143; // @[MapS.scala 23:83]
  wire  _T_144; // @[MapS.scala 23:83]
  wire  _T_145; // @[MapS.scala 23:83]
  wire  _T_146; // @[MapS.scala 23:83]
  wire  _T_147; // @[MapS.scala 23:83]
  wire  _T_148; // @[MapS.scala 23:83]
  wire  _T_149; // @[MapS.scala 23:83]
  wire  _T_150; // @[MapS.scala 23:83]
  wire  _T_151; // @[MapS.scala 23:83]
  wire  _T_152; // @[MapS.scala 23:83]
  wire  _T_153; // @[MapS.scala 23:83]
  wire  _T_154; // @[MapS.scala 23:83]
  wire  _T_155; // @[MapS.scala 23:83]
  wire  _T_156; // @[MapS.scala 23:83]
  wire  _T_157; // @[MapS.scala 23:83]
  wire  _T_158; // @[MapS.scala 23:83]
  wire  _T_159; // @[MapS.scala 23:83]
  wire  _T_160; // @[MapS.scala 23:83]
  wire  _T_161; // @[MapS.scala 23:83]
  wire  _T_162; // @[MapS.scala 23:83]
  wire  _T_163; // @[MapS.scala 23:83]
  wire  _T_164; // @[MapS.scala 23:83]
  wire  _T_165; // @[MapS.scala 23:83]
  wire  _T_166; // @[MapS.scala 23:83]
  wire  _T_167; // @[MapS.scala 23:83]
  wire  _T_168; // @[MapS.scala 23:83]
  wire  _T_169; // @[MapS.scala 23:83]
  wire  _T_170; // @[MapS.scala 23:83]
  wire  _T_171; // @[MapS.scala 23:83]
  wire  _T_172; // @[MapS.scala 23:83]
  wire  _T_173; // @[MapS.scala 23:83]
  wire  _T_174; // @[MapS.scala 23:83]
  wire  _T_175; // @[MapS.scala 23:83]
  wire  _T_176; // @[MapS.scala 23:83]
  wire  _T_177; // @[MapS.scala 23:83]
  wire  _T_178; // @[MapS.scala 23:83]
  wire  _T_179; // @[MapS.scala 23:83]
  wire  _T_180; // @[MapS.scala 23:83]
  wire  _T_181; // @[MapS.scala 23:83]
  wire  _T_182; // @[MapS.scala 23:83]
  wire  _T_183; // @[MapS.scala 23:83]
  wire  _T_184; // @[MapS.scala 23:83]
  wire  _T_185; // @[MapS.scala 23:83]
  wire  _T_186; // @[MapS.scala 23:83]
  wire  _T_187; // @[MapS.scala 23:83]
  wire  _T_188; // @[MapS.scala 23:83]
  wire  _T_189; // @[MapS.scala 23:83]
  wire  _T_190; // @[MapS.scala 23:83]
  wire  _T_191; // @[MapS.scala 23:83]
  wire  _T_192; // @[MapS.scala 23:83]
  wire  _T_193; // @[MapS.scala 23:83]
  wire  _T_194; // @[MapS.scala 23:83]
  wire  _T_195; // @[MapS.scala 23:83]
  wire  _T_196; // @[MapS.scala 23:83]
  wire  _T_197; // @[MapS.scala 23:83]
  Module_0 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I(fst_op_I),
    .O(fst_op_O)
  );
  Module_0 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I(other_ops_0_I),
    .O(other_ops_0_O)
  );
  Module_0 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I(other_ops_1_I),
    .O(other_ops_1_O)
  );
  Module_0 other_ops_2 ( // @[MapS.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I(other_ops_2_I),
    .O(other_ops_2_O)
  );
  Module_0 other_ops_3 ( // @[MapS.scala 10:86]
    .clock(other_ops_3_clock),
    .reset(other_ops_3_reset),
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I(other_ops_3_I),
    .O(other_ops_3_O)
  );
  Module_0 other_ops_4 ( // @[MapS.scala 10:86]
    .clock(other_ops_4_clock),
    .reset(other_ops_4_reset),
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I(other_ops_4_I),
    .O(other_ops_4_O)
  );
  Module_0 other_ops_5 ( // @[MapS.scala 10:86]
    .clock(other_ops_5_clock),
    .reset(other_ops_5_reset),
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I(other_ops_5_I),
    .O(other_ops_5_O)
  );
  Module_0 other_ops_6 ( // @[MapS.scala 10:86]
    .clock(other_ops_6_clock),
    .reset(other_ops_6_reset),
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I(other_ops_6_I),
    .O(other_ops_6_O)
  );
  Module_0 other_ops_7 ( // @[MapS.scala 10:86]
    .clock(other_ops_7_clock),
    .reset(other_ops_7_reset),
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I(other_ops_7_I),
    .O(other_ops_7_O)
  );
  Module_0 other_ops_8 ( // @[MapS.scala 10:86]
    .clock(other_ops_8_clock),
    .reset(other_ops_8_reset),
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I(other_ops_8_I),
    .O(other_ops_8_O)
  );
  Module_0 other_ops_9 ( // @[MapS.scala 10:86]
    .clock(other_ops_9_clock),
    .reset(other_ops_9_reset),
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I(other_ops_9_I),
    .O(other_ops_9_O)
  );
  Module_0 other_ops_10 ( // @[MapS.scala 10:86]
    .clock(other_ops_10_clock),
    .reset(other_ops_10_reset),
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I(other_ops_10_I),
    .O(other_ops_10_O)
  );
  Module_0 other_ops_11 ( // @[MapS.scala 10:86]
    .clock(other_ops_11_clock),
    .reset(other_ops_11_reset),
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I(other_ops_11_I),
    .O(other_ops_11_O)
  );
  Module_0 other_ops_12 ( // @[MapS.scala 10:86]
    .clock(other_ops_12_clock),
    .reset(other_ops_12_reset),
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I(other_ops_12_I),
    .O(other_ops_12_O)
  );
  Module_0 other_ops_13 ( // @[MapS.scala 10:86]
    .clock(other_ops_13_clock),
    .reset(other_ops_13_reset),
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I(other_ops_13_I),
    .O(other_ops_13_O)
  );
  Module_0 other_ops_14 ( // @[MapS.scala 10:86]
    .clock(other_ops_14_clock),
    .reset(other_ops_14_reset),
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I(other_ops_14_I),
    .O(other_ops_14_O)
  );
  Module_0 other_ops_15 ( // @[MapS.scala 10:86]
    .clock(other_ops_15_clock),
    .reset(other_ops_15_reset),
    .valid_up(other_ops_15_valid_up),
    .valid_down(other_ops_15_valid_down),
    .I(other_ops_15_I),
    .O(other_ops_15_O)
  );
  Module_0 other_ops_16 ( // @[MapS.scala 10:86]
    .clock(other_ops_16_clock),
    .reset(other_ops_16_reset),
    .valid_up(other_ops_16_valid_up),
    .valid_down(other_ops_16_valid_down),
    .I(other_ops_16_I),
    .O(other_ops_16_O)
  );
  Module_0 other_ops_17 ( // @[MapS.scala 10:86]
    .clock(other_ops_17_clock),
    .reset(other_ops_17_reset),
    .valid_up(other_ops_17_valid_up),
    .valid_down(other_ops_17_valid_down),
    .I(other_ops_17_I),
    .O(other_ops_17_O)
  );
  Module_0 other_ops_18 ( // @[MapS.scala 10:86]
    .clock(other_ops_18_clock),
    .reset(other_ops_18_reset),
    .valid_up(other_ops_18_valid_up),
    .valid_down(other_ops_18_valid_down),
    .I(other_ops_18_I),
    .O(other_ops_18_O)
  );
  Module_0 other_ops_19 ( // @[MapS.scala 10:86]
    .clock(other_ops_19_clock),
    .reset(other_ops_19_reset),
    .valid_up(other_ops_19_valid_up),
    .valid_down(other_ops_19_valid_down),
    .I(other_ops_19_I),
    .O(other_ops_19_O)
  );
  Module_0 other_ops_20 ( // @[MapS.scala 10:86]
    .clock(other_ops_20_clock),
    .reset(other_ops_20_reset),
    .valid_up(other_ops_20_valid_up),
    .valid_down(other_ops_20_valid_down),
    .I(other_ops_20_I),
    .O(other_ops_20_O)
  );
  Module_0 other_ops_21 ( // @[MapS.scala 10:86]
    .clock(other_ops_21_clock),
    .reset(other_ops_21_reset),
    .valid_up(other_ops_21_valid_up),
    .valid_down(other_ops_21_valid_down),
    .I(other_ops_21_I),
    .O(other_ops_21_O)
  );
  Module_0 other_ops_22 ( // @[MapS.scala 10:86]
    .clock(other_ops_22_clock),
    .reset(other_ops_22_reset),
    .valid_up(other_ops_22_valid_up),
    .valid_down(other_ops_22_valid_down),
    .I(other_ops_22_I),
    .O(other_ops_22_O)
  );
  Module_0 other_ops_23 ( // @[MapS.scala 10:86]
    .clock(other_ops_23_clock),
    .reset(other_ops_23_reset),
    .valid_up(other_ops_23_valid_up),
    .valid_down(other_ops_23_valid_down),
    .I(other_ops_23_I),
    .O(other_ops_23_O)
  );
  Module_0 other_ops_24 ( // @[MapS.scala 10:86]
    .clock(other_ops_24_clock),
    .reset(other_ops_24_reset),
    .valid_up(other_ops_24_valid_up),
    .valid_down(other_ops_24_valid_down),
    .I(other_ops_24_I),
    .O(other_ops_24_O)
  );
  Module_0 other_ops_25 ( // @[MapS.scala 10:86]
    .clock(other_ops_25_clock),
    .reset(other_ops_25_reset),
    .valid_up(other_ops_25_valid_up),
    .valid_down(other_ops_25_valid_down),
    .I(other_ops_25_I),
    .O(other_ops_25_O)
  );
  Module_0 other_ops_26 ( // @[MapS.scala 10:86]
    .clock(other_ops_26_clock),
    .reset(other_ops_26_reset),
    .valid_up(other_ops_26_valid_up),
    .valid_down(other_ops_26_valid_down),
    .I(other_ops_26_I),
    .O(other_ops_26_O)
  );
  Module_0 other_ops_27 ( // @[MapS.scala 10:86]
    .clock(other_ops_27_clock),
    .reset(other_ops_27_reset),
    .valid_up(other_ops_27_valid_up),
    .valid_down(other_ops_27_valid_down),
    .I(other_ops_27_I),
    .O(other_ops_27_O)
  );
  Module_0 other_ops_28 ( // @[MapS.scala 10:86]
    .clock(other_ops_28_clock),
    .reset(other_ops_28_reset),
    .valid_up(other_ops_28_valid_up),
    .valid_down(other_ops_28_valid_down),
    .I(other_ops_28_I),
    .O(other_ops_28_O)
  );
  Module_0 other_ops_29 ( // @[MapS.scala 10:86]
    .clock(other_ops_29_clock),
    .reset(other_ops_29_reset),
    .valid_up(other_ops_29_valid_up),
    .valid_down(other_ops_29_valid_down),
    .I(other_ops_29_I),
    .O(other_ops_29_O)
  );
  Module_0 other_ops_30 ( // @[MapS.scala 10:86]
    .clock(other_ops_30_clock),
    .reset(other_ops_30_reset),
    .valid_up(other_ops_30_valid_up),
    .valid_down(other_ops_30_valid_down),
    .I(other_ops_30_I),
    .O(other_ops_30_O)
  );
  Module_0 other_ops_31 ( // @[MapS.scala 10:86]
    .clock(other_ops_31_clock),
    .reset(other_ops_31_reset),
    .valid_up(other_ops_31_valid_up),
    .valid_down(other_ops_31_valid_down),
    .I(other_ops_31_I),
    .O(other_ops_31_O)
  );
  Module_0 other_ops_32 ( // @[MapS.scala 10:86]
    .clock(other_ops_32_clock),
    .reset(other_ops_32_reset),
    .valid_up(other_ops_32_valid_up),
    .valid_down(other_ops_32_valid_down),
    .I(other_ops_32_I),
    .O(other_ops_32_O)
  );
  Module_0 other_ops_33 ( // @[MapS.scala 10:86]
    .clock(other_ops_33_clock),
    .reset(other_ops_33_reset),
    .valid_up(other_ops_33_valid_up),
    .valid_down(other_ops_33_valid_down),
    .I(other_ops_33_I),
    .O(other_ops_33_O)
  );
  Module_0 other_ops_34 ( // @[MapS.scala 10:86]
    .clock(other_ops_34_clock),
    .reset(other_ops_34_reset),
    .valid_up(other_ops_34_valid_up),
    .valid_down(other_ops_34_valid_down),
    .I(other_ops_34_I),
    .O(other_ops_34_O)
  );
  Module_0 other_ops_35 ( // @[MapS.scala 10:86]
    .clock(other_ops_35_clock),
    .reset(other_ops_35_reset),
    .valid_up(other_ops_35_valid_up),
    .valid_down(other_ops_35_valid_down),
    .I(other_ops_35_I),
    .O(other_ops_35_O)
  );
  Module_0 other_ops_36 ( // @[MapS.scala 10:86]
    .clock(other_ops_36_clock),
    .reset(other_ops_36_reset),
    .valid_up(other_ops_36_valid_up),
    .valid_down(other_ops_36_valid_down),
    .I(other_ops_36_I),
    .O(other_ops_36_O)
  );
  Module_0 other_ops_37 ( // @[MapS.scala 10:86]
    .clock(other_ops_37_clock),
    .reset(other_ops_37_reset),
    .valid_up(other_ops_37_valid_up),
    .valid_down(other_ops_37_valid_down),
    .I(other_ops_37_I),
    .O(other_ops_37_O)
  );
  Module_0 other_ops_38 ( // @[MapS.scala 10:86]
    .clock(other_ops_38_clock),
    .reset(other_ops_38_reset),
    .valid_up(other_ops_38_valid_up),
    .valid_down(other_ops_38_valid_down),
    .I(other_ops_38_I),
    .O(other_ops_38_O)
  );
  Module_0 other_ops_39 ( // @[MapS.scala 10:86]
    .clock(other_ops_39_clock),
    .reset(other_ops_39_reset),
    .valid_up(other_ops_39_valid_up),
    .valid_down(other_ops_39_valid_down),
    .I(other_ops_39_I),
    .O(other_ops_39_O)
  );
  Module_0 other_ops_40 ( // @[MapS.scala 10:86]
    .clock(other_ops_40_clock),
    .reset(other_ops_40_reset),
    .valid_up(other_ops_40_valid_up),
    .valid_down(other_ops_40_valid_down),
    .I(other_ops_40_I),
    .O(other_ops_40_O)
  );
  Module_0 other_ops_41 ( // @[MapS.scala 10:86]
    .clock(other_ops_41_clock),
    .reset(other_ops_41_reset),
    .valid_up(other_ops_41_valid_up),
    .valid_down(other_ops_41_valid_down),
    .I(other_ops_41_I),
    .O(other_ops_41_O)
  );
  Module_0 other_ops_42 ( // @[MapS.scala 10:86]
    .clock(other_ops_42_clock),
    .reset(other_ops_42_reset),
    .valid_up(other_ops_42_valid_up),
    .valid_down(other_ops_42_valid_down),
    .I(other_ops_42_I),
    .O(other_ops_42_O)
  );
  Module_0 other_ops_43 ( // @[MapS.scala 10:86]
    .clock(other_ops_43_clock),
    .reset(other_ops_43_reset),
    .valid_up(other_ops_43_valid_up),
    .valid_down(other_ops_43_valid_down),
    .I(other_ops_43_I),
    .O(other_ops_43_O)
  );
  Module_0 other_ops_44 ( // @[MapS.scala 10:86]
    .clock(other_ops_44_clock),
    .reset(other_ops_44_reset),
    .valid_up(other_ops_44_valid_up),
    .valid_down(other_ops_44_valid_down),
    .I(other_ops_44_I),
    .O(other_ops_44_O)
  );
  Module_0 other_ops_45 ( // @[MapS.scala 10:86]
    .clock(other_ops_45_clock),
    .reset(other_ops_45_reset),
    .valid_up(other_ops_45_valid_up),
    .valid_down(other_ops_45_valid_down),
    .I(other_ops_45_I),
    .O(other_ops_45_O)
  );
  Module_0 other_ops_46 ( // @[MapS.scala 10:86]
    .clock(other_ops_46_clock),
    .reset(other_ops_46_reset),
    .valid_up(other_ops_46_valid_up),
    .valid_down(other_ops_46_valid_down),
    .I(other_ops_46_I),
    .O(other_ops_46_O)
  );
  Module_0 other_ops_47 ( // @[MapS.scala 10:86]
    .clock(other_ops_47_clock),
    .reset(other_ops_47_reset),
    .valid_up(other_ops_47_valid_up),
    .valid_down(other_ops_47_valid_down),
    .I(other_ops_47_I),
    .O(other_ops_47_O)
  );
  Module_0 other_ops_48 ( // @[MapS.scala 10:86]
    .clock(other_ops_48_clock),
    .reset(other_ops_48_reset),
    .valid_up(other_ops_48_valid_up),
    .valid_down(other_ops_48_valid_down),
    .I(other_ops_48_I),
    .O(other_ops_48_O)
  );
  Module_0 other_ops_49 ( // @[MapS.scala 10:86]
    .clock(other_ops_49_clock),
    .reset(other_ops_49_reset),
    .valid_up(other_ops_49_valid_up),
    .valid_down(other_ops_49_valid_down),
    .I(other_ops_49_I),
    .O(other_ops_49_O)
  );
  Module_0 other_ops_50 ( // @[MapS.scala 10:86]
    .clock(other_ops_50_clock),
    .reset(other_ops_50_reset),
    .valid_up(other_ops_50_valid_up),
    .valid_down(other_ops_50_valid_down),
    .I(other_ops_50_I),
    .O(other_ops_50_O)
  );
  Module_0 other_ops_51 ( // @[MapS.scala 10:86]
    .clock(other_ops_51_clock),
    .reset(other_ops_51_reset),
    .valid_up(other_ops_51_valid_up),
    .valid_down(other_ops_51_valid_down),
    .I(other_ops_51_I),
    .O(other_ops_51_O)
  );
  Module_0 other_ops_52 ( // @[MapS.scala 10:86]
    .clock(other_ops_52_clock),
    .reset(other_ops_52_reset),
    .valid_up(other_ops_52_valid_up),
    .valid_down(other_ops_52_valid_down),
    .I(other_ops_52_I),
    .O(other_ops_52_O)
  );
  Module_0 other_ops_53 ( // @[MapS.scala 10:86]
    .clock(other_ops_53_clock),
    .reset(other_ops_53_reset),
    .valid_up(other_ops_53_valid_up),
    .valid_down(other_ops_53_valid_down),
    .I(other_ops_53_I),
    .O(other_ops_53_O)
  );
  Module_0 other_ops_54 ( // @[MapS.scala 10:86]
    .clock(other_ops_54_clock),
    .reset(other_ops_54_reset),
    .valid_up(other_ops_54_valid_up),
    .valid_down(other_ops_54_valid_down),
    .I(other_ops_54_I),
    .O(other_ops_54_O)
  );
  Module_0 other_ops_55 ( // @[MapS.scala 10:86]
    .clock(other_ops_55_clock),
    .reset(other_ops_55_reset),
    .valid_up(other_ops_55_valid_up),
    .valid_down(other_ops_55_valid_down),
    .I(other_ops_55_I),
    .O(other_ops_55_O)
  );
  Module_0 other_ops_56 ( // @[MapS.scala 10:86]
    .clock(other_ops_56_clock),
    .reset(other_ops_56_reset),
    .valid_up(other_ops_56_valid_up),
    .valid_down(other_ops_56_valid_down),
    .I(other_ops_56_I),
    .O(other_ops_56_O)
  );
  Module_0 other_ops_57 ( // @[MapS.scala 10:86]
    .clock(other_ops_57_clock),
    .reset(other_ops_57_reset),
    .valid_up(other_ops_57_valid_up),
    .valid_down(other_ops_57_valid_down),
    .I(other_ops_57_I),
    .O(other_ops_57_O)
  );
  Module_0 other_ops_58 ( // @[MapS.scala 10:86]
    .clock(other_ops_58_clock),
    .reset(other_ops_58_reset),
    .valid_up(other_ops_58_valid_up),
    .valid_down(other_ops_58_valid_down),
    .I(other_ops_58_I),
    .O(other_ops_58_O)
  );
  Module_0 other_ops_59 ( // @[MapS.scala 10:86]
    .clock(other_ops_59_clock),
    .reset(other_ops_59_reset),
    .valid_up(other_ops_59_valid_up),
    .valid_down(other_ops_59_valid_down),
    .I(other_ops_59_I),
    .O(other_ops_59_O)
  );
  Module_0 other_ops_60 ( // @[MapS.scala 10:86]
    .clock(other_ops_60_clock),
    .reset(other_ops_60_reset),
    .valid_up(other_ops_60_valid_up),
    .valid_down(other_ops_60_valid_down),
    .I(other_ops_60_I),
    .O(other_ops_60_O)
  );
  Module_0 other_ops_61 ( // @[MapS.scala 10:86]
    .clock(other_ops_61_clock),
    .reset(other_ops_61_reset),
    .valid_up(other_ops_61_valid_up),
    .valid_down(other_ops_61_valid_down),
    .I(other_ops_61_I),
    .O(other_ops_61_O)
  );
  Module_0 other_ops_62 ( // @[MapS.scala 10:86]
    .clock(other_ops_62_clock),
    .reset(other_ops_62_reset),
    .valid_up(other_ops_62_valid_up),
    .valid_down(other_ops_62_valid_down),
    .I(other_ops_62_I),
    .O(other_ops_62_O)
  );
  Module_0 other_ops_63 ( // @[MapS.scala 10:86]
    .clock(other_ops_63_clock),
    .reset(other_ops_63_reset),
    .valid_up(other_ops_63_valid_up),
    .valid_down(other_ops_63_valid_down),
    .I(other_ops_63_I),
    .O(other_ops_63_O)
  );
  Module_0 other_ops_64 ( // @[MapS.scala 10:86]
    .clock(other_ops_64_clock),
    .reset(other_ops_64_reset),
    .valid_up(other_ops_64_valid_up),
    .valid_down(other_ops_64_valid_down),
    .I(other_ops_64_I),
    .O(other_ops_64_O)
  );
  Module_0 other_ops_65 ( // @[MapS.scala 10:86]
    .clock(other_ops_65_clock),
    .reset(other_ops_65_reset),
    .valid_up(other_ops_65_valid_up),
    .valid_down(other_ops_65_valid_down),
    .I(other_ops_65_I),
    .O(other_ops_65_O)
  );
  Module_0 other_ops_66 ( // @[MapS.scala 10:86]
    .clock(other_ops_66_clock),
    .reset(other_ops_66_reset),
    .valid_up(other_ops_66_valid_up),
    .valid_down(other_ops_66_valid_down),
    .I(other_ops_66_I),
    .O(other_ops_66_O)
  );
  Module_0 other_ops_67 ( // @[MapS.scala 10:86]
    .clock(other_ops_67_clock),
    .reset(other_ops_67_reset),
    .valid_up(other_ops_67_valid_up),
    .valid_down(other_ops_67_valid_down),
    .I(other_ops_67_I),
    .O(other_ops_67_O)
  );
  Module_0 other_ops_68 ( // @[MapS.scala 10:86]
    .clock(other_ops_68_clock),
    .reset(other_ops_68_reset),
    .valid_up(other_ops_68_valid_up),
    .valid_down(other_ops_68_valid_down),
    .I(other_ops_68_I),
    .O(other_ops_68_O)
  );
  Module_0 other_ops_69 ( // @[MapS.scala 10:86]
    .clock(other_ops_69_clock),
    .reset(other_ops_69_reset),
    .valid_up(other_ops_69_valid_up),
    .valid_down(other_ops_69_valid_down),
    .I(other_ops_69_I),
    .O(other_ops_69_O)
  );
  Module_0 other_ops_70 ( // @[MapS.scala 10:86]
    .clock(other_ops_70_clock),
    .reset(other_ops_70_reset),
    .valid_up(other_ops_70_valid_up),
    .valid_down(other_ops_70_valid_down),
    .I(other_ops_70_I),
    .O(other_ops_70_O)
  );
  Module_0 other_ops_71 ( // @[MapS.scala 10:86]
    .clock(other_ops_71_clock),
    .reset(other_ops_71_reset),
    .valid_up(other_ops_71_valid_up),
    .valid_down(other_ops_71_valid_down),
    .I(other_ops_71_I),
    .O(other_ops_71_O)
  );
  Module_0 other_ops_72 ( // @[MapS.scala 10:86]
    .clock(other_ops_72_clock),
    .reset(other_ops_72_reset),
    .valid_up(other_ops_72_valid_up),
    .valid_down(other_ops_72_valid_down),
    .I(other_ops_72_I),
    .O(other_ops_72_O)
  );
  Module_0 other_ops_73 ( // @[MapS.scala 10:86]
    .clock(other_ops_73_clock),
    .reset(other_ops_73_reset),
    .valid_up(other_ops_73_valid_up),
    .valid_down(other_ops_73_valid_down),
    .I(other_ops_73_I),
    .O(other_ops_73_O)
  );
  Module_0 other_ops_74 ( // @[MapS.scala 10:86]
    .clock(other_ops_74_clock),
    .reset(other_ops_74_reset),
    .valid_up(other_ops_74_valid_up),
    .valid_down(other_ops_74_valid_down),
    .I(other_ops_74_I),
    .O(other_ops_74_O)
  );
  Module_0 other_ops_75 ( // @[MapS.scala 10:86]
    .clock(other_ops_75_clock),
    .reset(other_ops_75_reset),
    .valid_up(other_ops_75_valid_up),
    .valid_down(other_ops_75_valid_down),
    .I(other_ops_75_I),
    .O(other_ops_75_O)
  );
  Module_0 other_ops_76 ( // @[MapS.scala 10:86]
    .clock(other_ops_76_clock),
    .reset(other_ops_76_reset),
    .valid_up(other_ops_76_valid_up),
    .valid_down(other_ops_76_valid_down),
    .I(other_ops_76_I),
    .O(other_ops_76_O)
  );
  Module_0 other_ops_77 ( // @[MapS.scala 10:86]
    .clock(other_ops_77_clock),
    .reset(other_ops_77_reset),
    .valid_up(other_ops_77_valid_up),
    .valid_down(other_ops_77_valid_down),
    .I(other_ops_77_I),
    .O(other_ops_77_O)
  );
  Module_0 other_ops_78 ( // @[MapS.scala 10:86]
    .clock(other_ops_78_clock),
    .reset(other_ops_78_reset),
    .valid_up(other_ops_78_valid_up),
    .valid_down(other_ops_78_valid_down),
    .I(other_ops_78_I),
    .O(other_ops_78_O)
  );
  Module_0 other_ops_79 ( // @[MapS.scala 10:86]
    .clock(other_ops_79_clock),
    .reset(other_ops_79_reset),
    .valid_up(other_ops_79_valid_up),
    .valid_down(other_ops_79_valid_down),
    .I(other_ops_79_I),
    .O(other_ops_79_O)
  );
  Module_0 other_ops_80 ( // @[MapS.scala 10:86]
    .clock(other_ops_80_clock),
    .reset(other_ops_80_reset),
    .valid_up(other_ops_80_valid_up),
    .valid_down(other_ops_80_valid_down),
    .I(other_ops_80_I),
    .O(other_ops_80_O)
  );
  Module_0 other_ops_81 ( // @[MapS.scala 10:86]
    .clock(other_ops_81_clock),
    .reset(other_ops_81_reset),
    .valid_up(other_ops_81_valid_up),
    .valid_down(other_ops_81_valid_down),
    .I(other_ops_81_I),
    .O(other_ops_81_O)
  );
  Module_0 other_ops_82 ( // @[MapS.scala 10:86]
    .clock(other_ops_82_clock),
    .reset(other_ops_82_reset),
    .valid_up(other_ops_82_valid_up),
    .valid_down(other_ops_82_valid_down),
    .I(other_ops_82_I),
    .O(other_ops_82_O)
  );
  Module_0 other_ops_83 ( // @[MapS.scala 10:86]
    .clock(other_ops_83_clock),
    .reset(other_ops_83_reset),
    .valid_up(other_ops_83_valid_up),
    .valid_down(other_ops_83_valid_down),
    .I(other_ops_83_I),
    .O(other_ops_83_O)
  );
  Module_0 other_ops_84 ( // @[MapS.scala 10:86]
    .clock(other_ops_84_clock),
    .reset(other_ops_84_reset),
    .valid_up(other_ops_84_valid_up),
    .valid_down(other_ops_84_valid_down),
    .I(other_ops_84_I),
    .O(other_ops_84_O)
  );
  Module_0 other_ops_85 ( // @[MapS.scala 10:86]
    .clock(other_ops_85_clock),
    .reset(other_ops_85_reset),
    .valid_up(other_ops_85_valid_up),
    .valid_down(other_ops_85_valid_down),
    .I(other_ops_85_I),
    .O(other_ops_85_O)
  );
  Module_0 other_ops_86 ( // @[MapS.scala 10:86]
    .clock(other_ops_86_clock),
    .reset(other_ops_86_reset),
    .valid_up(other_ops_86_valid_up),
    .valid_down(other_ops_86_valid_down),
    .I(other_ops_86_I),
    .O(other_ops_86_O)
  );
  Module_0 other_ops_87 ( // @[MapS.scala 10:86]
    .clock(other_ops_87_clock),
    .reset(other_ops_87_reset),
    .valid_up(other_ops_87_valid_up),
    .valid_down(other_ops_87_valid_down),
    .I(other_ops_87_I),
    .O(other_ops_87_O)
  );
  Module_0 other_ops_88 ( // @[MapS.scala 10:86]
    .clock(other_ops_88_clock),
    .reset(other_ops_88_reset),
    .valid_up(other_ops_88_valid_up),
    .valid_down(other_ops_88_valid_down),
    .I(other_ops_88_I),
    .O(other_ops_88_O)
  );
  Module_0 other_ops_89 ( // @[MapS.scala 10:86]
    .clock(other_ops_89_clock),
    .reset(other_ops_89_reset),
    .valid_up(other_ops_89_valid_up),
    .valid_down(other_ops_89_valid_down),
    .I(other_ops_89_I),
    .O(other_ops_89_O)
  );
  Module_0 other_ops_90 ( // @[MapS.scala 10:86]
    .clock(other_ops_90_clock),
    .reset(other_ops_90_reset),
    .valid_up(other_ops_90_valid_up),
    .valid_down(other_ops_90_valid_down),
    .I(other_ops_90_I),
    .O(other_ops_90_O)
  );
  Module_0 other_ops_91 ( // @[MapS.scala 10:86]
    .clock(other_ops_91_clock),
    .reset(other_ops_91_reset),
    .valid_up(other_ops_91_valid_up),
    .valid_down(other_ops_91_valid_down),
    .I(other_ops_91_I),
    .O(other_ops_91_O)
  );
  Module_0 other_ops_92 ( // @[MapS.scala 10:86]
    .clock(other_ops_92_clock),
    .reset(other_ops_92_reset),
    .valid_up(other_ops_92_valid_up),
    .valid_down(other_ops_92_valid_down),
    .I(other_ops_92_I),
    .O(other_ops_92_O)
  );
  Module_0 other_ops_93 ( // @[MapS.scala 10:86]
    .clock(other_ops_93_clock),
    .reset(other_ops_93_reset),
    .valid_up(other_ops_93_valid_up),
    .valid_down(other_ops_93_valid_down),
    .I(other_ops_93_I),
    .O(other_ops_93_O)
  );
  Module_0 other_ops_94 ( // @[MapS.scala 10:86]
    .clock(other_ops_94_clock),
    .reset(other_ops_94_reset),
    .valid_up(other_ops_94_valid_up),
    .valid_down(other_ops_94_valid_down),
    .I(other_ops_94_I),
    .O(other_ops_94_O)
  );
  Module_0 other_ops_95 ( // @[MapS.scala 10:86]
    .clock(other_ops_95_clock),
    .reset(other_ops_95_reset),
    .valid_up(other_ops_95_valid_up),
    .valid_down(other_ops_95_valid_down),
    .I(other_ops_95_I),
    .O(other_ops_95_O)
  );
  Module_0 other_ops_96 ( // @[MapS.scala 10:86]
    .clock(other_ops_96_clock),
    .reset(other_ops_96_reset),
    .valid_up(other_ops_96_valid_up),
    .valid_down(other_ops_96_valid_down),
    .I(other_ops_96_I),
    .O(other_ops_96_O)
  );
  Module_0 other_ops_97 ( // @[MapS.scala 10:86]
    .clock(other_ops_97_clock),
    .reset(other_ops_97_reset),
    .valid_up(other_ops_97_valid_up),
    .valid_down(other_ops_97_valid_down),
    .I(other_ops_97_I),
    .O(other_ops_97_O)
  );
  Module_0 other_ops_98 ( // @[MapS.scala 10:86]
    .clock(other_ops_98_clock),
    .reset(other_ops_98_reset),
    .valid_up(other_ops_98_valid_up),
    .valid_down(other_ops_98_valid_down),
    .I(other_ops_98_I),
    .O(other_ops_98_O)
  );
  Module_0 other_ops_99 ( // @[MapS.scala 10:86]
    .clock(other_ops_99_clock),
    .reset(other_ops_99_reset),
    .valid_up(other_ops_99_valid_up),
    .valid_down(other_ops_99_valid_down),
    .I(other_ops_99_I),
    .O(other_ops_99_O)
  );
  Module_0 other_ops_100 ( // @[MapS.scala 10:86]
    .clock(other_ops_100_clock),
    .reset(other_ops_100_reset),
    .valid_up(other_ops_100_valid_up),
    .valid_down(other_ops_100_valid_down),
    .I(other_ops_100_I),
    .O(other_ops_100_O)
  );
  Module_0 other_ops_101 ( // @[MapS.scala 10:86]
    .clock(other_ops_101_clock),
    .reset(other_ops_101_reset),
    .valid_up(other_ops_101_valid_up),
    .valid_down(other_ops_101_valid_down),
    .I(other_ops_101_I),
    .O(other_ops_101_O)
  );
  Module_0 other_ops_102 ( // @[MapS.scala 10:86]
    .clock(other_ops_102_clock),
    .reset(other_ops_102_reset),
    .valid_up(other_ops_102_valid_up),
    .valid_down(other_ops_102_valid_down),
    .I(other_ops_102_I),
    .O(other_ops_102_O)
  );
  Module_0 other_ops_103 ( // @[MapS.scala 10:86]
    .clock(other_ops_103_clock),
    .reset(other_ops_103_reset),
    .valid_up(other_ops_103_valid_up),
    .valid_down(other_ops_103_valid_down),
    .I(other_ops_103_I),
    .O(other_ops_103_O)
  );
  Module_0 other_ops_104 ( // @[MapS.scala 10:86]
    .clock(other_ops_104_clock),
    .reset(other_ops_104_reset),
    .valid_up(other_ops_104_valid_up),
    .valid_down(other_ops_104_valid_down),
    .I(other_ops_104_I),
    .O(other_ops_104_O)
  );
  Module_0 other_ops_105 ( // @[MapS.scala 10:86]
    .clock(other_ops_105_clock),
    .reset(other_ops_105_reset),
    .valid_up(other_ops_105_valid_up),
    .valid_down(other_ops_105_valid_down),
    .I(other_ops_105_I),
    .O(other_ops_105_O)
  );
  Module_0 other_ops_106 ( // @[MapS.scala 10:86]
    .clock(other_ops_106_clock),
    .reset(other_ops_106_reset),
    .valid_up(other_ops_106_valid_up),
    .valid_down(other_ops_106_valid_down),
    .I(other_ops_106_I),
    .O(other_ops_106_O)
  );
  Module_0 other_ops_107 ( // @[MapS.scala 10:86]
    .clock(other_ops_107_clock),
    .reset(other_ops_107_reset),
    .valid_up(other_ops_107_valid_up),
    .valid_down(other_ops_107_valid_down),
    .I(other_ops_107_I),
    .O(other_ops_107_O)
  );
  Module_0 other_ops_108 ( // @[MapS.scala 10:86]
    .clock(other_ops_108_clock),
    .reset(other_ops_108_reset),
    .valid_up(other_ops_108_valid_up),
    .valid_down(other_ops_108_valid_down),
    .I(other_ops_108_I),
    .O(other_ops_108_O)
  );
  Module_0 other_ops_109 ( // @[MapS.scala 10:86]
    .clock(other_ops_109_clock),
    .reset(other_ops_109_reset),
    .valid_up(other_ops_109_valid_up),
    .valid_down(other_ops_109_valid_down),
    .I(other_ops_109_I),
    .O(other_ops_109_O)
  );
  Module_0 other_ops_110 ( // @[MapS.scala 10:86]
    .clock(other_ops_110_clock),
    .reset(other_ops_110_reset),
    .valid_up(other_ops_110_valid_up),
    .valid_down(other_ops_110_valid_down),
    .I(other_ops_110_I),
    .O(other_ops_110_O)
  );
  Module_0 other_ops_111 ( // @[MapS.scala 10:86]
    .clock(other_ops_111_clock),
    .reset(other_ops_111_reset),
    .valid_up(other_ops_111_valid_up),
    .valid_down(other_ops_111_valid_down),
    .I(other_ops_111_I),
    .O(other_ops_111_O)
  );
  Module_0 other_ops_112 ( // @[MapS.scala 10:86]
    .clock(other_ops_112_clock),
    .reset(other_ops_112_reset),
    .valid_up(other_ops_112_valid_up),
    .valid_down(other_ops_112_valid_down),
    .I(other_ops_112_I),
    .O(other_ops_112_O)
  );
  Module_0 other_ops_113 ( // @[MapS.scala 10:86]
    .clock(other_ops_113_clock),
    .reset(other_ops_113_reset),
    .valid_up(other_ops_113_valid_up),
    .valid_down(other_ops_113_valid_down),
    .I(other_ops_113_I),
    .O(other_ops_113_O)
  );
  Module_0 other_ops_114 ( // @[MapS.scala 10:86]
    .clock(other_ops_114_clock),
    .reset(other_ops_114_reset),
    .valid_up(other_ops_114_valid_up),
    .valid_down(other_ops_114_valid_down),
    .I(other_ops_114_I),
    .O(other_ops_114_O)
  );
  Module_0 other_ops_115 ( // @[MapS.scala 10:86]
    .clock(other_ops_115_clock),
    .reset(other_ops_115_reset),
    .valid_up(other_ops_115_valid_up),
    .valid_down(other_ops_115_valid_down),
    .I(other_ops_115_I),
    .O(other_ops_115_O)
  );
  Module_0 other_ops_116 ( // @[MapS.scala 10:86]
    .clock(other_ops_116_clock),
    .reset(other_ops_116_reset),
    .valid_up(other_ops_116_valid_up),
    .valid_down(other_ops_116_valid_down),
    .I(other_ops_116_I),
    .O(other_ops_116_O)
  );
  Module_0 other_ops_117 ( // @[MapS.scala 10:86]
    .clock(other_ops_117_clock),
    .reset(other_ops_117_reset),
    .valid_up(other_ops_117_valid_up),
    .valid_down(other_ops_117_valid_down),
    .I(other_ops_117_I),
    .O(other_ops_117_O)
  );
  Module_0 other_ops_118 ( // @[MapS.scala 10:86]
    .clock(other_ops_118_clock),
    .reset(other_ops_118_reset),
    .valid_up(other_ops_118_valid_up),
    .valid_down(other_ops_118_valid_down),
    .I(other_ops_118_I),
    .O(other_ops_118_O)
  );
  Module_0 other_ops_119 ( // @[MapS.scala 10:86]
    .clock(other_ops_119_clock),
    .reset(other_ops_119_reset),
    .valid_up(other_ops_119_valid_up),
    .valid_down(other_ops_119_valid_down),
    .I(other_ops_119_I),
    .O(other_ops_119_O)
  );
  Module_0 other_ops_120 ( // @[MapS.scala 10:86]
    .clock(other_ops_120_clock),
    .reset(other_ops_120_reset),
    .valid_up(other_ops_120_valid_up),
    .valid_down(other_ops_120_valid_down),
    .I(other_ops_120_I),
    .O(other_ops_120_O)
  );
  Module_0 other_ops_121 ( // @[MapS.scala 10:86]
    .clock(other_ops_121_clock),
    .reset(other_ops_121_reset),
    .valid_up(other_ops_121_valid_up),
    .valid_down(other_ops_121_valid_down),
    .I(other_ops_121_I),
    .O(other_ops_121_O)
  );
  Module_0 other_ops_122 ( // @[MapS.scala 10:86]
    .clock(other_ops_122_clock),
    .reset(other_ops_122_reset),
    .valid_up(other_ops_122_valid_up),
    .valid_down(other_ops_122_valid_down),
    .I(other_ops_122_I),
    .O(other_ops_122_O)
  );
  Module_0 other_ops_123 ( // @[MapS.scala 10:86]
    .clock(other_ops_123_clock),
    .reset(other_ops_123_reset),
    .valid_up(other_ops_123_valid_up),
    .valid_down(other_ops_123_valid_down),
    .I(other_ops_123_I),
    .O(other_ops_123_O)
  );
  Module_0 other_ops_124 ( // @[MapS.scala 10:86]
    .clock(other_ops_124_clock),
    .reset(other_ops_124_reset),
    .valid_up(other_ops_124_valid_up),
    .valid_down(other_ops_124_valid_down),
    .I(other_ops_124_I),
    .O(other_ops_124_O)
  );
  Module_0 other_ops_125 ( // @[MapS.scala 10:86]
    .clock(other_ops_125_clock),
    .reset(other_ops_125_reset),
    .valid_up(other_ops_125_valid_up),
    .valid_down(other_ops_125_valid_down),
    .I(other_ops_125_I),
    .O(other_ops_125_O)
  );
  Module_0 other_ops_126 ( // @[MapS.scala 10:86]
    .clock(other_ops_126_clock),
    .reset(other_ops_126_reset),
    .valid_up(other_ops_126_valid_up),
    .valid_down(other_ops_126_valid_down),
    .I(other_ops_126_I),
    .O(other_ops_126_O)
  );
  Module_0 other_ops_127 ( // @[MapS.scala 10:86]
    .clock(other_ops_127_clock),
    .reset(other_ops_127_reset),
    .valid_up(other_ops_127_valid_up),
    .valid_down(other_ops_127_valid_down),
    .I(other_ops_127_I),
    .O(other_ops_127_O)
  );
  Module_0 other_ops_128 ( // @[MapS.scala 10:86]
    .clock(other_ops_128_clock),
    .reset(other_ops_128_reset),
    .valid_up(other_ops_128_valid_up),
    .valid_down(other_ops_128_valid_down),
    .I(other_ops_128_I),
    .O(other_ops_128_O)
  );
  Module_0 other_ops_129 ( // @[MapS.scala 10:86]
    .clock(other_ops_129_clock),
    .reset(other_ops_129_reset),
    .valid_up(other_ops_129_valid_up),
    .valid_down(other_ops_129_valid_down),
    .I(other_ops_129_I),
    .O(other_ops_129_O)
  );
  Module_0 other_ops_130 ( // @[MapS.scala 10:86]
    .clock(other_ops_130_clock),
    .reset(other_ops_130_reset),
    .valid_up(other_ops_130_valid_up),
    .valid_down(other_ops_130_valid_down),
    .I(other_ops_130_I),
    .O(other_ops_130_O)
  );
  Module_0 other_ops_131 ( // @[MapS.scala 10:86]
    .clock(other_ops_131_clock),
    .reset(other_ops_131_reset),
    .valid_up(other_ops_131_valid_up),
    .valid_down(other_ops_131_valid_down),
    .I(other_ops_131_I),
    .O(other_ops_131_O)
  );
  Module_0 other_ops_132 ( // @[MapS.scala 10:86]
    .clock(other_ops_132_clock),
    .reset(other_ops_132_reset),
    .valid_up(other_ops_132_valid_up),
    .valid_down(other_ops_132_valid_down),
    .I(other_ops_132_I),
    .O(other_ops_132_O)
  );
  Module_0 other_ops_133 ( // @[MapS.scala 10:86]
    .clock(other_ops_133_clock),
    .reset(other_ops_133_reset),
    .valid_up(other_ops_133_valid_up),
    .valid_down(other_ops_133_valid_down),
    .I(other_ops_133_I),
    .O(other_ops_133_O)
  );
  Module_0 other_ops_134 ( // @[MapS.scala 10:86]
    .clock(other_ops_134_clock),
    .reset(other_ops_134_reset),
    .valid_up(other_ops_134_valid_up),
    .valid_down(other_ops_134_valid_down),
    .I(other_ops_134_I),
    .O(other_ops_134_O)
  );
  Module_0 other_ops_135 ( // @[MapS.scala 10:86]
    .clock(other_ops_135_clock),
    .reset(other_ops_135_reset),
    .valid_up(other_ops_135_valid_up),
    .valid_down(other_ops_135_valid_down),
    .I(other_ops_135_I),
    .O(other_ops_135_O)
  );
  Module_0 other_ops_136 ( // @[MapS.scala 10:86]
    .clock(other_ops_136_clock),
    .reset(other_ops_136_reset),
    .valid_up(other_ops_136_valid_up),
    .valid_down(other_ops_136_valid_down),
    .I(other_ops_136_I),
    .O(other_ops_136_O)
  );
  Module_0 other_ops_137 ( // @[MapS.scala 10:86]
    .clock(other_ops_137_clock),
    .reset(other_ops_137_reset),
    .valid_up(other_ops_137_valid_up),
    .valid_down(other_ops_137_valid_down),
    .I(other_ops_137_I),
    .O(other_ops_137_O)
  );
  Module_0 other_ops_138 ( // @[MapS.scala 10:86]
    .clock(other_ops_138_clock),
    .reset(other_ops_138_reset),
    .valid_up(other_ops_138_valid_up),
    .valid_down(other_ops_138_valid_down),
    .I(other_ops_138_I),
    .O(other_ops_138_O)
  );
  Module_0 other_ops_139 ( // @[MapS.scala 10:86]
    .clock(other_ops_139_clock),
    .reset(other_ops_139_reset),
    .valid_up(other_ops_139_valid_up),
    .valid_down(other_ops_139_valid_down),
    .I(other_ops_139_I),
    .O(other_ops_139_O)
  );
  Module_0 other_ops_140 ( // @[MapS.scala 10:86]
    .clock(other_ops_140_clock),
    .reset(other_ops_140_reset),
    .valid_up(other_ops_140_valid_up),
    .valid_down(other_ops_140_valid_down),
    .I(other_ops_140_I),
    .O(other_ops_140_O)
  );
  Module_0 other_ops_141 ( // @[MapS.scala 10:86]
    .clock(other_ops_141_clock),
    .reset(other_ops_141_reset),
    .valid_up(other_ops_141_valid_up),
    .valid_down(other_ops_141_valid_down),
    .I(other_ops_141_I),
    .O(other_ops_141_O)
  );
  Module_0 other_ops_142 ( // @[MapS.scala 10:86]
    .clock(other_ops_142_clock),
    .reset(other_ops_142_reset),
    .valid_up(other_ops_142_valid_up),
    .valid_down(other_ops_142_valid_down),
    .I(other_ops_142_I),
    .O(other_ops_142_O)
  );
  Module_0 other_ops_143 ( // @[MapS.scala 10:86]
    .clock(other_ops_143_clock),
    .reset(other_ops_143_reset),
    .valid_up(other_ops_143_valid_up),
    .valid_down(other_ops_143_valid_down),
    .I(other_ops_143_I),
    .O(other_ops_143_O)
  );
  Module_0 other_ops_144 ( // @[MapS.scala 10:86]
    .clock(other_ops_144_clock),
    .reset(other_ops_144_reset),
    .valid_up(other_ops_144_valid_up),
    .valid_down(other_ops_144_valid_down),
    .I(other_ops_144_I),
    .O(other_ops_144_O)
  );
  Module_0 other_ops_145 ( // @[MapS.scala 10:86]
    .clock(other_ops_145_clock),
    .reset(other_ops_145_reset),
    .valid_up(other_ops_145_valid_up),
    .valid_down(other_ops_145_valid_down),
    .I(other_ops_145_I),
    .O(other_ops_145_O)
  );
  Module_0 other_ops_146 ( // @[MapS.scala 10:86]
    .clock(other_ops_146_clock),
    .reset(other_ops_146_reset),
    .valid_up(other_ops_146_valid_up),
    .valid_down(other_ops_146_valid_down),
    .I(other_ops_146_I),
    .O(other_ops_146_O)
  );
  Module_0 other_ops_147 ( // @[MapS.scala 10:86]
    .clock(other_ops_147_clock),
    .reset(other_ops_147_reset),
    .valid_up(other_ops_147_valid_up),
    .valid_down(other_ops_147_valid_down),
    .I(other_ops_147_I),
    .O(other_ops_147_O)
  );
  Module_0 other_ops_148 ( // @[MapS.scala 10:86]
    .clock(other_ops_148_clock),
    .reset(other_ops_148_reset),
    .valid_up(other_ops_148_valid_up),
    .valid_down(other_ops_148_valid_down),
    .I(other_ops_148_I),
    .O(other_ops_148_O)
  );
  Module_0 other_ops_149 ( // @[MapS.scala 10:86]
    .clock(other_ops_149_clock),
    .reset(other_ops_149_reset),
    .valid_up(other_ops_149_valid_up),
    .valid_down(other_ops_149_valid_down),
    .I(other_ops_149_I),
    .O(other_ops_149_O)
  );
  Module_0 other_ops_150 ( // @[MapS.scala 10:86]
    .clock(other_ops_150_clock),
    .reset(other_ops_150_reset),
    .valid_up(other_ops_150_valid_up),
    .valid_down(other_ops_150_valid_down),
    .I(other_ops_150_I),
    .O(other_ops_150_O)
  );
  Module_0 other_ops_151 ( // @[MapS.scala 10:86]
    .clock(other_ops_151_clock),
    .reset(other_ops_151_reset),
    .valid_up(other_ops_151_valid_up),
    .valid_down(other_ops_151_valid_down),
    .I(other_ops_151_I),
    .O(other_ops_151_O)
  );
  Module_0 other_ops_152 ( // @[MapS.scala 10:86]
    .clock(other_ops_152_clock),
    .reset(other_ops_152_reset),
    .valid_up(other_ops_152_valid_up),
    .valid_down(other_ops_152_valid_down),
    .I(other_ops_152_I),
    .O(other_ops_152_O)
  );
  Module_0 other_ops_153 ( // @[MapS.scala 10:86]
    .clock(other_ops_153_clock),
    .reset(other_ops_153_reset),
    .valid_up(other_ops_153_valid_up),
    .valid_down(other_ops_153_valid_down),
    .I(other_ops_153_I),
    .O(other_ops_153_O)
  );
  Module_0 other_ops_154 ( // @[MapS.scala 10:86]
    .clock(other_ops_154_clock),
    .reset(other_ops_154_reset),
    .valid_up(other_ops_154_valid_up),
    .valid_down(other_ops_154_valid_down),
    .I(other_ops_154_I),
    .O(other_ops_154_O)
  );
  Module_0 other_ops_155 ( // @[MapS.scala 10:86]
    .clock(other_ops_155_clock),
    .reset(other_ops_155_reset),
    .valid_up(other_ops_155_valid_up),
    .valid_down(other_ops_155_valid_down),
    .I(other_ops_155_I),
    .O(other_ops_155_O)
  );
  Module_0 other_ops_156 ( // @[MapS.scala 10:86]
    .clock(other_ops_156_clock),
    .reset(other_ops_156_reset),
    .valid_up(other_ops_156_valid_up),
    .valid_down(other_ops_156_valid_down),
    .I(other_ops_156_I),
    .O(other_ops_156_O)
  );
  Module_0 other_ops_157 ( // @[MapS.scala 10:86]
    .clock(other_ops_157_clock),
    .reset(other_ops_157_reset),
    .valid_up(other_ops_157_valid_up),
    .valid_down(other_ops_157_valid_down),
    .I(other_ops_157_I),
    .O(other_ops_157_O)
  );
  Module_0 other_ops_158 ( // @[MapS.scala 10:86]
    .clock(other_ops_158_clock),
    .reset(other_ops_158_reset),
    .valid_up(other_ops_158_valid_up),
    .valid_down(other_ops_158_valid_down),
    .I(other_ops_158_I),
    .O(other_ops_158_O)
  );
  Module_0 other_ops_159 ( // @[MapS.scala 10:86]
    .clock(other_ops_159_clock),
    .reset(other_ops_159_reset),
    .valid_up(other_ops_159_valid_up),
    .valid_down(other_ops_159_valid_down),
    .I(other_ops_159_I),
    .O(other_ops_159_O)
  );
  Module_0 other_ops_160 ( // @[MapS.scala 10:86]
    .clock(other_ops_160_clock),
    .reset(other_ops_160_reset),
    .valid_up(other_ops_160_valid_up),
    .valid_down(other_ops_160_valid_down),
    .I(other_ops_160_I),
    .O(other_ops_160_O)
  );
  Module_0 other_ops_161 ( // @[MapS.scala 10:86]
    .clock(other_ops_161_clock),
    .reset(other_ops_161_reset),
    .valid_up(other_ops_161_valid_up),
    .valid_down(other_ops_161_valid_down),
    .I(other_ops_161_I),
    .O(other_ops_161_O)
  );
  Module_0 other_ops_162 ( // @[MapS.scala 10:86]
    .clock(other_ops_162_clock),
    .reset(other_ops_162_reset),
    .valid_up(other_ops_162_valid_up),
    .valid_down(other_ops_162_valid_down),
    .I(other_ops_162_I),
    .O(other_ops_162_O)
  );
  Module_0 other_ops_163 ( // @[MapS.scala 10:86]
    .clock(other_ops_163_clock),
    .reset(other_ops_163_reset),
    .valid_up(other_ops_163_valid_up),
    .valid_down(other_ops_163_valid_down),
    .I(other_ops_163_I),
    .O(other_ops_163_O)
  );
  Module_0 other_ops_164 ( // @[MapS.scala 10:86]
    .clock(other_ops_164_clock),
    .reset(other_ops_164_reset),
    .valid_up(other_ops_164_valid_up),
    .valid_down(other_ops_164_valid_down),
    .I(other_ops_164_I),
    .O(other_ops_164_O)
  );
  Module_0 other_ops_165 ( // @[MapS.scala 10:86]
    .clock(other_ops_165_clock),
    .reset(other_ops_165_reset),
    .valid_up(other_ops_165_valid_up),
    .valid_down(other_ops_165_valid_down),
    .I(other_ops_165_I),
    .O(other_ops_165_O)
  );
  Module_0 other_ops_166 ( // @[MapS.scala 10:86]
    .clock(other_ops_166_clock),
    .reset(other_ops_166_reset),
    .valid_up(other_ops_166_valid_up),
    .valid_down(other_ops_166_valid_down),
    .I(other_ops_166_I),
    .O(other_ops_166_O)
  );
  Module_0 other_ops_167 ( // @[MapS.scala 10:86]
    .clock(other_ops_167_clock),
    .reset(other_ops_167_reset),
    .valid_up(other_ops_167_valid_up),
    .valid_down(other_ops_167_valid_down),
    .I(other_ops_167_I),
    .O(other_ops_167_O)
  );
  Module_0 other_ops_168 ( // @[MapS.scala 10:86]
    .clock(other_ops_168_clock),
    .reset(other_ops_168_reset),
    .valid_up(other_ops_168_valid_up),
    .valid_down(other_ops_168_valid_down),
    .I(other_ops_168_I),
    .O(other_ops_168_O)
  );
  Module_0 other_ops_169 ( // @[MapS.scala 10:86]
    .clock(other_ops_169_clock),
    .reset(other_ops_169_reset),
    .valid_up(other_ops_169_valid_up),
    .valid_down(other_ops_169_valid_down),
    .I(other_ops_169_I),
    .O(other_ops_169_O)
  );
  Module_0 other_ops_170 ( // @[MapS.scala 10:86]
    .clock(other_ops_170_clock),
    .reset(other_ops_170_reset),
    .valid_up(other_ops_170_valid_up),
    .valid_down(other_ops_170_valid_down),
    .I(other_ops_170_I),
    .O(other_ops_170_O)
  );
  Module_0 other_ops_171 ( // @[MapS.scala 10:86]
    .clock(other_ops_171_clock),
    .reset(other_ops_171_reset),
    .valid_up(other_ops_171_valid_up),
    .valid_down(other_ops_171_valid_down),
    .I(other_ops_171_I),
    .O(other_ops_171_O)
  );
  Module_0 other_ops_172 ( // @[MapS.scala 10:86]
    .clock(other_ops_172_clock),
    .reset(other_ops_172_reset),
    .valid_up(other_ops_172_valid_up),
    .valid_down(other_ops_172_valid_down),
    .I(other_ops_172_I),
    .O(other_ops_172_O)
  );
  Module_0 other_ops_173 ( // @[MapS.scala 10:86]
    .clock(other_ops_173_clock),
    .reset(other_ops_173_reset),
    .valid_up(other_ops_173_valid_up),
    .valid_down(other_ops_173_valid_down),
    .I(other_ops_173_I),
    .O(other_ops_173_O)
  );
  Module_0 other_ops_174 ( // @[MapS.scala 10:86]
    .clock(other_ops_174_clock),
    .reset(other_ops_174_reset),
    .valid_up(other_ops_174_valid_up),
    .valid_down(other_ops_174_valid_down),
    .I(other_ops_174_I),
    .O(other_ops_174_O)
  );
  Module_0 other_ops_175 ( // @[MapS.scala 10:86]
    .clock(other_ops_175_clock),
    .reset(other_ops_175_reset),
    .valid_up(other_ops_175_valid_up),
    .valid_down(other_ops_175_valid_down),
    .I(other_ops_175_I),
    .O(other_ops_175_O)
  );
  Module_0 other_ops_176 ( // @[MapS.scala 10:86]
    .clock(other_ops_176_clock),
    .reset(other_ops_176_reset),
    .valid_up(other_ops_176_valid_up),
    .valid_down(other_ops_176_valid_down),
    .I(other_ops_176_I),
    .O(other_ops_176_O)
  );
  Module_0 other_ops_177 ( // @[MapS.scala 10:86]
    .clock(other_ops_177_clock),
    .reset(other_ops_177_reset),
    .valid_up(other_ops_177_valid_up),
    .valid_down(other_ops_177_valid_down),
    .I(other_ops_177_I),
    .O(other_ops_177_O)
  );
  Module_0 other_ops_178 ( // @[MapS.scala 10:86]
    .clock(other_ops_178_clock),
    .reset(other_ops_178_reset),
    .valid_up(other_ops_178_valid_up),
    .valid_down(other_ops_178_valid_down),
    .I(other_ops_178_I),
    .O(other_ops_178_O)
  );
  Module_0 other_ops_179 ( // @[MapS.scala 10:86]
    .clock(other_ops_179_clock),
    .reset(other_ops_179_reset),
    .valid_up(other_ops_179_valid_up),
    .valid_down(other_ops_179_valid_down),
    .I(other_ops_179_I),
    .O(other_ops_179_O)
  );
  Module_0 other_ops_180 ( // @[MapS.scala 10:86]
    .clock(other_ops_180_clock),
    .reset(other_ops_180_reset),
    .valid_up(other_ops_180_valid_up),
    .valid_down(other_ops_180_valid_down),
    .I(other_ops_180_I),
    .O(other_ops_180_O)
  );
  Module_0 other_ops_181 ( // @[MapS.scala 10:86]
    .clock(other_ops_181_clock),
    .reset(other_ops_181_reset),
    .valid_up(other_ops_181_valid_up),
    .valid_down(other_ops_181_valid_down),
    .I(other_ops_181_I),
    .O(other_ops_181_O)
  );
  Module_0 other_ops_182 ( // @[MapS.scala 10:86]
    .clock(other_ops_182_clock),
    .reset(other_ops_182_reset),
    .valid_up(other_ops_182_valid_up),
    .valid_down(other_ops_182_valid_down),
    .I(other_ops_182_I),
    .O(other_ops_182_O)
  );
  Module_0 other_ops_183 ( // @[MapS.scala 10:86]
    .clock(other_ops_183_clock),
    .reset(other_ops_183_reset),
    .valid_up(other_ops_183_valid_up),
    .valid_down(other_ops_183_valid_down),
    .I(other_ops_183_I),
    .O(other_ops_183_O)
  );
  Module_0 other_ops_184 ( // @[MapS.scala 10:86]
    .clock(other_ops_184_clock),
    .reset(other_ops_184_reset),
    .valid_up(other_ops_184_valid_up),
    .valid_down(other_ops_184_valid_down),
    .I(other_ops_184_I),
    .O(other_ops_184_O)
  );
  Module_0 other_ops_185 ( // @[MapS.scala 10:86]
    .clock(other_ops_185_clock),
    .reset(other_ops_185_reset),
    .valid_up(other_ops_185_valid_up),
    .valid_down(other_ops_185_valid_down),
    .I(other_ops_185_I),
    .O(other_ops_185_O)
  );
  Module_0 other_ops_186 ( // @[MapS.scala 10:86]
    .clock(other_ops_186_clock),
    .reset(other_ops_186_reset),
    .valid_up(other_ops_186_valid_up),
    .valid_down(other_ops_186_valid_down),
    .I(other_ops_186_I),
    .O(other_ops_186_O)
  );
  Module_0 other_ops_187 ( // @[MapS.scala 10:86]
    .clock(other_ops_187_clock),
    .reset(other_ops_187_reset),
    .valid_up(other_ops_187_valid_up),
    .valid_down(other_ops_187_valid_down),
    .I(other_ops_187_I),
    .O(other_ops_187_O)
  );
  Module_0 other_ops_188 ( // @[MapS.scala 10:86]
    .clock(other_ops_188_clock),
    .reset(other_ops_188_reset),
    .valid_up(other_ops_188_valid_up),
    .valid_down(other_ops_188_valid_down),
    .I(other_ops_188_I),
    .O(other_ops_188_O)
  );
  Module_0 other_ops_189 ( // @[MapS.scala 10:86]
    .clock(other_ops_189_clock),
    .reset(other_ops_189_reset),
    .valid_up(other_ops_189_valid_up),
    .valid_down(other_ops_189_valid_down),
    .I(other_ops_189_I),
    .O(other_ops_189_O)
  );
  Module_0 other_ops_190 ( // @[MapS.scala 10:86]
    .clock(other_ops_190_clock),
    .reset(other_ops_190_reset),
    .valid_up(other_ops_190_valid_up),
    .valid_down(other_ops_190_valid_down),
    .I(other_ops_190_I),
    .O(other_ops_190_O)
  );
  Module_0 other_ops_191 ( // @[MapS.scala 10:86]
    .clock(other_ops_191_clock),
    .reset(other_ops_191_reset),
    .valid_up(other_ops_191_valid_up),
    .valid_down(other_ops_191_valid_down),
    .I(other_ops_191_I),
    .O(other_ops_191_O)
  );
  Module_0 other_ops_192 ( // @[MapS.scala 10:86]
    .clock(other_ops_192_clock),
    .reset(other_ops_192_reset),
    .valid_up(other_ops_192_valid_up),
    .valid_down(other_ops_192_valid_down),
    .I(other_ops_192_I),
    .O(other_ops_192_O)
  );
  Module_0 other_ops_193 ( // @[MapS.scala 10:86]
    .clock(other_ops_193_clock),
    .reset(other_ops_193_reset),
    .valid_up(other_ops_193_valid_up),
    .valid_down(other_ops_193_valid_down),
    .I(other_ops_193_I),
    .O(other_ops_193_O)
  );
  Module_0 other_ops_194 ( // @[MapS.scala 10:86]
    .clock(other_ops_194_clock),
    .reset(other_ops_194_reset),
    .valid_up(other_ops_194_valid_up),
    .valid_down(other_ops_194_valid_down),
    .I(other_ops_194_I),
    .O(other_ops_194_O)
  );
  Module_0 other_ops_195 ( // @[MapS.scala 10:86]
    .clock(other_ops_195_clock),
    .reset(other_ops_195_reset),
    .valid_up(other_ops_195_valid_up),
    .valid_down(other_ops_195_valid_down),
    .I(other_ops_195_I),
    .O(other_ops_195_O)
  );
  Module_0 other_ops_196 ( // @[MapS.scala 10:86]
    .clock(other_ops_196_clock),
    .reset(other_ops_196_reset),
    .valid_up(other_ops_196_valid_up),
    .valid_down(other_ops_196_valid_down),
    .I(other_ops_196_I),
    .O(other_ops_196_O)
  );
  Module_0 other_ops_197 ( // @[MapS.scala 10:86]
    .clock(other_ops_197_clock),
    .reset(other_ops_197_reset),
    .valid_up(other_ops_197_valid_up),
    .valid_down(other_ops_197_valid_down),
    .I(other_ops_197_I),
    .O(other_ops_197_O)
  );
  Module_0 other_ops_198 ( // @[MapS.scala 10:86]
    .clock(other_ops_198_clock),
    .reset(other_ops_198_reset),
    .valid_up(other_ops_198_valid_up),
    .valid_down(other_ops_198_valid_down),
    .I(other_ops_198_I),
    .O(other_ops_198_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign _T_14 = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:83]
  assign _T_15 = _T_14 & other_ops_15_valid_down; // @[MapS.scala 23:83]
  assign _T_16 = _T_15 & other_ops_16_valid_down; // @[MapS.scala 23:83]
  assign _T_17 = _T_16 & other_ops_17_valid_down; // @[MapS.scala 23:83]
  assign _T_18 = _T_17 & other_ops_18_valid_down; // @[MapS.scala 23:83]
  assign _T_19 = _T_18 & other_ops_19_valid_down; // @[MapS.scala 23:83]
  assign _T_20 = _T_19 & other_ops_20_valid_down; // @[MapS.scala 23:83]
  assign _T_21 = _T_20 & other_ops_21_valid_down; // @[MapS.scala 23:83]
  assign _T_22 = _T_21 & other_ops_22_valid_down; // @[MapS.scala 23:83]
  assign _T_23 = _T_22 & other_ops_23_valid_down; // @[MapS.scala 23:83]
  assign _T_24 = _T_23 & other_ops_24_valid_down; // @[MapS.scala 23:83]
  assign _T_25 = _T_24 & other_ops_25_valid_down; // @[MapS.scala 23:83]
  assign _T_26 = _T_25 & other_ops_26_valid_down; // @[MapS.scala 23:83]
  assign _T_27 = _T_26 & other_ops_27_valid_down; // @[MapS.scala 23:83]
  assign _T_28 = _T_27 & other_ops_28_valid_down; // @[MapS.scala 23:83]
  assign _T_29 = _T_28 & other_ops_29_valid_down; // @[MapS.scala 23:83]
  assign _T_30 = _T_29 & other_ops_30_valid_down; // @[MapS.scala 23:83]
  assign _T_31 = _T_30 & other_ops_31_valid_down; // @[MapS.scala 23:83]
  assign _T_32 = _T_31 & other_ops_32_valid_down; // @[MapS.scala 23:83]
  assign _T_33 = _T_32 & other_ops_33_valid_down; // @[MapS.scala 23:83]
  assign _T_34 = _T_33 & other_ops_34_valid_down; // @[MapS.scala 23:83]
  assign _T_35 = _T_34 & other_ops_35_valid_down; // @[MapS.scala 23:83]
  assign _T_36 = _T_35 & other_ops_36_valid_down; // @[MapS.scala 23:83]
  assign _T_37 = _T_36 & other_ops_37_valid_down; // @[MapS.scala 23:83]
  assign _T_38 = _T_37 & other_ops_38_valid_down; // @[MapS.scala 23:83]
  assign _T_39 = _T_38 & other_ops_39_valid_down; // @[MapS.scala 23:83]
  assign _T_40 = _T_39 & other_ops_40_valid_down; // @[MapS.scala 23:83]
  assign _T_41 = _T_40 & other_ops_41_valid_down; // @[MapS.scala 23:83]
  assign _T_42 = _T_41 & other_ops_42_valid_down; // @[MapS.scala 23:83]
  assign _T_43 = _T_42 & other_ops_43_valid_down; // @[MapS.scala 23:83]
  assign _T_44 = _T_43 & other_ops_44_valid_down; // @[MapS.scala 23:83]
  assign _T_45 = _T_44 & other_ops_45_valid_down; // @[MapS.scala 23:83]
  assign _T_46 = _T_45 & other_ops_46_valid_down; // @[MapS.scala 23:83]
  assign _T_47 = _T_46 & other_ops_47_valid_down; // @[MapS.scala 23:83]
  assign _T_48 = _T_47 & other_ops_48_valid_down; // @[MapS.scala 23:83]
  assign _T_49 = _T_48 & other_ops_49_valid_down; // @[MapS.scala 23:83]
  assign _T_50 = _T_49 & other_ops_50_valid_down; // @[MapS.scala 23:83]
  assign _T_51 = _T_50 & other_ops_51_valid_down; // @[MapS.scala 23:83]
  assign _T_52 = _T_51 & other_ops_52_valid_down; // @[MapS.scala 23:83]
  assign _T_53 = _T_52 & other_ops_53_valid_down; // @[MapS.scala 23:83]
  assign _T_54 = _T_53 & other_ops_54_valid_down; // @[MapS.scala 23:83]
  assign _T_55 = _T_54 & other_ops_55_valid_down; // @[MapS.scala 23:83]
  assign _T_56 = _T_55 & other_ops_56_valid_down; // @[MapS.scala 23:83]
  assign _T_57 = _T_56 & other_ops_57_valid_down; // @[MapS.scala 23:83]
  assign _T_58 = _T_57 & other_ops_58_valid_down; // @[MapS.scala 23:83]
  assign _T_59 = _T_58 & other_ops_59_valid_down; // @[MapS.scala 23:83]
  assign _T_60 = _T_59 & other_ops_60_valid_down; // @[MapS.scala 23:83]
  assign _T_61 = _T_60 & other_ops_61_valid_down; // @[MapS.scala 23:83]
  assign _T_62 = _T_61 & other_ops_62_valid_down; // @[MapS.scala 23:83]
  assign _T_63 = _T_62 & other_ops_63_valid_down; // @[MapS.scala 23:83]
  assign _T_64 = _T_63 & other_ops_64_valid_down; // @[MapS.scala 23:83]
  assign _T_65 = _T_64 & other_ops_65_valid_down; // @[MapS.scala 23:83]
  assign _T_66 = _T_65 & other_ops_66_valid_down; // @[MapS.scala 23:83]
  assign _T_67 = _T_66 & other_ops_67_valid_down; // @[MapS.scala 23:83]
  assign _T_68 = _T_67 & other_ops_68_valid_down; // @[MapS.scala 23:83]
  assign _T_69 = _T_68 & other_ops_69_valid_down; // @[MapS.scala 23:83]
  assign _T_70 = _T_69 & other_ops_70_valid_down; // @[MapS.scala 23:83]
  assign _T_71 = _T_70 & other_ops_71_valid_down; // @[MapS.scala 23:83]
  assign _T_72 = _T_71 & other_ops_72_valid_down; // @[MapS.scala 23:83]
  assign _T_73 = _T_72 & other_ops_73_valid_down; // @[MapS.scala 23:83]
  assign _T_74 = _T_73 & other_ops_74_valid_down; // @[MapS.scala 23:83]
  assign _T_75 = _T_74 & other_ops_75_valid_down; // @[MapS.scala 23:83]
  assign _T_76 = _T_75 & other_ops_76_valid_down; // @[MapS.scala 23:83]
  assign _T_77 = _T_76 & other_ops_77_valid_down; // @[MapS.scala 23:83]
  assign _T_78 = _T_77 & other_ops_78_valid_down; // @[MapS.scala 23:83]
  assign _T_79 = _T_78 & other_ops_79_valid_down; // @[MapS.scala 23:83]
  assign _T_80 = _T_79 & other_ops_80_valid_down; // @[MapS.scala 23:83]
  assign _T_81 = _T_80 & other_ops_81_valid_down; // @[MapS.scala 23:83]
  assign _T_82 = _T_81 & other_ops_82_valid_down; // @[MapS.scala 23:83]
  assign _T_83 = _T_82 & other_ops_83_valid_down; // @[MapS.scala 23:83]
  assign _T_84 = _T_83 & other_ops_84_valid_down; // @[MapS.scala 23:83]
  assign _T_85 = _T_84 & other_ops_85_valid_down; // @[MapS.scala 23:83]
  assign _T_86 = _T_85 & other_ops_86_valid_down; // @[MapS.scala 23:83]
  assign _T_87 = _T_86 & other_ops_87_valid_down; // @[MapS.scala 23:83]
  assign _T_88 = _T_87 & other_ops_88_valid_down; // @[MapS.scala 23:83]
  assign _T_89 = _T_88 & other_ops_89_valid_down; // @[MapS.scala 23:83]
  assign _T_90 = _T_89 & other_ops_90_valid_down; // @[MapS.scala 23:83]
  assign _T_91 = _T_90 & other_ops_91_valid_down; // @[MapS.scala 23:83]
  assign _T_92 = _T_91 & other_ops_92_valid_down; // @[MapS.scala 23:83]
  assign _T_93 = _T_92 & other_ops_93_valid_down; // @[MapS.scala 23:83]
  assign _T_94 = _T_93 & other_ops_94_valid_down; // @[MapS.scala 23:83]
  assign _T_95 = _T_94 & other_ops_95_valid_down; // @[MapS.scala 23:83]
  assign _T_96 = _T_95 & other_ops_96_valid_down; // @[MapS.scala 23:83]
  assign _T_97 = _T_96 & other_ops_97_valid_down; // @[MapS.scala 23:83]
  assign _T_98 = _T_97 & other_ops_98_valid_down; // @[MapS.scala 23:83]
  assign _T_99 = _T_98 & other_ops_99_valid_down; // @[MapS.scala 23:83]
  assign _T_100 = _T_99 & other_ops_100_valid_down; // @[MapS.scala 23:83]
  assign _T_101 = _T_100 & other_ops_101_valid_down; // @[MapS.scala 23:83]
  assign _T_102 = _T_101 & other_ops_102_valid_down; // @[MapS.scala 23:83]
  assign _T_103 = _T_102 & other_ops_103_valid_down; // @[MapS.scala 23:83]
  assign _T_104 = _T_103 & other_ops_104_valid_down; // @[MapS.scala 23:83]
  assign _T_105 = _T_104 & other_ops_105_valid_down; // @[MapS.scala 23:83]
  assign _T_106 = _T_105 & other_ops_106_valid_down; // @[MapS.scala 23:83]
  assign _T_107 = _T_106 & other_ops_107_valid_down; // @[MapS.scala 23:83]
  assign _T_108 = _T_107 & other_ops_108_valid_down; // @[MapS.scala 23:83]
  assign _T_109 = _T_108 & other_ops_109_valid_down; // @[MapS.scala 23:83]
  assign _T_110 = _T_109 & other_ops_110_valid_down; // @[MapS.scala 23:83]
  assign _T_111 = _T_110 & other_ops_111_valid_down; // @[MapS.scala 23:83]
  assign _T_112 = _T_111 & other_ops_112_valid_down; // @[MapS.scala 23:83]
  assign _T_113 = _T_112 & other_ops_113_valid_down; // @[MapS.scala 23:83]
  assign _T_114 = _T_113 & other_ops_114_valid_down; // @[MapS.scala 23:83]
  assign _T_115 = _T_114 & other_ops_115_valid_down; // @[MapS.scala 23:83]
  assign _T_116 = _T_115 & other_ops_116_valid_down; // @[MapS.scala 23:83]
  assign _T_117 = _T_116 & other_ops_117_valid_down; // @[MapS.scala 23:83]
  assign _T_118 = _T_117 & other_ops_118_valid_down; // @[MapS.scala 23:83]
  assign _T_119 = _T_118 & other_ops_119_valid_down; // @[MapS.scala 23:83]
  assign _T_120 = _T_119 & other_ops_120_valid_down; // @[MapS.scala 23:83]
  assign _T_121 = _T_120 & other_ops_121_valid_down; // @[MapS.scala 23:83]
  assign _T_122 = _T_121 & other_ops_122_valid_down; // @[MapS.scala 23:83]
  assign _T_123 = _T_122 & other_ops_123_valid_down; // @[MapS.scala 23:83]
  assign _T_124 = _T_123 & other_ops_124_valid_down; // @[MapS.scala 23:83]
  assign _T_125 = _T_124 & other_ops_125_valid_down; // @[MapS.scala 23:83]
  assign _T_126 = _T_125 & other_ops_126_valid_down; // @[MapS.scala 23:83]
  assign _T_127 = _T_126 & other_ops_127_valid_down; // @[MapS.scala 23:83]
  assign _T_128 = _T_127 & other_ops_128_valid_down; // @[MapS.scala 23:83]
  assign _T_129 = _T_128 & other_ops_129_valid_down; // @[MapS.scala 23:83]
  assign _T_130 = _T_129 & other_ops_130_valid_down; // @[MapS.scala 23:83]
  assign _T_131 = _T_130 & other_ops_131_valid_down; // @[MapS.scala 23:83]
  assign _T_132 = _T_131 & other_ops_132_valid_down; // @[MapS.scala 23:83]
  assign _T_133 = _T_132 & other_ops_133_valid_down; // @[MapS.scala 23:83]
  assign _T_134 = _T_133 & other_ops_134_valid_down; // @[MapS.scala 23:83]
  assign _T_135 = _T_134 & other_ops_135_valid_down; // @[MapS.scala 23:83]
  assign _T_136 = _T_135 & other_ops_136_valid_down; // @[MapS.scala 23:83]
  assign _T_137 = _T_136 & other_ops_137_valid_down; // @[MapS.scala 23:83]
  assign _T_138 = _T_137 & other_ops_138_valid_down; // @[MapS.scala 23:83]
  assign _T_139 = _T_138 & other_ops_139_valid_down; // @[MapS.scala 23:83]
  assign _T_140 = _T_139 & other_ops_140_valid_down; // @[MapS.scala 23:83]
  assign _T_141 = _T_140 & other_ops_141_valid_down; // @[MapS.scala 23:83]
  assign _T_142 = _T_141 & other_ops_142_valid_down; // @[MapS.scala 23:83]
  assign _T_143 = _T_142 & other_ops_143_valid_down; // @[MapS.scala 23:83]
  assign _T_144 = _T_143 & other_ops_144_valid_down; // @[MapS.scala 23:83]
  assign _T_145 = _T_144 & other_ops_145_valid_down; // @[MapS.scala 23:83]
  assign _T_146 = _T_145 & other_ops_146_valid_down; // @[MapS.scala 23:83]
  assign _T_147 = _T_146 & other_ops_147_valid_down; // @[MapS.scala 23:83]
  assign _T_148 = _T_147 & other_ops_148_valid_down; // @[MapS.scala 23:83]
  assign _T_149 = _T_148 & other_ops_149_valid_down; // @[MapS.scala 23:83]
  assign _T_150 = _T_149 & other_ops_150_valid_down; // @[MapS.scala 23:83]
  assign _T_151 = _T_150 & other_ops_151_valid_down; // @[MapS.scala 23:83]
  assign _T_152 = _T_151 & other_ops_152_valid_down; // @[MapS.scala 23:83]
  assign _T_153 = _T_152 & other_ops_153_valid_down; // @[MapS.scala 23:83]
  assign _T_154 = _T_153 & other_ops_154_valid_down; // @[MapS.scala 23:83]
  assign _T_155 = _T_154 & other_ops_155_valid_down; // @[MapS.scala 23:83]
  assign _T_156 = _T_155 & other_ops_156_valid_down; // @[MapS.scala 23:83]
  assign _T_157 = _T_156 & other_ops_157_valid_down; // @[MapS.scala 23:83]
  assign _T_158 = _T_157 & other_ops_158_valid_down; // @[MapS.scala 23:83]
  assign _T_159 = _T_158 & other_ops_159_valid_down; // @[MapS.scala 23:83]
  assign _T_160 = _T_159 & other_ops_160_valid_down; // @[MapS.scala 23:83]
  assign _T_161 = _T_160 & other_ops_161_valid_down; // @[MapS.scala 23:83]
  assign _T_162 = _T_161 & other_ops_162_valid_down; // @[MapS.scala 23:83]
  assign _T_163 = _T_162 & other_ops_163_valid_down; // @[MapS.scala 23:83]
  assign _T_164 = _T_163 & other_ops_164_valid_down; // @[MapS.scala 23:83]
  assign _T_165 = _T_164 & other_ops_165_valid_down; // @[MapS.scala 23:83]
  assign _T_166 = _T_165 & other_ops_166_valid_down; // @[MapS.scala 23:83]
  assign _T_167 = _T_166 & other_ops_167_valid_down; // @[MapS.scala 23:83]
  assign _T_168 = _T_167 & other_ops_168_valid_down; // @[MapS.scala 23:83]
  assign _T_169 = _T_168 & other_ops_169_valid_down; // @[MapS.scala 23:83]
  assign _T_170 = _T_169 & other_ops_170_valid_down; // @[MapS.scala 23:83]
  assign _T_171 = _T_170 & other_ops_171_valid_down; // @[MapS.scala 23:83]
  assign _T_172 = _T_171 & other_ops_172_valid_down; // @[MapS.scala 23:83]
  assign _T_173 = _T_172 & other_ops_173_valid_down; // @[MapS.scala 23:83]
  assign _T_174 = _T_173 & other_ops_174_valid_down; // @[MapS.scala 23:83]
  assign _T_175 = _T_174 & other_ops_175_valid_down; // @[MapS.scala 23:83]
  assign _T_176 = _T_175 & other_ops_176_valid_down; // @[MapS.scala 23:83]
  assign _T_177 = _T_176 & other_ops_177_valid_down; // @[MapS.scala 23:83]
  assign _T_178 = _T_177 & other_ops_178_valid_down; // @[MapS.scala 23:83]
  assign _T_179 = _T_178 & other_ops_179_valid_down; // @[MapS.scala 23:83]
  assign _T_180 = _T_179 & other_ops_180_valid_down; // @[MapS.scala 23:83]
  assign _T_181 = _T_180 & other_ops_181_valid_down; // @[MapS.scala 23:83]
  assign _T_182 = _T_181 & other_ops_182_valid_down; // @[MapS.scala 23:83]
  assign _T_183 = _T_182 & other_ops_183_valid_down; // @[MapS.scala 23:83]
  assign _T_184 = _T_183 & other_ops_184_valid_down; // @[MapS.scala 23:83]
  assign _T_185 = _T_184 & other_ops_185_valid_down; // @[MapS.scala 23:83]
  assign _T_186 = _T_185 & other_ops_186_valid_down; // @[MapS.scala 23:83]
  assign _T_187 = _T_186 & other_ops_187_valid_down; // @[MapS.scala 23:83]
  assign _T_188 = _T_187 & other_ops_188_valid_down; // @[MapS.scala 23:83]
  assign _T_189 = _T_188 & other_ops_189_valid_down; // @[MapS.scala 23:83]
  assign _T_190 = _T_189 & other_ops_190_valid_down; // @[MapS.scala 23:83]
  assign _T_191 = _T_190 & other_ops_191_valid_down; // @[MapS.scala 23:83]
  assign _T_192 = _T_191 & other_ops_192_valid_down; // @[MapS.scala 23:83]
  assign _T_193 = _T_192 & other_ops_193_valid_down; // @[MapS.scala 23:83]
  assign _T_194 = _T_193 & other_ops_194_valid_down; // @[MapS.scala 23:83]
  assign _T_195 = _T_194 & other_ops_195_valid_down; // @[MapS.scala 23:83]
  assign _T_196 = _T_195 & other_ops_196_valid_down; // @[MapS.scala 23:83]
  assign _T_197 = _T_196 & other_ops_197_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_197 & other_ops_198_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign O_3 = other_ops_2_O; // @[MapS.scala 21:12]
  assign O_4 = other_ops_3_O; // @[MapS.scala 21:12]
  assign O_5 = other_ops_4_O; // @[MapS.scala 21:12]
  assign O_6 = other_ops_5_O; // @[MapS.scala 21:12]
  assign O_7 = other_ops_6_O; // @[MapS.scala 21:12]
  assign O_8 = other_ops_7_O; // @[MapS.scala 21:12]
  assign O_9 = other_ops_8_O; // @[MapS.scala 21:12]
  assign O_10 = other_ops_9_O; // @[MapS.scala 21:12]
  assign O_11 = other_ops_10_O; // @[MapS.scala 21:12]
  assign O_12 = other_ops_11_O; // @[MapS.scala 21:12]
  assign O_13 = other_ops_12_O; // @[MapS.scala 21:12]
  assign O_14 = other_ops_13_O; // @[MapS.scala 21:12]
  assign O_15 = other_ops_14_O; // @[MapS.scala 21:12]
  assign O_16 = other_ops_15_O; // @[MapS.scala 21:12]
  assign O_17 = other_ops_16_O; // @[MapS.scala 21:12]
  assign O_18 = other_ops_17_O; // @[MapS.scala 21:12]
  assign O_19 = other_ops_18_O; // @[MapS.scala 21:12]
  assign O_20 = other_ops_19_O; // @[MapS.scala 21:12]
  assign O_21 = other_ops_20_O; // @[MapS.scala 21:12]
  assign O_22 = other_ops_21_O; // @[MapS.scala 21:12]
  assign O_23 = other_ops_22_O; // @[MapS.scala 21:12]
  assign O_24 = other_ops_23_O; // @[MapS.scala 21:12]
  assign O_25 = other_ops_24_O; // @[MapS.scala 21:12]
  assign O_26 = other_ops_25_O; // @[MapS.scala 21:12]
  assign O_27 = other_ops_26_O; // @[MapS.scala 21:12]
  assign O_28 = other_ops_27_O; // @[MapS.scala 21:12]
  assign O_29 = other_ops_28_O; // @[MapS.scala 21:12]
  assign O_30 = other_ops_29_O; // @[MapS.scala 21:12]
  assign O_31 = other_ops_30_O; // @[MapS.scala 21:12]
  assign O_32 = other_ops_31_O; // @[MapS.scala 21:12]
  assign O_33 = other_ops_32_O; // @[MapS.scala 21:12]
  assign O_34 = other_ops_33_O; // @[MapS.scala 21:12]
  assign O_35 = other_ops_34_O; // @[MapS.scala 21:12]
  assign O_36 = other_ops_35_O; // @[MapS.scala 21:12]
  assign O_37 = other_ops_36_O; // @[MapS.scala 21:12]
  assign O_38 = other_ops_37_O; // @[MapS.scala 21:12]
  assign O_39 = other_ops_38_O; // @[MapS.scala 21:12]
  assign O_40 = other_ops_39_O; // @[MapS.scala 21:12]
  assign O_41 = other_ops_40_O; // @[MapS.scala 21:12]
  assign O_42 = other_ops_41_O; // @[MapS.scala 21:12]
  assign O_43 = other_ops_42_O; // @[MapS.scala 21:12]
  assign O_44 = other_ops_43_O; // @[MapS.scala 21:12]
  assign O_45 = other_ops_44_O; // @[MapS.scala 21:12]
  assign O_46 = other_ops_45_O; // @[MapS.scala 21:12]
  assign O_47 = other_ops_46_O; // @[MapS.scala 21:12]
  assign O_48 = other_ops_47_O; // @[MapS.scala 21:12]
  assign O_49 = other_ops_48_O; // @[MapS.scala 21:12]
  assign O_50 = other_ops_49_O; // @[MapS.scala 21:12]
  assign O_51 = other_ops_50_O; // @[MapS.scala 21:12]
  assign O_52 = other_ops_51_O; // @[MapS.scala 21:12]
  assign O_53 = other_ops_52_O; // @[MapS.scala 21:12]
  assign O_54 = other_ops_53_O; // @[MapS.scala 21:12]
  assign O_55 = other_ops_54_O; // @[MapS.scala 21:12]
  assign O_56 = other_ops_55_O; // @[MapS.scala 21:12]
  assign O_57 = other_ops_56_O; // @[MapS.scala 21:12]
  assign O_58 = other_ops_57_O; // @[MapS.scala 21:12]
  assign O_59 = other_ops_58_O; // @[MapS.scala 21:12]
  assign O_60 = other_ops_59_O; // @[MapS.scala 21:12]
  assign O_61 = other_ops_60_O; // @[MapS.scala 21:12]
  assign O_62 = other_ops_61_O; // @[MapS.scala 21:12]
  assign O_63 = other_ops_62_O; // @[MapS.scala 21:12]
  assign O_64 = other_ops_63_O; // @[MapS.scala 21:12]
  assign O_65 = other_ops_64_O; // @[MapS.scala 21:12]
  assign O_66 = other_ops_65_O; // @[MapS.scala 21:12]
  assign O_67 = other_ops_66_O; // @[MapS.scala 21:12]
  assign O_68 = other_ops_67_O; // @[MapS.scala 21:12]
  assign O_69 = other_ops_68_O; // @[MapS.scala 21:12]
  assign O_70 = other_ops_69_O; // @[MapS.scala 21:12]
  assign O_71 = other_ops_70_O; // @[MapS.scala 21:12]
  assign O_72 = other_ops_71_O; // @[MapS.scala 21:12]
  assign O_73 = other_ops_72_O; // @[MapS.scala 21:12]
  assign O_74 = other_ops_73_O; // @[MapS.scala 21:12]
  assign O_75 = other_ops_74_O; // @[MapS.scala 21:12]
  assign O_76 = other_ops_75_O; // @[MapS.scala 21:12]
  assign O_77 = other_ops_76_O; // @[MapS.scala 21:12]
  assign O_78 = other_ops_77_O; // @[MapS.scala 21:12]
  assign O_79 = other_ops_78_O; // @[MapS.scala 21:12]
  assign O_80 = other_ops_79_O; // @[MapS.scala 21:12]
  assign O_81 = other_ops_80_O; // @[MapS.scala 21:12]
  assign O_82 = other_ops_81_O; // @[MapS.scala 21:12]
  assign O_83 = other_ops_82_O; // @[MapS.scala 21:12]
  assign O_84 = other_ops_83_O; // @[MapS.scala 21:12]
  assign O_85 = other_ops_84_O; // @[MapS.scala 21:12]
  assign O_86 = other_ops_85_O; // @[MapS.scala 21:12]
  assign O_87 = other_ops_86_O; // @[MapS.scala 21:12]
  assign O_88 = other_ops_87_O; // @[MapS.scala 21:12]
  assign O_89 = other_ops_88_O; // @[MapS.scala 21:12]
  assign O_90 = other_ops_89_O; // @[MapS.scala 21:12]
  assign O_91 = other_ops_90_O; // @[MapS.scala 21:12]
  assign O_92 = other_ops_91_O; // @[MapS.scala 21:12]
  assign O_93 = other_ops_92_O; // @[MapS.scala 21:12]
  assign O_94 = other_ops_93_O; // @[MapS.scala 21:12]
  assign O_95 = other_ops_94_O; // @[MapS.scala 21:12]
  assign O_96 = other_ops_95_O; // @[MapS.scala 21:12]
  assign O_97 = other_ops_96_O; // @[MapS.scala 21:12]
  assign O_98 = other_ops_97_O; // @[MapS.scala 21:12]
  assign O_99 = other_ops_98_O; // @[MapS.scala 21:12]
  assign O_100 = other_ops_99_O; // @[MapS.scala 21:12]
  assign O_101 = other_ops_100_O; // @[MapS.scala 21:12]
  assign O_102 = other_ops_101_O; // @[MapS.scala 21:12]
  assign O_103 = other_ops_102_O; // @[MapS.scala 21:12]
  assign O_104 = other_ops_103_O; // @[MapS.scala 21:12]
  assign O_105 = other_ops_104_O; // @[MapS.scala 21:12]
  assign O_106 = other_ops_105_O; // @[MapS.scala 21:12]
  assign O_107 = other_ops_106_O; // @[MapS.scala 21:12]
  assign O_108 = other_ops_107_O; // @[MapS.scala 21:12]
  assign O_109 = other_ops_108_O; // @[MapS.scala 21:12]
  assign O_110 = other_ops_109_O; // @[MapS.scala 21:12]
  assign O_111 = other_ops_110_O; // @[MapS.scala 21:12]
  assign O_112 = other_ops_111_O; // @[MapS.scala 21:12]
  assign O_113 = other_ops_112_O; // @[MapS.scala 21:12]
  assign O_114 = other_ops_113_O; // @[MapS.scala 21:12]
  assign O_115 = other_ops_114_O; // @[MapS.scala 21:12]
  assign O_116 = other_ops_115_O; // @[MapS.scala 21:12]
  assign O_117 = other_ops_116_O; // @[MapS.scala 21:12]
  assign O_118 = other_ops_117_O; // @[MapS.scala 21:12]
  assign O_119 = other_ops_118_O; // @[MapS.scala 21:12]
  assign O_120 = other_ops_119_O; // @[MapS.scala 21:12]
  assign O_121 = other_ops_120_O; // @[MapS.scala 21:12]
  assign O_122 = other_ops_121_O; // @[MapS.scala 21:12]
  assign O_123 = other_ops_122_O; // @[MapS.scala 21:12]
  assign O_124 = other_ops_123_O; // @[MapS.scala 21:12]
  assign O_125 = other_ops_124_O; // @[MapS.scala 21:12]
  assign O_126 = other_ops_125_O; // @[MapS.scala 21:12]
  assign O_127 = other_ops_126_O; // @[MapS.scala 21:12]
  assign O_128 = other_ops_127_O; // @[MapS.scala 21:12]
  assign O_129 = other_ops_128_O; // @[MapS.scala 21:12]
  assign O_130 = other_ops_129_O; // @[MapS.scala 21:12]
  assign O_131 = other_ops_130_O; // @[MapS.scala 21:12]
  assign O_132 = other_ops_131_O; // @[MapS.scala 21:12]
  assign O_133 = other_ops_132_O; // @[MapS.scala 21:12]
  assign O_134 = other_ops_133_O; // @[MapS.scala 21:12]
  assign O_135 = other_ops_134_O; // @[MapS.scala 21:12]
  assign O_136 = other_ops_135_O; // @[MapS.scala 21:12]
  assign O_137 = other_ops_136_O; // @[MapS.scala 21:12]
  assign O_138 = other_ops_137_O; // @[MapS.scala 21:12]
  assign O_139 = other_ops_138_O; // @[MapS.scala 21:12]
  assign O_140 = other_ops_139_O; // @[MapS.scala 21:12]
  assign O_141 = other_ops_140_O; // @[MapS.scala 21:12]
  assign O_142 = other_ops_141_O; // @[MapS.scala 21:12]
  assign O_143 = other_ops_142_O; // @[MapS.scala 21:12]
  assign O_144 = other_ops_143_O; // @[MapS.scala 21:12]
  assign O_145 = other_ops_144_O; // @[MapS.scala 21:12]
  assign O_146 = other_ops_145_O; // @[MapS.scala 21:12]
  assign O_147 = other_ops_146_O; // @[MapS.scala 21:12]
  assign O_148 = other_ops_147_O; // @[MapS.scala 21:12]
  assign O_149 = other_ops_148_O; // @[MapS.scala 21:12]
  assign O_150 = other_ops_149_O; // @[MapS.scala 21:12]
  assign O_151 = other_ops_150_O; // @[MapS.scala 21:12]
  assign O_152 = other_ops_151_O; // @[MapS.scala 21:12]
  assign O_153 = other_ops_152_O; // @[MapS.scala 21:12]
  assign O_154 = other_ops_153_O; // @[MapS.scala 21:12]
  assign O_155 = other_ops_154_O; // @[MapS.scala 21:12]
  assign O_156 = other_ops_155_O; // @[MapS.scala 21:12]
  assign O_157 = other_ops_156_O; // @[MapS.scala 21:12]
  assign O_158 = other_ops_157_O; // @[MapS.scala 21:12]
  assign O_159 = other_ops_158_O; // @[MapS.scala 21:12]
  assign O_160 = other_ops_159_O; // @[MapS.scala 21:12]
  assign O_161 = other_ops_160_O; // @[MapS.scala 21:12]
  assign O_162 = other_ops_161_O; // @[MapS.scala 21:12]
  assign O_163 = other_ops_162_O; // @[MapS.scala 21:12]
  assign O_164 = other_ops_163_O; // @[MapS.scala 21:12]
  assign O_165 = other_ops_164_O; // @[MapS.scala 21:12]
  assign O_166 = other_ops_165_O; // @[MapS.scala 21:12]
  assign O_167 = other_ops_166_O; // @[MapS.scala 21:12]
  assign O_168 = other_ops_167_O; // @[MapS.scala 21:12]
  assign O_169 = other_ops_168_O; // @[MapS.scala 21:12]
  assign O_170 = other_ops_169_O; // @[MapS.scala 21:12]
  assign O_171 = other_ops_170_O; // @[MapS.scala 21:12]
  assign O_172 = other_ops_171_O; // @[MapS.scala 21:12]
  assign O_173 = other_ops_172_O; // @[MapS.scala 21:12]
  assign O_174 = other_ops_173_O; // @[MapS.scala 21:12]
  assign O_175 = other_ops_174_O; // @[MapS.scala 21:12]
  assign O_176 = other_ops_175_O; // @[MapS.scala 21:12]
  assign O_177 = other_ops_176_O; // @[MapS.scala 21:12]
  assign O_178 = other_ops_177_O; // @[MapS.scala 21:12]
  assign O_179 = other_ops_178_O; // @[MapS.scala 21:12]
  assign O_180 = other_ops_179_O; // @[MapS.scala 21:12]
  assign O_181 = other_ops_180_O; // @[MapS.scala 21:12]
  assign O_182 = other_ops_181_O; // @[MapS.scala 21:12]
  assign O_183 = other_ops_182_O; // @[MapS.scala 21:12]
  assign O_184 = other_ops_183_O; // @[MapS.scala 21:12]
  assign O_185 = other_ops_184_O; // @[MapS.scala 21:12]
  assign O_186 = other_ops_185_O; // @[MapS.scala 21:12]
  assign O_187 = other_ops_186_O; // @[MapS.scala 21:12]
  assign O_188 = other_ops_187_O; // @[MapS.scala 21:12]
  assign O_189 = other_ops_188_O; // @[MapS.scala 21:12]
  assign O_190 = other_ops_189_O; // @[MapS.scala 21:12]
  assign O_191 = other_ops_190_O; // @[MapS.scala 21:12]
  assign O_192 = other_ops_191_O; // @[MapS.scala 21:12]
  assign O_193 = other_ops_192_O; // @[MapS.scala 21:12]
  assign O_194 = other_ops_193_O; // @[MapS.scala 21:12]
  assign O_195 = other_ops_194_O; // @[MapS.scala 21:12]
  assign O_196 = other_ops_195_O; // @[MapS.scala 21:12]
  assign O_197 = other_ops_196_O; // @[MapS.scala 21:12]
  assign O_198 = other_ops_197_O; // @[MapS.scala 21:12]
  assign O_199 = other_ops_198_O; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I = I_0; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I = I_1; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I = I_2; // @[MapS.scala 20:41]
  assign other_ops_2_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_2_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I = I_3; // @[MapS.scala 20:41]
  assign other_ops_3_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_3_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I = I_4; // @[MapS.scala 20:41]
  assign other_ops_4_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_4_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I = I_5; // @[MapS.scala 20:41]
  assign other_ops_5_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_5_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I = I_6; // @[MapS.scala 20:41]
  assign other_ops_6_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_6_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I = I_7; // @[MapS.scala 20:41]
  assign other_ops_7_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_7_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I = I_8; // @[MapS.scala 20:41]
  assign other_ops_8_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_8_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I = I_9; // @[MapS.scala 20:41]
  assign other_ops_9_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_9_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I = I_10; // @[MapS.scala 20:41]
  assign other_ops_10_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_10_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I = I_11; // @[MapS.scala 20:41]
  assign other_ops_11_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_11_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I = I_12; // @[MapS.scala 20:41]
  assign other_ops_12_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_12_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I = I_13; // @[MapS.scala 20:41]
  assign other_ops_13_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_13_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I = I_14; // @[MapS.scala 20:41]
  assign other_ops_14_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_14_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I = I_15; // @[MapS.scala 20:41]
  assign other_ops_15_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_15_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_15_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_15_I = I_16; // @[MapS.scala 20:41]
  assign other_ops_16_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_16_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_16_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_16_I = I_17; // @[MapS.scala 20:41]
  assign other_ops_17_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_17_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_17_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_17_I = I_18; // @[MapS.scala 20:41]
  assign other_ops_18_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_18_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_18_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_18_I = I_19; // @[MapS.scala 20:41]
  assign other_ops_19_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_19_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_19_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_19_I = I_20; // @[MapS.scala 20:41]
  assign other_ops_20_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_20_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_20_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_20_I = I_21; // @[MapS.scala 20:41]
  assign other_ops_21_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_21_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_21_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_21_I = I_22; // @[MapS.scala 20:41]
  assign other_ops_22_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_22_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_22_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_22_I = I_23; // @[MapS.scala 20:41]
  assign other_ops_23_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_23_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_23_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_23_I = I_24; // @[MapS.scala 20:41]
  assign other_ops_24_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_24_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_24_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_24_I = I_25; // @[MapS.scala 20:41]
  assign other_ops_25_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_25_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_25_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_25_I = I_26; // @[MapS.scala 20:41]
  assign other_ops_26_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_26_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_26_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_26_I = I_27; // @[MapS.scala 20:41]
  assign other_ops_27_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_27_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_27_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_27_I = I_28; // @[MapS.scala 20:41]
  assign other_ops_28_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_28_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_28_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_28_I = I_29; // @[MapS.scala 20:41]
  assign other_ops_29_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_29_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_29_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_29_I = I_30; // @[MapS.scala 20:41]
  assign other_ops_30_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_30_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_30_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_30_I = I_31; // @[MapS.scala 20:41]
  assign other_ops_31_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_31_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_31_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_31_I = I_32; // @[MapS.scala 20:41]
  assign other_ops_32_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_32_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_32_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_32_I = I_33; // @[MapS.scala 20:41]
  assign other_ops_33_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_33_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_33_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_33_I = I_34; // @[MapS.scala 20:41]
  assign other_ops_34_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_34_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_34_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_34_I = I_35; // @[MapS.scala 20:41]
  assign other_ops_35_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_35_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_35_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_35_I = I_36; // @[MapS.scala 20:41]
  assign other_ops_36_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_36_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_36_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_36_I = I_37; // @[MapS.scala 20:41]
  assign other_ops_37_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_37_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_37_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_37_I = I_38; // @[MapS.scala 20:41]
  assign other_ops_38_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_38_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_38_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_38_I = I_39; // @[MapS.scala 20:41]
  assign other_ops_39_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_39_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_39_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_39_I = I_40; // @[MapS.scala 20:41]
  assign other_ops_40_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_40_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_40_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_40_I = I_41; // @[MapS.scala 20:41]
  assign other_ops_41_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_41_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_41_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_41_I = I_42; // @[MapS.scala 20:41]
  assign other_ops_42_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_42_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_42_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_42_I = I_43; // @[MapS.scala 20:41]
  assign other_ops_43_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_43_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_43_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_43_I = I_44; // @[MapS.scala 20:41]
  assign other_ops_44_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_44_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_44_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_44_I = I_45; // @[MapS.scala 20:41]
  assign other_ops_45_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_45_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_45_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_45_I = I_46; // @[MapS.scala 20:41]
  assign other_ops_46_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_46_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_46_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_46_I = I_47; // @[MapS.scala 20:41]
  assign other_ops_47_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_47_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_47_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_47_I = I_48; // @[MapS.scala 20:41]
  assign other_ops_48_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_48_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_48_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_48_I = I_49; // @[MapS.scala 20:41]
  assign other_ops_49_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_49_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_49_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_49_I = I_50; // @[MapS.scala 20:41]
  assign other_ops_50_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_50_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_50_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_50_I = I_51; // @[MapS.scala 20:41]
  assign other_ops_51_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_51_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_51_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_51_I = I_52; // @[MapS.scala 20:41]
  assign other_ops_52_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_52_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_52_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_52_I = I_53; // @[MapS.scala 20:41]
  assign other_ops_53_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_53_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_53_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_53_I = I_54; // @[MapS.scala 20:41]
  assign other_ops_54_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_54_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_54_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_54_I = I_55; // @[MapS.scala 20:41]
  assign other_ops_55_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_55_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_55_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_55_I = I_56; // @[MapS.scala 20:41]
  assign other_ops_56_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_56_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_56_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_56_I = I_57; // @[MapS.scala 20:41]
  assign other_ops_57_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_57_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_57_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_57_I = I_58; // @[MapS.scala 20:41]
  assign other_ops_58_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_58_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_58_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_58_I = I_59; // @[MapS.scala 20:41]
  assign other_ops_59_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_59_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_59_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_59_I = I_60; // @[MapS.scala 20:41]
  assign other_ops_60_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_60_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_60_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_60_I = I_61; // @[MapS.scala 20:41]
  assign other_ops_61_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_61_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_61_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_61_I = I_62; // @[MapS.scala 20:41]
  assign other_ops_62_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_62_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_62_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_62_I = I_63; // @[MapS.scala 20:41]
  assign other_ops_63_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_63_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_63_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_63_I = I_64; // @[MapS.scala 20:41]
  assign other_ops_64_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_64_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_64_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_64_I = I_65; // @[MapS.scala 20:41]
  assign other_ops_65_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_65_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_65_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_65_I = I_66; // @[MapS.scala 20:41]
  assign other_ops_66_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_66_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_66_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_66_I = I_67; // @[MapS.scala 20:41]
  assign other_ops_67_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_67_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_67_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_67_I = I_68; // @[MapS.scala 20:41]
  assign other_ops_68_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_68_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_68_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_68_I = I_69; // @[MapS.scala 20:41]
  assign other_ops_69_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_69_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_69_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_69_I = I_70; // @[MapS.scala 20:41]
  assign other_ops_70_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_70_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_70_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_70_I = I_71; // @[MapS.scala 20:41]
  assign other_ops_71_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_71_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_71_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_71_I = I_72; // @[MapS.scala 20:41]
  assign other_ops_72_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_72_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_72_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_72_I = I_73; // @[MapS.scala 20:41]
  assign other_ops_73_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_73_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_73_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_73_I = I_74; // @[MapS.scala 20:41]
  assign other_ops_74_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_74_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_74_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_74_I = I_75; // @[MapS.scala 20:41]
  assign other_ops_75_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_75_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_75_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_75_I = I_76; // @[MapS.scala 20:41]
  assign other_ops_76_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_76_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_76_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_76_I = I_77; // @[MapS.scala 20:41]
  assign other_ops_77_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_77_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_77_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_77_I = I_78; // @[MapS.scala 20:41]
  assign other_ops_78_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_78_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_78_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_78_I = I_79; // @[MapS.scala 20:41]
  assign other_ops_79_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_79_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_79_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_79_I = I_80; // @[MapS.scala 20:41]
  assign other_ops_80_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_80_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_80_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_80_I = I_81; // @[MapS.scala 20:41]
  assign other_ops_81_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_81_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_81_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_81_I = I_82; // @[MapS.scala 20:41]
  assign other_ops_82_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_82_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_82_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_82_I = I_83; // @[MapS.scala 20:41]
  assign other_ops_83_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_83_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_83_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_83_I = I_84; // @[MapS.scala 20:41]
  assign other_ops_84_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_84_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_84_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_84_I = I_85; // @[MapS.scala 20:41]
  assign other_ops_85_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_85_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_85_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_85_I = I_86; // @[MapS.scala 20:41]
  assign other_ops_86_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_86_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_86_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_86_I = I_87; // @[MapS.scala 20:41]
  assign other_ops_87_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_87_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_87_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_87_I = I_88; // @[MapS.scala 20:41]
  assign other_ops_88_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_88_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_88_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_88_I = I_89; // @[MapS.scala 20:41]
  assign other_ops_89_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_89_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_89_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_89_I = I_90; // @[MapS.scala 20:41]
  assign other_ops_90_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_90_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_90_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_90_I = I_91; // @[MapS.scala 20:41]
  assign other_ops_91_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_91_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_91_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_91_I = I_92; // @[MapS.scala 20:41]
  assign other_ops_92_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_92_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_92_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_92_I = I_93; // @[MapS.scala 20:41]
  assign other_ops_93_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_93_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_93_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_93_I = I_94; // @[MapS.scala 20:41]
  assign other_ops_94_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_94_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_94_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_94_I = I_95; // @[MapS.scala 20:41]
  assign other_ops_95_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_95_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_95_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_95_I = I_96; // @[MapS.scala 20:41]
  assign other_ops_96_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_96_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_96_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_96_I = I_97; // @[MapS.scala 20:41]
  assign other_ops_97_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_97_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_97_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_97_I = I_98; // @[MapS.scala 20:41]
  assign other_ops_98_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_98_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_98_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_98_I = I_99; // @[MapS.scala 20:41]
  assign other_ops_99_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_99_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_99_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_99_I = I_100; // @[MapS.scala 20:41]
  assign other_ops_100_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_100_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_100_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_100_I = I_101; // @[MapS.scala 20:41]
  assign other_ops_101_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_101_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_101_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_101_I = I_102; // @[MapS.scala 20:41]
  assign other_ops_102_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_102_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_102_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_102_I = I_103; // @[MapS.scala 20:41]
  assign other_ops_103_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_103_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_103_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_103_I = I_104; // @[MapS.scala 20:41]
  assign other_ops_104_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_104_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_104_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_104_I = I_105; // @[MapS.scala 20:41]
  assign other_ops_105_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_105_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_105_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_105_I = I_106; // @[MapS.scala 20:41]
  assign other_ops_106_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_106_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_106_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_106_I = I_107; // @[MapS.scala 20:41]
  assign other_ops_107_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_107_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_107_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_107_I = I_108; // @[MapS.scala 20:41]
  assign other_ops_108_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_108_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_108_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_108_I = I_109; // @[MapS.scala 20:41]
  assign other_ops_109_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_109_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_109_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_109_I = I_110; // @[MapS.scala 20:41]
  assign other_ops_110_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_110_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_110_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_110_I = I_111; // @[MapS.scala 20:41]
  assign other_ops_111_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_111_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_111_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_111_I = I_112; // @[MapS.scala 20:41]
  assign other_ops_112_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_112_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_112_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_112_I = I_113; // @[MapS.scala 20:41]
  assign other_ops_113_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_113_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_113_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_113_I = I_114; // @[MapS.scala 20:41]
  assign other_ops_114_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_114_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_114_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_114_I = I_115; // @[MapS.scala 20:41]
  assign other_ops_115_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_115_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_115_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_115_I = I_116; // @[MapS.scala 20:41]
  assign other_ops_116_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_116_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_116_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_116_I = I_117; // @[MapS.scala 20:41]
  assign other_ops_117_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_117_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_117_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_117_I = I_118; // @[MapS.scala 20:41]
  assign other_ops_118_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_118_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_118_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_118_I = I_119; // @[MapS.scala 20:41]
  assign other_ops_119_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_119_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_119_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_119_I = I_120; // @[MapS.scala 20:41]
  assign other_ops_120_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_120_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_120_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_120_I = I_121; // @[MapS.scala 20:41]
  assign other_ops_121_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_121_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_121_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_121_I = I_122; // @[MapS.scala 20:41]
  assign other_ops_122_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_122_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_122_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_122_I = I_123; // @[MapS.scala 20:41]
  assign other_ops_123_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_123_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_123_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_123_I = I_124; // @[MapS.scala 20:41]
  assign other_ops_124_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_124_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_124_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_124_I = I_125; // @[MapS.scala 20:41]
  assign other_ops_125_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_125_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_125_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_125_I = I_126; // @[MapS.scala 20:41]
  assign other_ops_126_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_126_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_126_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_126_I = I_127; // @[MapS.scala 20:41]
  assign other_ops_127_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_127_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_127_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_127_I = I_128; // @[MapS.scala 20:41]
  assign other_ops_128_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_128_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_128_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_128_I = I_129; // @[MapS.scala 20:41]
  assign other_ops_129_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_129_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_129_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_129_I = I_130; // @[MapS.scala 20:41]
  assign other_ops_130_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_130_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_130_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_130_I = I_131; // @[MapS.scala 20:41]
  assign other_ops_131_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_131_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_131_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_131_I = I_132; // @[MapS.scala 20:41]
  assign other_ops_132_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_132_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_132_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_132_I = I_133; // @[MapS.scala 20:41]
  assign other_ops_133_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_133_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_133_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_133_I = I_134; // @[MapS.scala 20:41]
  assign other_ops_134_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_134_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_134_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_134_I = I_135; // @[MapS.scala 20:41]
  assign other_ops_135_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_135_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_135_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_135_I = I_136; // @[MapS.scala 20:41]
  assign other_ops_136_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_136_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_136_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_136_I = I_137; // @[MapS.scala 20:41]
  assign other_ops_137_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_137_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_137_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_137_I = I_138; // @[MapS.scala 20:41]
  assign other_ops_138_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_138_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_138_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_138_I = I_139; // @[MapS.scala 20:41]
  assign other_ops_139_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_139_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_139_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_139_I = I_140; // @[MapS.scala 20:41]
  assign other_ops_140_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_140_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_140_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_140_I = I_141; // @[MapS.scala 20:41]
  assign other_ops_141_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_141_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_141_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_141_I = I_142; // @[MapS.scala 20:41]
  assign other_ops_142_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_142_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_142_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_142_I = I_143; // @[MapS.scala 20:41]
  assign other_ops_143_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_143_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_143_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_143_I = I_144; // @[MapS.scala 20:41]
  assign other_ops_144_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_144_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_144_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_144_I = I_145; // @[MapS.scala 20:41]
  assign other_ops_145_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_145_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_145_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_145_I = I_146; // @[MapS.scala 20:41]
  assign other_ops_146_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_146_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_146_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_146_I = I_147; // @[MapS.scala 20:41]
  assign other_ops_147_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_147_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_147_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_147_I = I_148; // @[MapS.scala 20:41]
  assign other_ops_148_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_148_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_148_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_148_I = I_149; // @[MapS.scala 20:41]
  assign other_ops_149_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_149_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_149_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_149_I = I_150; // @[MapS.scala 20:41]
  assign other_ops_150_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_150_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_150_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_150_I = I_151; // @[MapS.scala 20:41]
  assign other_ops_151_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_151_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_151_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_151_I = I_152; // @[MapS.scala 20:41]
  assign other_ops_152_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_152_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_152_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_152_I = I_153; // @[MapS.scala 20:41]
  assign other_ops_153_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_153_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_153_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_153_I = I_154; // @[MapS.scala 20:41]
  assign other_ops_154_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_154_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_154_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_154_I = I_155; // @[MapS.scala 20:41]
  assign other_ops_155_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_155_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_155_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_155_I = I_156; // @[MapS.scala 20:41]
  assign other_ops_156_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_156_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_156_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_156_I = I_157; // @[MapS.scala 20:41]
  assign other_ops_157_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_157_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_157_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_157_I = I_158; // @[MapS.scala 20:41]
  assign other_ops_158_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_158_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_158_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_158_I = I_159; // @[MapS.scala 20:41]
  assign other_ops_159_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_159_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_159_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_159_I = I_160; // @[MapS.scala 20:41]
  assign other_ops_160_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_160_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_160_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_160_I = I_161; // @[MapS.scala 20:41]
  assign other_ops_161_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_161_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_161_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_161_I = I_162; // @[MapS.scala 20:41]
  assign other_ops_162_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_162_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_162_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_162_I = I_163; // @[MapS.scala 20:41]
  assign other_ops_163_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_163_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_163_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_163_I = I_164; // @[MapS.scala 20:41]
  assign other_ops_164_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_164_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_164_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_164_I = I_165; // @[MapS.scala 20:41]
  assign other_ops_165_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_165_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_165_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_165_I = I_166; // @[MapS.scala 20:41]
  assign other_ops_166_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_166_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_166_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_166_I = I_167; // @[MapS.scala 20:41]
  assign other_ops_167_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_167_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_167_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_167_I = I_168; // @[MapS.scala 20:41]
  assign other_ops_168_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_168_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_168_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_168_I = I_169; // @[MapS.scala 20:41]
  assign other_ops_169_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_169_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_169_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_169_I = I_170; // @[MapS.scala 20:41]
  assign other_ops_170_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_170_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_170_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_170_I = I_171; // @[MapS.scala 20:41]
  assign other_ops_171_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_171_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_171_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_171_I = I_172; // @[MapS.scala 20:41]
  assign other_ops_172_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_172_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_172_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_172_I = I_173; // @[MapS.scala 20:41]
  assign other_ops_173_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_173_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_173_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_173_I = I_174; // @[MapS.scala 20:41]
  assign other_ops_174_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_174_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_174_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_174_I = I_175; // @[MapS.scala 20:41]
  assign other_ops_175_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_175_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_175_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_175_I = I_176; // @[MapS.scala 20:41]
  assign other_ops_176_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_176_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_176_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_176_I = I_177; // @[MapS.scala 20:41]
  assign other_ops_177_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_177_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_177_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_177_I = I_178; // @[MapS.scala 20:41]
  assign other_ops_178_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_178_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_178_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_178_I = I_179; // @[MapS.scala 20:41]
  assign other_ops_179_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_179_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_179_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_179_I = I_180; // @[MapS.scala 20:41]
  assign other_ops_180_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_180_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_180_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_180_I = I_181; // @[MapS.scala 20:41]
  assign other_ops_181_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_181_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_181_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_181_I = I_182; // @[MapS.scala 20:41]
  assign other_ops_182_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_182_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_182_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_182_I = I_183; // @[MapS.scala 20:41]
  assign other_ops_183_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_183_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_183_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_183_I = I_184; // @[MapS.scala 20:41]
  assign other_ops_184_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_184_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_184_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_184_I = I_185; // @[MapS.scala 20:41]
  assign other_ops_185_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_185_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_185_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_185_I = I_186; // @[MapS.scala 20:41]
  assign other_ops_186_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_186_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_186_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_186_I = I_187; // @[MapS.scala 20:41]
  assign other_ops_187_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_187_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_187_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_187_I = I_188; // @[MapS.scala 20:41]
  assign other_ops_188_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_188_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_188_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_188_I = I_189; // @[MapS.scala 20:41]
  assign other_ops_189_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_189_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_189_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_189_I = I_190; // @[MapS.scala 20:41]
  assign other_ops_190_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_190_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_190_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_190_I = I_191; // @[MapS.scala 20:41]
  assign other_ops_191_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_191_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_191_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_191_I = I_192; // @[MapS.scala 20:41]
  assign other_ops_192_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_192_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_192_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_192_I = I_193; // @[MapS.scala 20:41]
  assign other_ops_193_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_193_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_193_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_193_I = I_194; // @[MapS.scala 20:41]
  assign other_ops_194_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_194_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_194_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_194_I = I_195; // @[MapS.scala 20:41]
  assign other_ops_195_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_195_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_195_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_195_I = I_196; // @[MapS.scala 20:41]
  assign other_ops_196_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_196_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_196_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_196_I = I_197; // @[MapS.scala 20:41]
  assign other_ops_197_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_197_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_197_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_197_I = I_198; // @[MapS.scala 20:41]
  assign other_ops_198_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_198_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_198_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_198_I = I_199; // @[MapS.scala 20:41]
endmodule
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  input  [7:0] I_4,
  input  [7:0] I_5,
  input  [7:0] I_6,
  input  [7:0] I_7,
  input  [7:0] I_8,
  input  [7:0] I_9,
  input  [7:0] I_10,
  input  [7:0] I_11,
  input  [7:0] I_12,
  input  [7:0] I_13,
  input  [7:0] I_14,
  input  [7:0] I_15,
  input  [7:0] I_16,
  input  [7:0] I_17,
  input  [7:0] I_18,
  input  [7:0] I_19,
  input  [7:0] I_20,
  input  [7:0] I_21,
  input  [7:0] I_22,
  input  [7:0] I_23,
  input  [7:0] I_24,
  input  [7:0] I_25,
  input  [7:0] I_26,
  input  [7:0] I_27,
  input  [7:0] I_28,
  input  [7:0] I_29,
  input  [7:0] I_30,
  input  [7:0] I_31,
  input  [7:0] I_32,
  input  [7:0] I_33,
  input  [7:0] I_34,
  input  [7:0] I_35,
  input  [7:0] I_36,
  input  [7:0] I_37,
  input  [7:0] I_38,
  input  [7:0] I_39,
  input  [7:0] I_40,
  input  [7:0] I_41,
  input  [7:0] I_42,
  input  [7:0] I_43,
  input  [7:0] I_44,
  input  [7:0] I_45,
  input  [7:0] I_46,
  input  [7:0] I_47,
  input  [7:0] I_48,
  input  [7:0] I_49,
  input  [7:0] I_50,
  input  [7:0] I_51,
  input  [7:0] I_52,
  input  [7:0] I_53,
  input  [7:0] I_54,
  input  [7:0] I_55,
  input  [7:0] I_56,
  input  [7:0] I_57,
  input  [7:0] I_58,
  input  [7:0] I_59,
  input  [7:0] I_60,
  input  [7:0] I_61,
  input  [7:0] I_62,
  input  [7:0] I_63,
  input  [7:0] I_64,
  input  [7:0] I_65,
  input  [7:0] I_66,
  input  [7:0] I_67,
  input  [7:0] I_68,
  input  [7:0] I_69,
  input  [7:0] I_70,
  input  [7:0] I_71,
  input  [7:0] I_72,
  input  [7:0] I_73,
  input  [7:0] I_74,
  input  [7:0] I_75,
  input  [7:0] I_76,
  input  [7:0] I_77,
  input  [7:0] I_78,
  input  [7:0] I_79,
  input  [7:0] I_80,
  input  [7:0] I_81,
  input  [7:0] I_82,
  input  [7:0] I_83,
  input  [7:0] I_84,
  input  [7:0] I_85,
  input  [7:0] I_86,
  input  [7:0] I_87,
  input  [7:0] I_88,
  input  [7:0] I_89,
  input  [7:0] I_90,
  input  [7:0] I_91,
  input  [7:0] I_92,
  input  [7:0] I_93,
  input  [7:0] I_94,
  input  [7:0] I_95,
  input  [7:0] I_96,
  input  [7:0] I_97,
  input  [7:0] I_98,
  input  [7:0] I_99,
  input  [7:0] I_100,
  input  [7:0] I_101,
  input  [7:0] I_102,
  input  [7:0] I_103,
  input  [7:0] I_104,
  input  [7:0] I_105,
  input  [7:0] I_106,
  input  [7:0] I_107,
  input  [7:0] I_108,
  input  [7:0] I_109,
  input  [7:0] I_110,
  input  [7:0] I_111,
  input  [7:0] I_112,
  input  [7:0] I_113,
  input  [7:0] I_114,
  input  [7:0] I_115,
  input  [7:0] I_116,
  input  [7:0] I_117,
  input  [7:0] I_118,
  input  [7:0] I_119,
  input  [7:0] I_120,
  input  [7:0] I_121,
  input  [7:0] I_122,
  input  [7:0] I_123,
  input  [7:0] I_124,
  input  [7:0] I_125,
  input  [7:0] I_126,
  input  [7:0] I_127,
  input  [7:0] I_128,
  input  [7:0] I_129,
  input  [7:0] I_130,
  input  [7:0] I_131,
  input  [7:0] I_132,
  input  [7:0] I_133,
  input  [7:0] I_134,
  input  [7:0] I_135,
  input  [7:0] I_136,
  input  [7:0] I_137,
  input  [7:0] I_138,
  input  [7:0] I_139,
  input  [7:0] I_140,
  input  [7:0] I_141,
  input  [7:0] I_142,
  input  [7:0] I_143,
  input  [7:0] I_144,
  input  [7:0] I_145,
  input  [7:0] I_146,
  input  [7:0] I_147,
  input  [7:0] I_148,
  input  [7:0] I_149,
  input  [7:0] I_150,
  input  [7:0] I_151,
  input  [7:0] I_152,
  input  [7:0] I_153,
  input  [7:0] I_154,
  input  [7:0] I_155,
  input  [7:0] I_156,
  input  [7:0] I_157,
  input  [7:0] I_158,
  input  [7:0] I_159,
  input  [7:0] I_160,
  input  [7:0] I_161,
  input  [7:0] I_162,
  input  [7:0] I_163,
  input  [7:0] I_164,
  input  [7:0] I_165,
  input  [7:0] I_166,
  input  [7:0] I_167,
  input  [7:0] I_168,
  input  [7:0] I_169,
  input  [7:0] I_170,
  input  [7:0] I_171,
  input  [7:0] I_172,
  input  [7:0] I_173,
  input  [7:0] I_174,
  input  [7:0] I_175,
  input  [7:0] I_176,
  input  [7:0] I_177,
  input  [7:0] I_178,
  input  [7:0] I_179,
  input  [7:0] I_180,
  input  [7:0] I_181,
  input  [7:0] I_182,
  input  [7:0] I_183,
  input  [7:0] I_184,
  input  [7:0] I_185,
  input  [7:0] I_186,
  input  [7:0] I_187,
  input  [7:0] I_188,
  input  [7:0] I_189,
  input  [7:0] I_190,
  input  [7:0] I_191,
  input  [7:0] I_192,
  input  [7:0] I_193,
  input  [7:0] I_194,
  input  [7:0] I_195,
  input  [7:0] I_196,
  input  [7:0] I_197,
  input  [7:0] I_198,
  input  [7:0] I_199,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15,
  output [7:0] O_16,
  output [7:0] O_17,
  output [7:0] O_18,
  output [7:0] O_19,
  output [7:0] O_20,
  output [7:0] O_21,
  output [7:0] O_22,
  output [7:0] O_23,
  output [7:0] O_24,
  output [7:0] O_25,
  output [7:0] O_26,
  output [7:0] O_27,
  output [7:0] O_28,
  output [7:0] O_29,
  output [7:0] O_30,
  output [7:0] O_31,
  output [7:0] O_32,
  output [7:0] O_33,
  output [7:0] O_34,
  output [7:0] O_35,
  output [7:0] O_36,
  output [7:0] O_37,
  output [7:0] O_38,
  output [7:0] O_39,
  output [7:0] O_40,
  output [7:0] O_41,
  output [7:0] O_42,
  output [7:0] O_43,
  output [7:0] O_44,
  output [7:0] O_45,
  output [7:0] O_46,
  output [7:0] O_47,
  output [7:0] O_48,
  output [7:0] O_49,
  output [7:0] O_50,
  output [7:0] O_51,
  output [7:0] O_52,
  output [7:0] O_53,
  output [7:0] O_54,
  output [7:0] O_55,
  output [7:0] O_56,
  output [7:0] O_57,
  output [7:0] O_58,
  output [7:0] O_59,
  output [7:0] O_60,
  output [7:0] O_61,
  output [7:0] O_62,
  output [7:0] O_63,
  output [7:0] O_64,
  output [7:0] O_65,
  output [7:0] O_66,
  output [7:0] O_67,
  output [7:0] O_68,
  output [7:0] O_69,
  output [7:0] O_70,
  output [7:0] O_71,
  output [7:0] O_72,
  output [7:0] O_73,
  output [7:0] O_74,
  output [7:0] O_75,
  output [7:0] O_76,
  output [7:0] O_77,
  output [7:0] O_78,
  output [7:0] O_79,
  output [7:0] O_80,
  output [7:0] O_81,
  output [7:0] O_82,
  output [7:0] O_83,
  output [7:0] O_84,
  output [7:0] O_85,
  output [7:0] O_86,
  output [7:0] O_87,
  output [7:0] O_88,
  output [7:0] O_89,
  output [7:0] O_90,
  output [7:0] O_91,
  output [7:0] O_92,
  output [7:0] O_93,
  output [7:0] O_94,
  output [7:0] O_95,
  output [7:0] O_96,
  output [7:0] O_97,
  output [7:0] O_98,
  output [7:0] O_99,
  output [7:0] O_100,
  output [7:0] O_101,
  output [7:0] O_102,
  output [7:0] O_103,
  output [7:0] O_104,
  output [7:0] O_105,
  output [7:0] O_106,
  output [7:0] O_107,
  output [7:0] O_108,
  output [7:0] O_109,
  output [7:0] O_110,
  output [7:0] O_111,
  output [7:0] O_112,
  output [7:0] O_113,
  output [7:0] O_114,
  output [7:0] O_115,
  output [7:0] O_116,
  output [7:0] O_117,
  output [7:0] O_118,
  output [7:0] O_119,
  output [7:0] O_120,
  output [7:0] O_121,
  output [7:0] O_122,
  output [7:0] O_123,
  output [7:0] O_124,
  output [7:0] O_125,
  output [7:0] O_126,
  output [7:0] O_127,
  output [7:0] O_128,
  output [7:0] O_129,
  output [7:0] O_130,
  output [7:0] O_131,
  output [7:0] O_132,
  output [7:0] O_133,
  output [7:0] O_134,
  output [7:0] O_135,
  output [7:0] O_136,
  output [7:0] O_137,
  output [7:0] O_138,
  output [7:0] O_139,
  output [7:0] O_140,
  output [7:0] O_141,
  output [7:0] O_142,
  output [7:0] O_143,
  output [7:0] O_144,
  output [7:0] O_145,
  output [7:0] O_146,
  output [7:0] O_147,
  output [7:0] O_148,
  output [7:0] O_149,
  output [7:0] O_150,
  output [7:0] O_151,
  output [7:0] O_152,
  output [7:0] O_153,
  output [7:0] O_154,
  output [7:0] O_155,
  output [7:0] O_156,
  output [7:0] O_157,
  output [7:0] O_158,
  output [7:0] O_159,
  output [7:0] O_160,
  output [7:0] O_161,
  output [7:0] O_162,
  output [7:0] O_163,
  output [7:0] O_164,
  output [7:0] O_165,
  output [7:0] O_166,
  output [7:0] O_167,
  output [7:0] O_168,
  output [7:0] O_169,
  output [7:0] O_170,
  output [7:0] O_171,
  output [7:0] O_172,
  output [7:0] O_173,
  output [7:0] O_174,
  output [7:0] O_175,
  output [7:0] O_176,
  output [7:0] O_177,
  output [7:0] O_178,
  output [7:0] O_179,
  output [7:0] O_180,
  output [7:0] O_181,
  output [7:0] O_182,
  output [7:0] O_183,
  output [7:0] O_184,
  output [7:0] O_185,
  output [7:0] O_186,
  output [7:0] O_187,
  output [7:0] O_188,
  output [7:0] O_189,
  output [7:0] O_190,
  output [7:0] O_191,
  output [7:0] O_192,
  output [7:0] O_193,
  output [7:0] O_194,
  output [7:0] O_195,
  output [7:0] O_196,
  output [7:0] O_197,
  output [7:0] O_198,
  output [7:0] O_199
);
  wire  n1_clock; // @[Top.scala 32:20]
  wire  n1_reset; // @[Top.scala 32:20]
  wire  n1_valid_up; // @[Top.scala 32:20]
  wire  n1_valid_down; // @[Top.scala 32:20]
  wire [7:0] n1_I_0; // @[Top.scala 32:20]
  wire [7:0] n1_I_1; // @[Top.scala 32:20]
  wire [7:0] n1_I_2; // @[Top.scala 32:20]
  wire [7:0] n1_I_3; // @[Top.scala 32:20]
  wire [7:0] n1_I_4; // @[Top.scala 32:20]
  wire [7:0] n1_I_5; // @[Top.scala 32:20]
  wire [7:0] n1_I_6; // @[Top.scala 32:20]
  wire [7:0] n1_I_7; // @[Top.scala 32:20]
  wire [7:0] n1_I_8; // @[Top.scala 32:20]
  wire [7:0] n1_I_9; // @[Top.scala 32:20]
  wire [7:0] n1_I_10; // @[Top.scala 32:20]
  wire [7:0] n1_I_11; // @[Top.scala 32:20]
  wire [7:0] n1_I_12; // @[Top.scala 32:20]
  wire [7:0] n1_I_13; // @[Top.scala 32:20]
  wire [7:0] n1_I_14; // @[Top.scala 32:20]
  wire [7:0] n1_I_15; // @[Top.scala 32:20]
  wire [7:0] n1_I_16; // @[Top.scala 32:20]
  wire [7:0] n1_I_17; // @[Top.scala 32:20]
  wire [7:0] n1_I_18; // @[Top.scala 32:20]
  wire [7:0] n1_I_19; // @[Top.scala 32:20]
  wire [7:0] n1_I_20; // @[Top.scala 32:20]
  wire [7:0] n1_I_21; // @[Top.scala 32:20]
  wire [7:0] n1_I_22; // @[Top.scala 32:20]
  wire [7:0] n1_I_23; // @[Top.scala 32:20]
  wire [7:0] n1_I_24; // @[Top.scala 32:20]
  wire [7:0] n1_I_25; // @[Top.scala 32:20]
  wire [7:0] n1_I_26; // @[Top.scala 32:20]
  wire [7:0] n1_I_27; // @[Top.scala 32:20]
  wire [7:0] n1_I_28; // @[Top.scala 32:20]
  wire [7:0] n1_I_29; // @[Top.scala 32:20]
  wire [7:0] n1_I_30; // @[Top.scala 32:20]
  wire [7:0] n1_I_31; // @[Top.scala 32:20]
  wire [7:0] n1_I_32; // @[Top.scala 32:20]
  wire [7:0] n1_I_33; // @[Top.scala 32:20]
  wire [7:0] n1_I_34; // @[Top.scala 32:20]
  wire [7:0] n1_I_35; // @[Top.scala 32:20]
  wire [7:0] n1_I_36; // @[Top.scala 32:20]
  wire [7:0] n1_I_37; // @[Top.scala 32:20]
  wire [7:0] n1_I_38; // @[Top.scala 32:20]
  wire [7:0] n1_I_39; // @[Top.scala 32:20]
  wire [7:0] n1_I_40; // @[Top.scala 32:20]
  wire [7:0] n1_I_41; // @[Top.scala 32:20]
  wire [7:0] n1_I_42; // @[Top.scala 32:20]
  wire [7:0] n1_I_43; // @[Top.scala 32:20]
  wire [7:0] n1_I_44; // @[Top.scala 32:20]
  wire [7:0] n1_I_45; // @[Top.scala 32:20]
  wire [7:0] n1_I_46; // @[Top.scala 32:20]
  wire [7:0] n1_I_47; // @[Top.scala 32:20]
  wire [7:0] n1_I_48; // @[Top.scala 32:20]
  wire [7:0] n1_I_49; // @[Top.scala 32:20]
  wire [7:0] n1_I_50; // @[Top.scala 32:20]
  wire [7:0] n1_I_51; // @[Top.scala 32:20]
  wire [7:0] n1_I_52; // @[Top.scala 32:20]
  wire [7:0] n1_I_53; // @[Top.scala 32:20]
  wire [7:0] n1_I_54; // @[Top.scala 32:20]
  wire [7:0] n1_I_55; // @[Top.scala 32:20]
  wire [7:0] n1_I_56; // @[Top.scala 32:20]
  wire [7:0] n1_I_57; // @[Top.scala 32:20]
  wire [7:0] n1_I_58; // @[Top.scala 32:20]
  wire [7:0] n1_I_59; // @[Top.scala 32:20]
  wire [7:0] n1_I_60; // @[Top.scala 32:20]
  wire [7:0] n1_I_61; // @[Top.scala 32:20]
  wire [7:0] n1_I_62; // @[Top.scala 32:20]
  wire [7:0] n1_I_63; // @[Top.scala 32:20]
  wire [7:0] n1_I_64; // @[Top.scala 32:20]
  wire [7:0] n1_I_65; // @[Top.scala 32:20]
  wire [7:0] n1_I_66; // @[Top.scala 32:20]
  wire [7:0] n1_I_67; // @[Top.scala 32:20]
  wire [7:0] n1_I_68; // @[Top.scala 32:20]
  wire [7:0] n1_I_69; // @[Top.scala 32:20]
  wire [7:0] n1_I_70; // @[Top.scala 32:20]
  wire [7:0] n1_I_71; // @[Top.scala 32:20]
  wire [7:0] n1_I_72; // @[Top.scala 32:20]
  wire [7:0] n1_I_73; // @[Top.scala 32:20]
  wire [7:0] n1_I_74; // @[Top.scala 32:20]
  wire [7:0] n1_I_75; // @[Top.scala 32:20]
  wire [7:0] n1_I_76; // @[Top.scala 32:20]
  wire [7:0] n1_I_77; // @[Top.scala 32:20]
  wire [7:0] n1_I_78; // @[Top.scala 32:20]
  wire [7:0] n1_I_79; // @[Top.scala 32:20]
  wire [7:0] n1_I_80; // @[Top.scala 32:20]
  wire [7:0] n1_I_81; // @[Top.scala 32:20]
  wire [7:0] n1_I_82; // @[Top.scala 32:20]
  wire [7:0] n1_I_83; // @[Top.scala 32:20]
  wire [7:0] n1_I_84; // @[Top.scala 32:20]
  wire [7:0] n1_I_85; // @[Top.scala 32:20]
  wire [7:0] n1_I_86; // @[Top.scala 32:20]
  wire [7:0] n1_I_87; // @[Top.scala 32:20]
  wire [7:0] n1_I_88; // @[Top.scala 32:20]
  wire [7:0] n1_I_89; // @[Top.scala 32:20]
  wire [7:0] n1_I_90; // @[Top.scala 32:20]
  wire [7:0] n1_I_91; // @[Top.scala 32:20]
  wire [7:0] n1_I_92; // @[Top.scala 32:20]
  wire [7:0] n1_I_93; // @[Top.scala 32:20]
  wire [7:0] n1_I_94; // @[Top.scala 32:20]
  wire [7:0] n1_I_95; // @[Top.scala 32:20]
  wire [7:0] n1_I_96; // @[Top.scala 32:20]
  wire [7:0] n1_I_97; // @[Top.scala 32:20]
  wire [7:0] n1_I_98; // @[Top.scala 32:20]
  wire [7:0] n1_I_99; // @[Top.scala 32:20]
  wire [7:0] n1_I_100; // @[Top.scala 32:20]
  wire [7:0] n1_I_101; // @[Top.scala 32:20]
  wire [7:0] n1_I_102; // @[Top.scala 32:20]
  wire [7:0] n1_I_103; // @[Top.scala 32:20]
  wire [7:0] n1_I_104; // @[Top.scala 32:20]
  wire [7:0] n1_I_105; // @[Top.scala 32:20]
  wire [7:0] n1_I_106; // @[Top.scala 32:20]
  wire [7:0] n1_I_107; // @[Top.scala 32:20]
  wire [7:0] n1_I_108; // @[Top.scala 32:20]
  wire [7:0] n1_I_109; // @[Top.scala 32:20]
  wire [7:0] n1_I_110; // @[Top.scala 32:20]
  wire [7:0] n1_I_111; // @[Top.scala 32:20]
  wire [7:0] n1_I_112; // @[Top.scala 32:20]
  wire [7:0] n1_I_113; // @[Top.scala 32:20]
  wire [7:0] n1_I_114; // @[Top.scala 32:20]
  wire [7:0] n1_I_115; // @[Top.scala 32:20]
  wire [7:0] n1_I_116; // @[Top.scala 32:20]
  wire [7:0] n1_I_117; // @[Top.scala 32:20]
  wire [7:0] n1_I_118; // @[Top.scala 32:20]
  wire [7:0] n1_I_119; // @[Top.scala 32:20]
  wire [7:0] n1_I_120; // @[Top.scala 32:20]
  wire [7:0] n1_I_121; // @[Top.scala 32:20]
  wire [7:0] n1_I_122; // @[Top.scala 32:20]
  wire [7:0] n1_I_123; // @[Top.scala 32:20]
  wire [7:0] n1_I_124; // @[Top.scala 32:20]
  wire [7:0] n1_I_125; // @[Top.scala 32:20]
  wire [7:0] n1_I_126; // @[Top.scala 32:20]
  wire [7:0] n1_I_127; // @[Top.scala 32:20]
  wire [7:0] n1_I_128; // @[Top.scala 32:20]
  wire [7:0] n1_I_129; // @[Top.scala 32:20]
  wire [7:0] n1_I_130; // @[Top.scala 32:20]
  wire [7:0] n1_I_131; // @[Top.scala 32:20]
  wire [7:0] n1_I_132; // @[Top.scala 32:20]
  wire [7:0] n1_I_133; // @[Top.scala 32:20]
  wire [7:0] n1_I_134; // @[Top.scala 32:20]
  wire [7:0] n1_I_135; // @[Top.scala 32:20]
  wire [7:0] n1_I_136; // @[Top.scala 32:20]
  wire [7:0] n1_I_137; // @[Top.scala 32:20]
  wire [7:0] n1_I_138; // @[Top.scala 32:20]
  wire [7:0] n1_I_139; // @[Top.scala 32:20]
  wire [7:0] n1_I_140; // @[Top.scala 32:20]
  wire [7:0] n1_I_141; // @[Top.scala 32:20]
  wire [7:0] n1_I_142; // @[Top.scala 32:20]
  wire [7:0] n1_I_143; // @[Top.scala 32:20]
  wire [7:0] n1_I_144; // @[Top.scala 32:20]
  wire [7:0] n1_I_145; // @[Top.scala 32:20]
  wire [7:0] n1_I_146; // @[Top.scala 32:20]
  wire [7:0] n1_I_147; // @[Top.scala 32:20]
  wire [7:0] n1_I_148; // @[Top.scala 32:20]
  wire [7:0] n1_I_149; // @[Top.scala 32:20]
  wire [7:0] n1_I_150; // @[Top.scala 32:20]
  wire [7:0] n1_I_151; // @[Top.scala 32:20]
  wire [7:0] n1_I_152; // @[Top.scala 32:20]
  wire [7:0] n1_I_153; // @[Top.scala 32:20]
  wire [7:0] n1_I_154; // @[Top.scala 32:20]
  wire [7:0] n1_I_155; // @[Top.scala 32:20]
  wire [7:0] n1_I_156; // @[Top.scala 32:20]
  wire [7:0] n1_I_157; // @[Top.scala 32:20]
  wire [7:0] n1_I_158; // @[Top.scala 32:20]
  wire [7:0] n1_I_159; // @[Top.scala 32:20]
  wire [7:0] n1_I_160; // @[Top.scala 32:20]
  wire [7:0] n1_I_161; // @[Top.scala 32:20]
  wire [7:0] n1_I_162; // @[Top.scala 32:20]
  wire [7:0] n1_I_163; // @[Top.scala 32:20]
  wire [7:0] n1_I_164; // @[Top.scala 32:20]
  wire [7:0] n1_I_165; // @[Top.scala 32:20]
  wire [7:0] n1_I_166; // @[Top.scala 32:20]
  wire [7:0] n1_I_167; // @[Top.scala 32:20]
  wire [7:0] n1_I_168; // @[Top.scala 32:20]
  wire [7:0] n1_I_169; // @[Top.scala 32:20]
  wire [7:0] n1_I_170; // @[Top.scala 32:20]
  wire [7:0] n1_I_171; // @[Top.scala 32:20]
  wire [7:0] n1_I_172; // @[Top.scala 32:20]
  wire [7:0] n1_I_173; // @[Top.scala 32:20]
  wire [7:0] n1_I_174; // @[Top.scala 32:20]
  wire [7:0] n1_I_175; // @[Top.scala 32:20]
  wire [7:0] n1_I_176; // @[Top.scala 32:20]
  wire [7:0] n1_I_177; // @[Top.scala 32:20]
  wire [7:0] n1_I_178; // @[Top.scala 32:20]
  wire [7:0] n1_I_179; // @[Top.scala 32:20]
  wire [7:0] n1_I_180; // @[Top.scala 32:20]
  wire [7:0] n1_I_181; // @[Top.scala 32:20]
  wire [7:0] n1_I_182; // @[Top.scala 32:20]
  wire [7:0] n1_I_183; // @[Top.scala 32:20]
  wire [7:0] n1_I_184; // @[Top.scala 32:20]
  wire [7:0] n1_I_185; // @[Top.scala 32:20]
  wire [7:0] n1_I_186; // @[Top.scala 32:20]
  wire [7:0] n1_I_187; // @[Top.scala 32:20]
  wire [7:0] n1_I_188; // @[Top.scala 32:20]
  wire [7:0] n1_I_189; // @[Top.scala 32:20]
  wire [7:0] n1_I_190; // @[Top.scala 32:20]
  wire [7:0] n1_I_191; // @[Top.scala 32:20]
  wire [7:0] n1_I_192; // @[Top.scala 32:20]
  wire [7:0] n1_I_193; // @[Top.scala 32:20]
  wire [7:0] n1_I_194; // @[Top.scala 32:20]
  wire [7:0] n1_I_195; // @[Top.scala 32:20]
  wire [7:0] n1_I_196; // @[Top.scala 32:20]
  wire [7:0] n1_I_197; // @[Top.scala 32:20]
  wire [7:0] n1_I_198; // @[Top.scala 32:20]
  wire [7:0] n1_I_199; // @[Top.scala 32:20]
  wire [7:0] n1_O_0; // @[Top.scala 32:20]
  wire [7:0] n1_O_1; // @[Top.scala 32:20]
  wire [7:0] n1_O_2; // @[Top.scala 32:20]
  wire [7:0] n1_O_3; // @[Top.scala 32:20]
  wire [7:0] n1_O_4; // @[Top.scala 32:20]
  wire [7:0] n1_O_5; // @[Top.scala 32:20]
  wire [7:0] n1_O_6; // @[Top.scala 32:20]
  wire [7:0] n1_O_7; // @[Top.scala 32:20]
  wire [7:0] n1_O_8; // @[Top.scala 32:20]
  wire [7:0] n1_O_9; // @[Top.scala 32:20]
  wire [7:0] n1_O_10; // @[Top.scala 32:20]
  wire [7:0] n1_O_11; // @[Top.scala 32:20]
  wire [7:0] n1_O_12; // @[Top.scala 32:20]
  wire [7:0] n1_O_13; // @[Top.scala 32:20]
  wire [7:0] n1_O_14; // @[Top.scala 32:20]
  wire [7:0] n1_O_15; // @[Top.scala 32:20]
  wire [7:0] n1_O_16; // @[Top.scala 32:20]
  wire [7:0] n1_O_17; // @[Top.scala 32:20]
  wire [7:0] n1_O_18; // @[Top.scala 32:20]
  wire [7:0] n1_O_19; // @[Top.scala 32:20]
  wire [7:0] n1_O_20; // @[Top.scala 32:20]
  wire [7:0] n1_O_21; // @[Top.scala 32:20]
  wire [7:0] n1_O_22; // @[Top.scala 32:20]
  wire [7:0] n1_O_23; // @[Top.scala 32:20]
  wire [7:0] n1_O_24; // @[Top.scala 32:20]
  wire [7:0] n1_O_25; // @[Top.scala 32:20]
  wire [7:0] n1_O_26; // @[Top.scala 32:20]
  wire [7:0] n1_O_27; // @[Top.scala 32:20]
  wire [7:0] n1_O_28; // @[Top.scala 32:20]
  wire [7:0] n1_O_29; // @[Top.scala 32:20]
  wire [7:0] n1_O_30; // @[Top.scala 32:20]
  wire [7:0] n1_O_31; // @[Top.scala 32:20]
  wire [7:0] n1_O_32; // @[Top.scala 32:20]
  wire [7:0] n1_O_33; // @[Top.scala 32:20]
  wire [7:0] n1_O_34; // @[Top.scala 32:20]
  wire [7:0] n1_O_35; // @[Top.scala 32:20]
  wire [7:0] n1_O_36; // @[Top.scala 32:20]
  wire [7:0] n1_O_37; // @[Top.scala 32:20]
  wire [7:0] n1_O_38; // @[Top.scala 32:20]
  wire [7:0] n1_O_39; // @[Top.scala 32:20]
  wire [7:0] n1_O_40; // @[Top.scala 32:20]
  wire [7:0] n1_O_41; // @[Top.scala 32:20]
  wire [7:0] n1_O_42; // @[Top.scala 32:20]
  wire [7:0] n1_O_43; // @[Top.scala 32:20]
  wire [7:0] n1_O_44; // @[Top.scala 32:20]
  wire [7:0] n1_O_45; // @[Top.scala 32:20]
  wire [7:0] n1_O_46; // @[Top.scala 32:20]
  wire [7:0] n1_O_47; // @[Top.scala 32:20]
  wire [7:0] n1_O_48; // @[Top.scala 32:20]
  wire [7:0] n1_O_49; // @[Top.scala 32:20]
  wire [7:0] n1_O_50; // @[Top.scala 32:20]
  wire [7:0] n1_O_51; // @[Top.scala 32:20]
  wire [7:0] n1_O_52; // @[Top.scala 32:20]
  wire [7:0] n1_O_53; // @[Top.scala 32:20]
  wire [7:0] n1_O_54; // @[Top.scala 32:20]
  wire [7:0] n1_O_55; // @[Top.scala 32:20]
  wire [7:0] n1_O_56; // @[Top.scala 32:20]
  wire [7:0] n1_O_57; // @[Top.scala 32:20]
  wire [7:0] n1_O_58; // @[Top.scala 32:20]
  wire [7:0] n1_O_59; // @[Top.scala 32:20]
  wire [7:0] n1_O_60; // @[Top.scala 32:20]
  wire [7:0] n1_O_61; // @[Top.scala 32:20]
  wire [7:0] n1_O_62; // @[Top.scala 32:20]
  wire [7:0] n1_O_63; // @[Top.scala 32:20]
  wire [7:0] n1_O_64; // @[Top.scala 32:20]
  wire [7:0] n1_O_65; // @[Top.scala 32:20]
  wire [7:0] n1_O_66; // @[Top.scala 32:20]
  wire [7:0] n1_O_67; // @[Top.scala 32:20]
  wire [7:0] n1_O_68; // @[Top.scala 32:20]
  wire [7:0] n1_O_69; // @[Top.scala 32:20]
  wire [7:0] n1_O_70; // @[Top.scala 32:20]
  wire [7:0] n1_O_71; // @[Top.scala 32:20]
  wire [7:0] n1_O_72; // @[Top.scala 32:20]
  wire [7:0] n1_O_73; // @[Top.scala 32:20]
  wire [7:0] n1_O_74; // @[Top.scala 32:20]
  wire [7:0] n1_O_75; // @[Top.scala 32:20]
  wire [7:0] n1_O_76; // @[Top.scala 32:20]
  wire [7:0] n1_O_77; // @[Top.scala 32:20]
  wire [7:0] n1_O_78; // @[Top.scala 32:20]
  wire [7:0] n1_O_79; // @[Top.scala 32:20]
  wire [7:0] n1_O_80; // @[Top.scala 32:20]
  wire [7:0] n1_O_81; // @[Top.scala 32:20]
  wire [7:0] n1_O_82; // @[Top.scala 32:20]
  wire [7:0] n1_O_83; // @[Top.scala 32:20]
  wire [7:0] n1_O_84; // @[Top.scala 32:20]
  wire [7:0] n1_O_85; // @[Top.scala 32:20]
  wire [7:0] n1_O_86; // @[Top.scala 32:20]
  wire [7:0] n1_O_87; // @[Top.scala 32:20]
  wire [7:0] n1_O_88; // @[Top.scala 32:20]
  wire [7:0] n1_O_89; // @[Top.scala 32:20]
  wire [7:0] n1_O_90; // @[Top.scala 32:20]
  wire [7:0] n1_O_91; // @[Top.scala 32:20]
  wire [7:0] n1_O_92; // @[Top.scala 32:20]
  wire [7:0] n1_O_93; // @[Top.scala 32:20]
  wire [7:0] n1_O_94; // @[Top.scala 32:20]
  wire [7:0] n1_O_95; // @[Top.scala 32:20]
  wire [7:0] n1_O_96; // @[Top.scala 32:20]
  wire [7:0] n1_O_97; // @[Top.scala 32:20]
  wire [7:0] n1_O_98; // @[Top.scala 32:20]
  wire [7:0] n1_O_99; // @[Top.scala 32:20]
  wire [7:0] n1_O_100; // @[Top.scala 32:20]
  wire [7:0] n1_O_101; // @[Top.scala 32:20]
  wire [7:0] n1_O_102; // @[Top.scala 32:20]
  wire [7:0] n1_O_103; // @[Top.scala 32:20]
  wire [7:0] n1_O_104; // @[Top.scala 32:20]
  wire [7:0] n1_O_105; // @[Top.scala 32:20]
  wire [7:0] n1_O_106; // @[Top.scala 32:20]
  wire [7:0] n1_O_107; // @[Top.scala 32:20]
  wire [7:0] n1_O_108; // @[Top.scala 32:20]
  wire [7:0] n1_O_109; // @[Top.scala 32:20]
  wire [7:0] n1_O_110; // @[Top.scala 32:20]
  wire [7:0] n1_O_111; // @[Top.scala 32:20]
  wire [7:0] n1_O_112; // @[Top.scala 32:20]
  wire [7:0] n1_O_113; // @[Top.scala 32:20]
  wire [7:0] n1_O_114; // @[Top.scala 32:20]
  wire [7:0] n1_O_115; // @[Top.scala 32:20]
  wire [7:0] n1_O_116; // @[Top.scala 32:20]
  wire [7:0] n1_O_117; // @[Top.scala 32:20]
  wire [7:0] n1_O_118; // @[Top.scala 32:20]
  wire [7:0] n1_O_119; // @[Top.scala 32:20]
  wire [7:0] n1_O_120; // @[Top.scala 32:20]
  wire [7:0] n1_O_121; // @[Top.scala 32:20]
  wire [7:0] n1_O_122; // @[Top.scala 32:20]
  wire [7:0] n1_O_123; // @[Top.scala 32:20]
  wire [7:0] n1_O_124; // @[Top.scala 32:20]
  wire [7:0] n1_O_125; // @[Top.scala 32:20]
  wire [7:0] n1_O_126; // @[Top.scala 32:20]
  wire [7:0] n1_O_127; // @[Top.scala 32:20]
  wire [7:0] n1_O_128; // @[Top.scala 32:20]
  wire [7:0] n1_O_129; // @[Top.scala 32:20]
  wire [7:0] n1_O_130; // @[Top.scala 32:20]
  wire [7:0] n1_O_131; // @[Top.scala 32:20]
  wire [7:0] n1_O_132; // @[Top.scala 32:20]
  wire [7:0] n1_O_133; // @[Top.scala 32:20]
  wire [7:0] n1_O_134; // @[Top.scala 32:20]
  wire [7:0] n1_O_135; // @[Top.scala 32:20]
  wire [7:0] n1_O_136; // @[Top.scala 32:20]
  wire [7:0] n1_O_137; // @[Top.scala 32:20]
  wire [7:0] n1_O_138; // @[Top.scala 32:20]
  wire [7:0] n1_O_139; // @[Top.scala 32:20]
  wire [7:0] n1_O_140; // @[Top.scala 32:20]
  wire [7:0] n1_O_141; // @[Top.scala 32:20]
  wire [7:0] n1_O_142; // @[Top.scala 32:20]
  wire [7:0] n1_O_143; // @[Top.scala 32:20]
  wire [7:0] n1_O_144; // @[Top.scala 32:20]
  wire [7:0] n1_O_145; // @[Top.scala 32:20]
  wire [7:0] n1_O_146; // @[Top.scala 32:20]
  wire [7:0] n1_O_147; // @[Top.scala 32:20]
  wire [7:0] n1_O_148; // @[Top.scala 32:20]
  wire [7:0] n1_O_149; // @[Top.scala 32:20]
  wire [7:0] n1_O_150; // @[Top.scala 32:20]
  wire [7:0] n1_O_151; // @[Top.scala 32:20]
  wire [7:0] n1_O_152; // @[Top.scala 32:20]
  wire [7:0] n1_O_153; // @[Top.scala 32:20]
  wire [7:0] n1_O_154; // @[Top.scala 32:20]
  wire [7:0] n1_O_155; // @[Top.scala 32:20]
  wire [7:0] n1_O_156; // @[Top.scala 32:20]
  wire [7:0] n1_O_157; // @[Top.scala 32:20]
  wire [7:0] n1_O_158; // @[Top.scala 32:20]
  wire [7:0] n1_O_159; // @[Top.scala 32:20]
  wire [7:0] n1_O_160; // @[Top.scala 32:20]
  wire [7:0] n1_O_161; // @[Top.scala 32:20]
  wire [7:0] n1_O_162; // @[Top.scala 32:20]
  wire [7:0] n1_O_163; // @[Top.scala 32:20]
  wire [7:0] n1_O_164; // @[Top.scala 32:20]
  wire [7:0] n1_O_165; // @[Top.scala 32:20]
  wire [7:0] n1_O_166; // @[Top.scala 32:20]
  wire [7:0] n1_O_167; // @[Top.scala 32:20]
  wire [7:0] n1_O_168; // @[Top.scala 32:20]
  wire [7:0] n1_O_169; // @[Top.scala 32:20]
  wire [7:0] n1_O_170; // @[Top.scala 32:20]
  wire [7:0] n1_O_171; // @[Top.scala 32:20]
  wire [7:0] n1_O_172; // @[Top.scala 32:20]
  wire [7:0] n1_O_173; // @[Top.scala 32:20]
  wire [7:0] n1_O_174; // @[Top.scala 32:20]
  wire [7:0] n1_O_175; // @[Top.scala 32:20]
  wire [7:0] n1_O_176; // @[Top.scala 32:20]
  wire [7:0] n1_O_177; // @[Top.scala 32:20]
  wire [7:0] n1_O_178; // @[Top.scala 32:20]
  wire [7:0] n1_O_179; // @[Top.scala 32:20]
  wire [7:0] n1_O_180; // @[Top.scala 32:20]
  wire [7:0] n1_O_181; // @[Top.scala 32:20]
  wire [7:0] n1_O_182; // @[Top.scala 32:20]
  wire [7:0] n1_O_183; // @[Top.scala 32:20]
  wire [7:0] n1_O_184; // @[Top.scala 32:20]
  wire [7:0] n1_O_185; // @[Top.scala 32:20]
  wire [7:0] n1_O_186; // @[Top.scala 32:20]
  wire [7:0] n1_O_187; // @[Top.scala 32:20]
  wire [7:0] n1_O_188; // @[Top.scala 32:20]
  wire [7:0] n1_O_189; // @[Top.scala 32:20]
  wire [7:0] n1_O_190; // @[Top.scala 32:20]
  wire [7:0] n1_O_191; // @[Top.scala 32:20]
  wire [7:0] n1_O_192; // @[Top.scala 32:20]
  wire [7:0] n1_O_193; // @[Top.scala 32:20]
  wire [7:0] n1_O_194; // @[Top.scala 32:20]
  wire [7:0] n1_O_195; // @[Top.scala 32:20]
  wire [7:0] n1_O_196; // @[Top.scala 32:20]
  wire [7:0] n1_O_197; // @[Top.scala 32:20]
  wire [7:0] n1_O_198; // @[Top.scala 32:20]
  wire [7:0] n1_O_199; // @[Top.scala 32:20]
  wire  n7_clock; // @[Top.scala 35:20]
  wire  n7_reset; // @[Top.scala 35:20]
  wire  n7_valid_up; // @[Top.scala 35:20]
  wire  n7_valid_down; // @[Top.scala 35:20]
  wire [7:0] n7_I_0; // @[Top.scala 35:20]
  wire [7:0] n7_I_1; // @[Top.scala 35:20]
  wire [7:0] n7_I_2; // @[Top.scala 35:20]
  wire [7:0] n7_I_3; // @[Top.scala 35:20]
  wire [7:0] n7_I_4; // @[Top.scala 35:20]
  wire [7:0] n7_I_5; // @[Top.scala 35:20]
  wire [7:0] n7_I_6; // @[Top.scala 35:20]
  wire [7:0] n7_I_7; // @[Top.scala 35:20]
  wire [7:0] n7_I_8; // @[Top.scala 35:20]
  wire [7:0] n7_I_9; // @[Top.scala 35:20]
  wire [7:0] n7_I_10; // @[Top.scala 35:20]
  wire [7:0] n7_I_11; // @[Top.scala 35:20]
  wire [7:0] n7_I_12; // @[Top.scala 35:20]
  wire [7:0] n7_I_13; // @[Top.scala 35:20]
  wire [7:0] n7_I_14; // @[Top.scala 35:20]
  wire [7:0] n7_I_15; // @[Top.scala 35:20]
  wire [7:0] n7_I_16; // @[Top.scala 35:20]
  wire [7:0] n7_I_17; // @[Top.scala 35:20]
  wire [7:0] n7_I_18; // @[Top.scala 35:20]
  wire [7:0] n7_I_19; // @[Top.scala 35:20]
  wire [7:0] n7_I_20; // @[Top.scala 35:20]
  wire [7:0] n7_I_21; // @[Top.scala 35:20]
  wire [7:0] n7_I_22; // @[Top.scala 35:20]
  wire [7:0] n7_I_23; // @[Top.scala 35:20]
  wire [7:0] n7_I_24; // @[Top.scala 35:20]
  wire [7:0] n7_I_25; // @[Top.scala 35:20]
  wire [7:0] n7_I_26; // @[Top.scala 35:20]
  wire [7:0] n7_I_27; // @[Top.scala 35:20]
  wire [7:0] n7_I_28; // @[Top.scala 35:20]
  wire [7:0] n7_I_29; // @[Top.scala 35:20]
  wire [7:0] n7_I_30; // @[Top.scala 35:20]
  wire [7:0] n7_I_31; // @[Top.scala 35:20]
  wire [7:0] n7_I_32; // @[Top.scala 35:20]
  wire [7:0] n7_I_33; // @[Top.scala 35:20]
  wire [7:0] n7_I_34; // @[Top.scala 35:20]
  wire [7:0] n7_I_35; // @[Top.scala 35:20]
  wire [7:0] n7_I_36; // @[Top.scala 35:20]
  wire [7:0] n7_I_37; // @[Top.scala 35:20]
  wire [7:0] n7_I_38; // @[Top.scala 35:20]
  wire [7:0] n7_I_39; // @[Top.scala 35:20]
  wire [7:0] n7_I_40; // @[Top.scala 35:20]
  wire [7:0] n7_I_41; // @[Top.scala 35:20]
  wire [7:0] n7_I_42; // @[Top.scala 35:20]
  wire [7:0] n7_I_43; // @[Top.scala 35:20]
  wire [7:0] n7_I_44; // @[Top.scala 35:20]
  wire [7:0] n7_I_45; // @[Top.scala 35:20]
  wire [7:0] n7_I_46; // @[Top.scala 35:20]
  wire [7:0] n7_I_47; // @[Top.scala 35:20]
  wire [7:0] n7_I_48; // @[Top.scala 35:20]
  wire [7:0] n7_I_49; // @[Top.scala 35:20]
  wire [7:0] n7_I_50; // @[Top.scala 35:20]
  wire [7:0] n7_I_51; // @[Top.scala 35:20]
  wire [7:0] n7_I_52; // @[Top.scala 35:20]
  wire [7:0] n7_I_53; // @[Top.scala 35:20]
  wire [7:0] n7_I_54; // @[Top.scala 35:20]
  wire [7:0] n7_I_55; // @[Top.scala 35:20]
  wire [7:0] n7_I_56; // @[Top.scala 35:20]
  wire [7:0] n7_I_57; // @[Top.scala 35:20]
  wire [7:0] n7_I_58; // @[Top.scala 35:20]
  wire [7:0] n7_I_59; // @[Top.scala 35:20]
  wire [7:0] n7_I_60; // @[Top.scala 35:20]
  wire [7:0] n7_I_61; // @[Top.scala 35:20]
  wire [7:0] n7_I_62; // @[Top.scala 35:20]
  wire [7:0] n7_I_63; // @[Top.scala 35:20]
  wire [7:0] n7_I_64; // @[Top.scala 35:20]
  wire [7:0] n7_I_65; // @[Top.scala 35:20]
  wire [7:0] n7_I_66; // @[Top.scala 35:20]
  wire [7:0] n7_I_67; // @[Top.scala 35:20]
  wire [7:0] n7_I_68; // @[Top.scala 35:20]
  wire [7:0] n7_I_69; // @[Top.scala 35:20]
  wire [7:0] n7_I_70; // @[Top.scala 35:20]
  wire [7:0] n7_I_71; // @[Top.scala 35:20]
  wire [7:0] n7_I_72; // @[Top.scala 35:20]
  wire [7:0] n7_I_73; // @[Top.scala 35:20]
  wire [7:0] n7_I_74; // @[Top.scala 35:20]
  wire [7:0] n7_I_75; // @[Top.scala 35:20]
  wire [7:0] n7_I_76; // @[Top.scala 35:20]
  wire [7:0] n7_I_77; // @[Top.scala 35:20]
  wire [7:0] n7_I_78; // @[Top.scala 35:20]
  wire [7:0] n7_I_79; // @[Top.scala 35:20]
  wire [7:0] n7_I_80; // @[Top.scala 35:20]
  wire [7:0] n7_I_81; // @[Top.scala 35:20]
  wire [7:0] n7_I_82; // @[Top.scala 35:20]
  wire [7:0] n7_I_83; // @[Top.scala 35:20]
  wire [7:0] n7_I_84; // @[Top.scala 35:20]
  wire [7:0] n7_I_85; // @[Top.scala 35:20]
  wire [7:0] n7_I_86; // @[Top.scala 35:20]
  wire [7:0] n7_I_87; // @[Top.scala 35:20]
  wire [7:0] n7_I_88; // @[Top.scala 35:20]
  wire [7:0] n7_I_89; // @[Top.scala 35:20]
  wire [7:0] n7_I_90; // @[Top.scala 35:20]
  wire [7:0] n7_I_91; // @[Top.scala 35:20]
  wire [7:0] n7_I_92; // @[Top.scala 35:20]
  wire [7:0] n7_I_93; // @[Top.scala 35:20]
  wire [7:0] n7_I_94; // @[Top.scala 35:20]
  wire [7:0] n7_I_95; // @[Top.scala 35:20]
  wire [7:0] n7_I_96; // @[Top.scala 35:20]
  wire [7:0] n7_I_97; // @[Top.scala 35:20]
  wire [7:0] n7_I_98; // @[Top.scala 35:20]
  wire [7:0] n7_I_99; // @[Top.scala 35:20]
  wire [7:0] n7_I_100; // @[Top.scala 35:20]
  wire [7:0] n7_I_101; // @[Top.scala 35:20]
  wire [7:0] n7_I_102; // @[Top.scala 35:20]
  wire [7:0] n7_I_103; // @[Top.scala 35:20]
  wire [7:0] n7_I_104; // @[Top.scala 35:20]
  wire [7:0] n7_I_105; // @[Top.scala 35:20]
  wire [7:0] n7_I_106; // @[Top.scala 35:20]
  wire [7:0] n7_I_107; // @[Top.scala 35:20]
  wire [7:0] n7_I_108; // @[Top.scala 35:20]
  wire [7:0] n7_I_109; // @[Top.scala 35:20]
  wire [7:0] n7_I_110; // @[Top.scala 35:20]
  wire [7:0] n7_I_111; // @[Top.scala 35:20]
  wire [7:0] n7_I_112; // @[Top.scala 35:20]
  wire [7:0] n7_I_113; // @[Top.scala 35:20]
  wire [7:0] n7_I_114; // @[Top.scala 35:20]
  wire [7:0] n7_I_115; // @[Top.scala 35:20]
  wire [7:0] n7_I_116; // @[Top.scala 35:20]
  wire [7:0] n7_I_117; // @[Top.scala 35:20]
  wire [7:0] n7_I_118; // @[Top.scala 35:20]
  wire [7:0] n7_I_119; // @[Top.scala 35:20]
  wire [7:0] n7_I_120; // @[Top.scala 35:20]
  wire [7:0] n7_I_121; // @[Top.scala 35:20]
  wire [7:0] n7_I_122; // @[Top.scala 35:20]
  wire [7:0] n7_I_123; // @[Top.scala 35:20]
  wire [7:0] n7_I_124; // @[Top.scala 35:20]
  wire [7:0] n7_I_125; // @[Top.scala 35:20]
  wire [7:0] n7_I_126; // @[Top.scala 35:20]
  wire [7:0] n7_I_127; // @[Top.scala 35:20]
  wire [7:0] n7_I_128; // @[Top.scala 35:20]
  wire [7:0] n7_I_129; // @[Top.scala 35:20]
  wire [7:0] n7_I_130; // @[Top.scala 35:20]
  wire [7:0] n7_I_131; // @[Top.scala 35:20]
  wire [7:0] n7_I_132; // @[Top.scala 35:20]
  wire [7:0] n7_I_133; // @[Top.scala 35:20]
  wire [7:0] n7_I_134; // @[Top.scala 35:20]
  wire [7:0] n7_I_135; // @[Top.scala 35:20]
  wire [7:0] n7_I_136; // @[Top.scala 35:20]
  wire [7:0] n7_I_137; // @[Top.scala 35:20]
  wire [7:0] n7_I_138; // @[Top.scala 35:20]
  wire [7:0] n7_I_139; // @[Top.scala 35:20]
  wire [7:0] n7_I_140; // @[Top.scala 35:20]
  wire [7:0] n7_I_141; // @[Top.scala 35:20]
  wire [7:0] n7_I_142; // @[Top.scala 35:20]
  wire [7:0] n7_I_143; // @[Top.scala 35:20]
  wire [7:0] n7_I_144; // @[Top.scala 35:20]
  wire [7:0] n7_I_145; // @[Top.scala 35:20]
  wire [7:0] n7_I_146; // @[Top.scala 35:20]
  wire [7:0] n7_I_147; // @[Top.scala 35:20]
  wire [7:0] n7_I_148; // @[Top.scala 35:20]
  wire [7:0] n7_I_149; // @[Top.scala 35:20]
  wire [7:0] n7_I_150; // @[Top.scala 35:20]
  wire [7:0] n7_I_151; // @[Top.scala 35:20]
  wire [7:0] n7_I_152; // @[Top.scala 35:20]
  wire [7:0] n7_I_153; // @[Top.scala 35:20]
  wire [7:0] n7_I_154; // @[Top.scala 35:20]
  wire [7:0] n7_I_155; // @[Top.scala 35:20]
  wire [7:0] n7_I_156; // @[Top.scala 35:20]
  wire [7:0] n7_I_157; // @[Top.scala 35:20]
  wire [7:0] n7_I_158; // @[Top.scala 35:20]
  wire [7:0] n7_I_159; // @[Top.scala 35:20]
  wire [7:0] n7_I_160; // @[Top.scala 35:20]
  wire [7:0] n7_I_161; // @[Top.scala 35:20]
  wire [7:0] n7_I_162; // @[Top.scala 35:20]
  wire [7:0] n7_I_163; // @[Top.scala 35:20]
  wire [7:0] n7_I_164; // @[Top.scala 35:20]
  wire [7:0] n7_I_165; // @[Top.scala 35:20]
  wire [7:0] n7_I_166; // @[Top.scala 35:20]
  wire [7:0] n7_I_167; // @[Top.scala 35:20]
  wire [7:0] n7_I_168; // @[Top.scala 35:20]
  wire [7:0] n7_I_169; // @[Top.scala 35:20]
  wire [7:0] n7_I_170; // @[Top.scala 35:20]
  wire [7:0] n7_I_171; // @[Top.scala 35:20]
  wire [7:0] n7_I_172; // @[Top.scala 35:20]
  wire [7:0] n7_I_173; // @[Top.scala 35:20]
  wire [7:0] n7_I_174; // @[Top.scala 35:20]
  wire [7:0] n7_I_175; // @[Top.scala 35:20]
  wire [7:0] n7_I_176; // @[Top.scala 35:20]
  wire [7:0] n7_I_177; // @[Top.scala 35:20]
  wire [7:0] n7_I_178; // @[Top.scala 35:20]
  wire [7:0] n7_I_179; // @[Top.scala 35:20]
  wire [7:0] n7_I_180; // @[Top.scala 35:20]
  wire [7:0] n7_I_181; // @[Top.scala 35:20]
  wire [7:0] n7_I_182; // @[Top.scala 35:20]
  wire [7:0] n7_I_183; // @[Top.scala 35:20]
  wire [7:0] n7_I_184; // @[Top.scala 35:20]
  wire [7:0] n7_I_185; // @[Top.scala 35:20]
  wire [7:0] n7_I_186; // @[Top.scala 35:20]
  wire [7:0] n7_I_187; // @[Top.scala 35:20]
  wire [7:0] n7_I_188; // @[Top.scala 35:20]
  wire [7:0] n7_I_189; // @[Top.scala 35:20]
  wire [7:0] n7_I_190; // @[Top.scala 35:20]
  wire [7:0] n7_I_191; // @[Top.scala 35:20]
  wire [7:0] n7_I_192; // @[Top.scala 35:20]
  wire [7:0] n7_I_193; // @[Top.scala 35:20]
  wire [7:0] n7_I_194; // @[Top.scala 35:20]
  wire [7:0] n7_I_195; // @[Top.scala 35:20]
  wire [7:0] n7_I_196; // @[Top.scala 35:20]
  wire [7:0] n7_I_197; // @[Top.scala 35:20]
  wire [7:0] n7_I_198; // @[Top.scala 35:20]
  wire [7:0] n7_I_199; // @[Top.scala 35:20]
  wire [7:0] n7_O_0; // @[Top.scala 35:20]
  wire [7:0] n7_O_1; // @[Top.scala 35:20]
  wire [7:0] n7_O_2; // @[Top.scala 35:20]
  wire [7:0] n7_O_3; // @[Top.scala 35:20]
  wire [7:0] n7_O_4; // @[Top.scala 35:20]
  wire [7:0] n7_O_5; // @[Top.scala 35:20]
  wire [7:0] n7_O_6; // @[Top.scala 35:20]
  wire [7:0] n7_O_7; // @[Top.scala 35:20]
  wire [7:0] n7_O_8; // @[Top.scala 35:20]
  wire [7:0] n7_O_9; // @[Top.scala 35:20]
  wire [7:0] n7_O_10; // @[Top.scala 35:20]
  wire [7:0] n7_O_11; // @[Top.scala 35:20]
  wire [7:0] n7_O_12; // @[Top.scala 35:20]
  wire [7:0] n7_O_13; // @[Top.scala 35:20]
  wire [7:0] n7_O_14; // @[Top.scala 35:20]
  wire [7:0] n7_O_15; // @[Top.scala 35:20]
  wire [7:0] n7_O_16; // @[Top.scala 35:20]
  wire [7:0] n7_O_17; // @[Top.scala 35:20]
  wire [7:0] n7_O_18; // @[Top.scala 35:20]
  wire [7:0] n7_O_19; // @[Top.scala 35:20]
  wire [7:0] n7_O_20; // @[Top.scala 35:20]
  wire [7:0] n7_O_21; // @[Top.scala 35:20]
  wire [7:0] n7_O_22; // @[Top.scala 35:20]
  wire [7:0] n7_O_23; // @[Top.scala 35:20]
  wire [7:0] n7_O_24; // @[Top.scala 35:20]
  wire [7:0] n7_O_25; // @[Top.scala 35:20]
  wire [7:0] n7_O_26; // @[Top.scala 35:20]
  wire [7:0] n7_O_27; // @[Top.scala 35:20]
  wire [7:0] n7_O_28; // @[Top.scala 35:20]
  wire [7:0] n7_O_29; // @[Top.scala 35:20]
  wire [7:0] n7_O_30; // @[Top.scala 35:20]
  wire [7:0] n7_O_31; // @[Top.scala 35:20]
  wire [7:0] n7_O_32; // @[Top.scala 35:20]
  wire [7:0] n7_O_33; // @[Top.scala 35:20]
  wire [7:0] n7_O_34; // @[Top.scala 35:20]
  wire [7:0] n7_O_35; // @[Top.scala 35:20]
  wire [7:0] n7_O_36; // @[Top.scala 35:20]
  wire [7:0] n7_O_37; // @[Top.scala 35:20]
  wire [7:0] n7_O_38; // @[Top.scala 35:20]
  wire [7:0] n7_O_39; // @[Top.scala 35:20]
  wire [7:0] n7_O_40; // @[Top.scala 35:20]
  wire [7:0] n7_O_41; // @[Top.scala 35:20]
  wire [7:0] n7_O_42; // @[Top.scala 35:20]
  wire [7:0] n7_O_43; // @[Top.scala 35:20]
  wire [7:0] n7_O_44; // @[Top.scala 35:20]
  wire [7:0] n7_O_45; // @[Top.scala 35:20]
  wire [7:0] n7_O_46; // @[Top.scala 35:20]
  wire [7:0] n7_O_47; // @[Top.scala 35:20]
  wire [7:0] n7_O_48; // @[Top.scala 35:20]
  wire [7:0] n7_O_49; // @[Top.scala 35:20]
  wire [7:0] n7_O_50; // @[Top.scala 35:20]
  wire [7:0] n7_O_51; // @[Top.scala 35:20]
  wire [7:0] n7_O_52; // @[Top.scala 35:20]
  wire [7:0] n7_O_53; // @[Top.scala 35:20]
  wire [7:0] n7_O_54; // @[Top.scala 35:20]
  wire [7:0] n7_O_55; // @[Top.scala 35:20]
  wire [7:0] n7_O_56; // @[Top.scala 35:20]
  wire [7:0] n7_O_57; // @[Top.scala 35:20]
  wire [7:0] n7_O_58; // @[Top.scala 35:20]
  wire [7:0] n7_O_59; // @[Top.scala 35:20]
  wire [7:0] n7_O_60; // @[Top.scala 35:20]
  wire [7:0] n7_O_61; // @[Top.scala 35:20]
  wire [7:0] n7_O_62; // @[Top.scala 35:20]
  wire [7:0] n7_O_63; // @[Top.scala 35:20]
  wire [7:0] n7_O_64; // @[Top.scala 35:20]
  wire [7:0] n7_O_65; // @[Top.scala 35:20]
  wire [7:0] n7_O_66; // @[Top.scala 35:20]
  wire [7:0] n7_O_67; // @[Top.scala 35:20]
  wire [7:0] n7_O_68; // @[Top.scala 35:20]
  wire [7:0] n7_O_69; // @[Top.scala 35:20]
  wire [7:0] n7_O_70; // @[Top.scala 35:20]
  wire [7:0] n7_O_71; // @[Top.scala 35:20]
  wire [7:0] n7_O_72; // @[Top.scala 35:20]
  wire [7:0] n7_O_73; // @[Top.scala 35:20]
  wire [7:0] n7_O_74; // @[Top.scala 35:20]
  wire [7:0] n7_O_75; // @[Top.scala 35:20]
  wire [7:0] n7_O_76; // @[Top.scala 35:20]
  wire [7:0] n7_O_77; // @[Top.scala 35:20]
  wire [7:0] n7_O_78; // @[Top.scala 35:20]
  wire [7:0] n7_O_79; // @[Top.scala 35:20]
  wire [7:0] n7_O_80; // @[Top.scala 35:20]
  wire [7:0] n7_O_81; // @[Top.scala 35:20]
  wire [7:0] n7_O_82; // @[Top.scala 35:20]
  wire [7:0] n7_O_83; // @[Top.scala 35:20]
  wire [7:0] n7_O_84; // @[Top.scala 35:20]
  wire [7:0] n7_O_85; // @[Top.scala 35:20]
  wire [7:0] n7_O_86; // @[Top.scala 35:20]
  wire [7:0] n7_O_87; // @[Top.scala 35:20]
  wire [7:0] n7_O_88; // @[Top.scala 35:20]
  wire [7:0] n7_O_89; // @[Top.scala 35:20]
  wire [7:0] n7_O_90; // @[Top.scala 35:20]
  wire [7:0] n7_O_91; // @[Top.scala 35:20]
  wire [7:0] n7_O_92; // @[Top.scala 35:20]
  wire [7:0] n7_O_93; // @[Top.scala 35:20]
  wire [7:0] n7_O_94; // @[Top.scala 35:20]
  wire [7:0] n7_O_95; // @[Top.scala 35:20]
  wire [7:0] n7_O_96; // @[Top.scala 35:20]
  wire [7:0] n7_O_97; // @[Top.scala 35:20]
  wire [7:0] n7_O_98; // @[Top.scala 35:20]
  wire [7:0] n7_O_99; // @[Top.scala 35:20]
  wire [7:0] n7_O_100; // @[Top.scala 35:20]
  wire [7:0] n7_O_101; // @[Top.scala 35:20]
  wire [7:0] n7_O_102; // @[Top.scala 35:20]
  wire [7:0] n7_O_103; // @[Top.scala 35:20]
  wire [7:0] n7_O_104; // @[Top.scala 35:20]
  wire [7:0] n7_O_105; // @[Top.scala 35:20]
  wire [7:0] n7_O_106; // @[Top.scala 35:20]
  wire [7:0] n7_O_107; // @[Top.scala 35:20]
  wire [7:0] n7_O_108; // @[Top.scala 35:20]
  wire [7:0] n7_O_109; // @[Top.scala 35:20]
  wire [7:0] n7_O_110; // @[Top.scala 35:20]
  wire [7:0] n7_O_111; // @[Top.scala 35:20]
  wire [7:0] n7_O_112; // @[Top.scala 35:20]
  wire [7:0] n7_O_113; // @[Top.scala 35:20]
  wire [7:0] n7_O_114; // @[Top.scala 35:20]
  wire [7:0] n7_O_115; // @[Top.scala 35:20]
  wire [7:0] n7_O_116; // @[Top.scala 35:20]
  wire [7:0] n7_O_117; // @[Top.scala 35:20]
  wire [7:0] n7_O_118; // @[Top.scala 35:20]
  wire [7:0] n7_O_119; // @[Top.scala 35:20]
  wire [7:0] n7_O_120; // @[Top.scala 35:20]
  wire [7:0] n7_O_121; // @[Top.scala 35:20]
  wire [7:0] n7_O_122; // @[Top.scala 35:20]
  wire [7:0] n7_O_123; // @[Top.scala 35:20]
  wire [7:0] n7_O_124; // @[Top.scala 35:20]
  wire [7:0] n7_O_125; // @[Top.scala 35:20]
  wire [7:0] n7_O_126; // @[Top.scala 35:20]
  wire [7:0] n7_O_127; // @[Top.scala 35:20]
  wire [7:0] n7_O_128; // @[Top.scala 35:20]
  wire [7:0] n7_O_129; // @[Top.scala 35:20]
  wire [7:0] n7_O_130; // @[Top.scala 35:20]
  wire [7:0] n7_O_131; // @[Top.scala 35:20]
  wire [7:0] n7_O_132; // @[Top.scala 35:20]
  wire [7:0] n7_O_133; // @[Top.scala 35:20]
  wire [7:0] n7_O_134; // @[Top.scala 35:20]
  wire [7:0] n7_O_135; // @[Top.scala 35:20]
  wire [7:0] n7_O_136; // @[Top.scala 35:20]
  wire [7:0] n7_O_137; // @[Top.scala 35:20]
  wire [7:0] n7_O_138; // @[Top.scala 35:20]
  wire [7:0] n7_O_139; // @[Top.scala 35:20]
  wire [7:0] n7_O_140; // @[Top.scala 35:20]
  wire [7:0] n7_O_141; // @[Top.scala 35:20]
  wire [7:0] n7_O_142; // @[Top.scala 35:20]
  wire [7:0] n7_O_143; // @[Top.scala 35:20]
  wire [7:0] n7_O_144; // @[Top.scala 35:20]
  wire [7:0] n7_O_145; // @[Top.scala 35:20]
  wire [7:0] n7_O_146; // @[Top.scala 35:20]
  wire [7:0] n7_O_147; // @[Top.scala 35:20]
  wire [7:0] n7_O_148; // @[Top.scala 35:20]
  wire [7:0] n7_O_149; // @[Top.scala 35:20]
  wire [7:0] n7_O_150; // @[Top.scala 35:20]
  wire [7:0] n7_O_151; // @[Top.scala 35:20]
  wire [7:0] n7_O_152; // @[Top.scala 35:20]
  wire [7:0] n7_O_153; // @[Top.scala 35:20]
  wire [7:0] n7_O_154; // @[Top.scala 35:20]
  wire [7:0] n7_O_155; // @[Top.scala 35:20]
  wire [7:0] n7_O_156; // @[Top.scala 35:20]
  wire [7:0] n7_O_157; // @[Top.scala 35:20]
  wire [7:0] n7_O_158; // @[Top.scala 35:20]
  wire [7:0] n7_O_159; // @[Top.scala 35:20]
  wire [7:0] n7_O_160; // @[Top.scala 35:20]
  wire [7:0] n7_O_161; // @[Top.scala 35:20]
  wire [7:0] n7_O_162; // @[Top.scala 35:20]
  wire [7:0] n7_O_163; // @[Top.scala 35:20]
  wire [7:0] n7_O_164; // @[Top.scala 35:20]
  wire [7:0] n7_O_165; // @[Top.scala 35:20]
  wire [7:0] n7_O_166; // @[Top.scala 35:20]
  wire [7:0] n7_O_167; // @[Top.scala 35:20]
  wire [7:0] n7_O_168; // @[Top.scala 35:20]
  wire [7:0] n7_O_169; // @[Top.scala 35:20]
  wire [7:0] n7_O_170; // @[Top.scala 35:20]
  wire [7:0] n7_O_171; // @[Top.scala 35:20]
  wire [7:0] n7_O_172; // @[Top.scala 35:20]
  wire [7:0] n7_O_173; // @[Top.scala 35:20]
  wire [7:0] n7_O_174; // @[Top.scala 35:20]
  wire [7:0] n7_O_175; // @[Top.scala 35:20]
  wire [7:0] n7_O_176; // @[Top.scala 35:20]
  wire [7:0] n7_O_177; // @[Top.scala 35:20]
  wire [7:0] n7_O_178; // @[Top.scala 35:20]
  wire [7:0] n7_O_179; // @[Top.scala 35:20]
  wire [7:0] n7_O_180; // @[Top.scala 35:20]
  wire [7:0] n7_O_181; // @[Top.scala 35:20]
  wire [7:0] n7_O_182; // @[Top.scala 35:20]
  wire [7:0] n7_O_183; // @[Top.scala 35:20]
  wire [7:0] n7_O_184; // @[Top.scala 35:20]
  wire [7:0] n7_O_185; // @[Top.scala 35:20]
  wire [7:0] n7_O_186; // @[Top.scala 35:20]
  wire [7:0] n7_O_187; // @[Top.scala 35:20]
  wire [7:0] n7_O_188; // @[Top.scala 35:20]
  wire [7:0] n7_O_189; // @[Top.scala 35:20]
  wire [7:0] n7_O_190; // @[Top.scala 35:20]
  wire [7:0] n7_O_191; // @[Top.scala 35:20]
  wire [7:0] n7_O_192; // @[Top.scala 35:20]
  wire [7:0] n7_O_193; // @[Top.scala 35:20]
  wire [7:0] n7_O_194; // @[Top.scala 35:20]
  wire [7:0] n7_O_195; // @[Top.scala 35:20]
  wire [7:0] n7_O_196; // @[Top.scala 35:20]
  wire [7:0] n7_O_197; // @[Top.scala 35:20]
  wire [7:0] n7_O_198; // @[Top.scala 35:20]
  wire [7:0] n7_O_199; // @[Top.scala 35:20]
  wire  n8_clock; // @[Top.scala 38:20]
  wire  n8_reset; // @[Top.scala 38:20]
  wire  n8_valid_up; // @[Top.scala 38:20]
  wire  n8_valid_down; // @[Top.scala 38:20]
  wire [7:0] n8_I_0; // @[Top.scala 38:20]
  wire [7:0] n8_I_1; // @[Top.scala 38:20]
  wire [7:0] n8_I_2; // @[Top.scala 38:20]
  wire [7:0] n8_I_3; // @[Top.scala 38:20]
  wire [7:0] n8_I_4; // @[Top.scala 38:20]
  wire [7:0] n8_I_5; // @[Top.scala 38:20]
  wire [7:0] n8_I_6; // @[Top.scala 38:20]
  wire [7:0] n8_I_7; // @[Top.scala 38:20]
  wire [7:0] n8_I_8; // @[Top.scala 38:20]
  wire [7:0] n8_I_9; // @[Top.scala 38:20]
  wire [7:0] n8_I_10; // @[Top.scala 38:20]
  wire [7:0] n8_I_11; // @[Top.scala 38:20]
  wire [7:0] n8_I_12; // @[Top.scala 38:20]
  wire [7:0] n8_I_13; // @[Top.scala 38:20]
  wire [7:0] n8_I_14; // @[Top.scala 38:20]
  wire [7:0] n8_I_15; // @[Top.scala 38:20]
  wire [7:0] n8_I_16; // @[Top.scala 38:20]
  wire [7:0] n8_I_17; // @[Top.scala 38:20]
  wire [7:0] n8_I_18; // @[Top.scala 38:20]
  wire [7:0] n8_I_19; // @[Top.scala 38:20]
  wire [7:0] n8_I_20; // @[Top.scala 38:20]
  wire [7:0] n8_I_21; // @[Top.scala 38:20]
  wire [7:0] n8_I_22; // @[Top.scala 38:20]
  wire [7:0] n8_I_23; // @[Top.scala 38:20]
  wire [7:0] n8_I_24; // @[Top.scala 38:20]
  wire [7:0] n8_I_25; // @[Top.scala 38:20]
  wire [7:0] n8_I_26; // @[Top.scala 38:20]
  wire [7:0] n8_I_27; // @[Top.scala 38:20]
  wire [7:0] n8_I_28; // @[Top.scala 38:20]
  wire [7:0] n8_I_29; // @[Top.scala 38:20]
  wire [7:0] n8_I_30; // @[Top.scala 38:20]
  wire [7:0] n8_I_31; // @[Top.scala 38:20]
  wire [7:0] n8_I_32; // @[Top.scala 38:20]
  wire [7:0] n8_I_33; // @[Top.scala 38:20]
  wire [7:0] n8_I_34; // @[Top.scala 38:20]
  wire [7:0] n8_I_35; // @[Top.scala 38:20]
  wire [7:0] n8_I_36; // @[Top.scala 38:20]
  wire [7:0] n8_I_37; // @[Top.scala 38:20]
  wire [7:0] n8_I_38; // @[Top.scala 38:20]
  wire [7:0] n8_I_39; // @[Top.scala 38:20]
  wire [7:0] n8_I_40; // @[Top.scala 38:20]
  wire [7:0] n8_I_41; // @[Top.scala 38:20]
  wire [7:0] n8_I_42; // @[Top.scala 38:20]
  wire [7:0] n8_I_43; // @[Top.scala 38:20]
  wire [7:0] n8_I_44; // @[Top.scala 38:20]
  wire [7:0] n8_I_45; // @[Top.scala 38:20]
  wire [7:0] n8_I_46; // @[Top.scala 38:20]
  wire [7:0] n8_I_47; // @[Top.scala 38:20]
  wire [7:0] n8_I_48; // @[Top.scala 38:20]
  wire [7:0] n8_I_49; // @[Top.scala 38:20]
  wire [7:0] n8_I_50; // @[Top.scala 38:20]
  wire [7:0] n8_I_51; // @[Top.scala 38:20]
  wire [7:0] n8_I_52; // @[Top.scala 38:20]
  wire [7:0] n8_I_53; // @[Top.scala 38:20]
  wire [7:0] n8_I_54; // @[Top.scala 38:20]
  wire [7:0] n8_I_55; // @[Top.scala 38:20]
  wire [7:0] n8_I_56; // @[Top.scala 38:20]
  wire [7:0] n8_I_57; // @[Top.scala 38:20]
  wire [7:0] n8_I_58; // @[Top.scala 38:20]
  wire [7:0] n8_I_59; // @[Top.scala 38:20]
  wire [7:0] n8_I_60; // @[Top.scala 38:20]
  wire [7:0] n8_I_61; // @[Top.scala 38:20]
  wire [7:0] n8_I_62; // @[Top.scala 38:20]
  wire [7:0] n8_I_63; // @[Top.scala 38:20]
  wire [7:0] n8_I_64; // @[Top.scala 38:20]
  wire [7:0] n8_I_65; // @[Top.scala 38:20]
  wire [7:0] n8_I_66; // @[Top.scala 38:20]
  wire [7:0] n8_I_67; // @[Top.scala 38:20]
  wire [7:0] n8_I_68; // @[Top.scala 38:20]
  wire [7:0] n8_I_69; // @[Top.scala 38:20]
  wire [7:0] n8_I_70; // @[Top.scala 38:20]
  wire [7:0] n8_I_71; // @[Top.scala 38:20]
  wire [7:0] n8_I_72; // @[Top.scala 38:20]
  wire [7:0] n8_I_73; // @[Top.scala 38:20]
  wire [7:0] n8_I_74; // @[Top.scala 38:20]
  wire [7:0] n8_I_75; // @[Top.scala 38:20]
  wire [7:0] n8_I_76; // @[Top.scala 38:20]
  wire [7:0] n8_I_77; // @[Top.scala 38:20]
  wire [7:0] n8_I_78; // @[Top.scala 38:20]
  wire [7:0] n8_I_79; // @[Top.scala 38:20]
  wire [7:0] n8_I_80; // @[Top.scala 38:20]
  wire [7:0] n8_I_81; // @[Top.scala 38:20]
  wire [7:0] n8_I_82; // @[Top.scala 38:20]
  wire [7:0] n8_I_83; // @[Top.scala 38:20]
  wire [7:0] n8_I_84; // @[Top.scala 38:20]
  wire [7:0] n8_I_85; // @[Top.scala 38:20]
  wire [7:0] n8_I_86; // @[Top.scala 38:20]
  wire [7:0] n8_I_87; // @[Top.scala 38:20]
  wire [7:0] n8_I_88; // @[Top.scala 38:20]
  wire [7:0] n8_I_89; // @[Top.scala 38:20]
  wire [7:0] n8_I_90; // @[Top.scala 38:20]
  wire [7:0] n8_I_91; // @[Top.scala 38:20]
  wire [7:0] n8_I_92; // @[Top.scala 38:20]
  wire [7:0] n8_I_93; // @[Top.scala 38:20]
  wire [7:0] n8_I_94; // @[Top.scala 38:20]
  wire [7:0] n8_I_95; // @[Top.scala 38:20]
  wire [7:0] n8_I_96; // @[Top.scala 38:20]
  wire [7:0] n8_I_97; // @[Top.scala 38:20]
  wire [7:0] n8_I_98; // @[Top.scala 38:20]
  wire [7:0] n8_I_99; // @[Top.scala 38:20]
  wire [7:0] n8_I_100; // @[Top.scala 38:20]
  wire [7:0] n8_I_101; // @[Top.scala 38:20]
  wire [7:0] n8_I_102; // @[Top.scala 38:20]
  wire [7:0] n8_I_103; // @[Top.scala 38:20]
  wire [7:0] n8_I_104; // @[Top.scala 38:20]
  wire [7:0] n8_I_105; // @[Top.scala 38:20]
  wire [7:0] n8_I_106; // @[Top.scala 38:20]
  wire [7:0] n8_I_107; // @[Top.scala 38:20]
  wire [7:0] n8_I_108; // @[Top.scala 38:20]
  wire [7:0] n8_I_109; // @[Top.scala 38:20]
  wire [7:0] n8_I_110; // @[Top.scala 38:20]
  wire [7:0] n8_I_111; // @[Top.scala 38:20]
  wire [7:0] n8_I_112; // @[Top.scala 38:20]
  wire [7:0] n8_I_113; // @[Top.scala 38:20]
  wire [7:0] n8_I_114; // @[Top.scala 38:20]
  wire [7:0] n8_I_115; // @[Top.scala 38:20]
  wire [7:0] n8_I_116; // @[Top.scala 38:20]
  wire [7:0] n8_I_117; // @[Top.scala 38:20]
  wire [7:0] n8_I_118; // @[Top.scala 38:20]
  wire [7:0] n8_I_119; // @[Top.scala 38:20]
  wire [7:0] n8_I_120; // @[Top.scala 38:20]
  wire [7:0] n8_I_121; // @[Top.scala 38:20]
  wire [7:0] n8_I_122; // @[Top.scala 38:20]
  wire [7:0] n8_I_123; // @[Top.scala 38:20]
  wire [7:0] n8_I_124; // @[Top.scala 38:20]
  wire [7:0] n8_I_125; // @[Top.scala 38:20]
  wire [7:0] n8_I_126; // @[Top.scala 38:20]
  wire [7:0] n8_I_127; // @[Top.scala 38:20]
  wire [7:0] n8_I_128; // @[Top.scala 38:20]
  wire [7:0] n8_I_129; // @[Top.scala 38:20]
  wire [7:0] n8_I_130; // @[Top.scala 38:20]
  wire [7:0] n8_I_131; // @[Top.scala 38:20]
  wire [7:0] n8_I_132; // @[Top.scala 38:20]
  wire [7:0] n8_I_133; // @[Top.scala 38:20]
  wire [7:0] n8_I_134; // @[Top.scala 38:20]
  wire [7:0] n8_I_135; // @[Top.scala 38:20]
  wire [7:0] n8_I_136; // @[Top.scala 38:20]
  wire [7:0] n8_I_137; // @[Top.scala 38:20]
  wire [7:0] n8_I_138; // @[Top.scala 38:20]
  wire [7:0] n8_I_139; // @[Top.scala 38:20]
  wire [7:0] n8_I_140; // @[Top.scala 38:20]
  wire [7:0] n8_I_141; // @[Top.scala 38:20]
  wire [7:0] n8_I_142; // @[Top.scala 38:20]
  wire [7:0] n8_I_143; // @[Top.scala 38:20]
  wire [7:0] n8_I_144; // @[Top.scala 38:20]
  wire [7:0] n8_I_145; // @[Top.scala 38:20]
  wire [7:0] n8_I_146; // @[Top.scala 38:20]
  wire [7:0] n8_I_147; // @[Top.scala 38:20]
  wire [7:0] n8_I_148; // @[Top.scala 38:20]
  wire [7:0] n8_I_149; // @[Top.scala 38:20]
  wire [7:0] n8_I_150; // @[Top.scala 38:20]
  wire [7:0] n8_I_151; // @[Top.scala 38:20]
  wire [7:0] n8_I_152; // @[Top.scala 38:20]
  wire [7:0] n8_I_153; // @[Top.scala 38:20]
  wire [7:0] n8_I_154; // @[Top.scala 38:20]
  wire [7:0] n8_I_155; // @[Top.scala 38:20]
  wire [7:0] n8_I_156; // @[Top.scala 38:20]
  wire [7:0] n8_I_157; // @[Top.scala 38:20]
  wire [7:0] n8_I_158; // @[Top.scala 38:20]
  wire [7:0] n8_I_159; // @[Top.scala 38:20]
  wire [7:0] n8_I_160; // @[Top.scala 38:20]
  wire [7:0] n8_I_161; // @[Top.scala 38:20]
  wire [7:0] n8_I_162; // @[Top.scala 38:20]
  wire [7:0] n8_I_163; // @[Top.scala 38:20]
  wire [7:0] n8_I_164; // @[Top.scala 38:20]
  wire [7:0] n8_I_165; // @[Top.scala 38:20]
  wire [7:0] n8_I_166; // @[Top.scala 38:20]
  wire [7:0] n8_I_167; // @[Top.scala 38:20]
  wire [7:0] n8_I_168; // @[Top.scala 38:20]
  wire [7:0] n8_I_169; // @[Top.scala 38:20]
  wire [7:0] n8_I_170; // @[Top.scala 38:20]
  wire [7:0] n8_I_171; // @[Top.scala 38:20]
  wire [7:0] n8_I_172; // @[Top.scala 38:20]
  wire [7:0] n8_I_173; // @[Top.scala 38:20]
  wire [7:0] n8_I_174; // @[Top.scala 38:20]
  wire [7:0] n8_I_175; // @[Top.scala 38:20]
  wire [7:0] n8_I_176; // @[Top.scala 38:20]
  wire [7:0] n8_I_177; // @[Top.scala 38:20]
  wire [7:0] n8_I_178; // @[Top.scala 38:20]
  wire [7:0] n8_I_179; // @[Top.scala 38:20]
  wire [7:0] n8_I_180; // @[Top.scala 38:20]
  wire [7:0] n8_I_181; // @[Top.scala 38:20]
  wire [7:0] n8_I_182; // @[Top.scala 38:20]
  wire [7:0] n8_I_183; // @[Top.scala 38:20]
  wire [7:0] n8_I_184; // @[Top.scala 38:20]
  wire [7:0] n8_I_185; // @[Top.scala 38:20]
  wire [7:0] n8_I_186; // @[Top.scala 38:20]
  wire [7:0] n8_I_187; // @[Top.scala 38:20]
  wire [7:0] n8_I_188; // @[Top.scala 38:20]
  wire [7:0] n8_I_189; // @[Top.scala 38:20]
  wire [7:0] n8_I_190; // @[Top.scala 38:20]
  wire [7:0] n8_I_191; // @[Top.scala 38:20]
  wire [7:0] n8_I_192; // @[Top.scala 38:20]
  wire [7:0] n8_I_193; // @[Top.scala 38:20]
  wire [7:0] n8_I_194; // @[Top.scala 38:20]
  wire [7:0] n8_I_195; // @[Top.scala 38:20]
  wire [7:0] n8_I_196; // @[Top.scala 38:20]
  wire [7:0] n8_I_197; // @[Top.scala 38:20]
  wire [7:0] n8_I_198; // @[Top.scala 38:20]
  wire [7:0] n8_I_199; // @[Top.scala 38:20]
  wire [7:0] n8_O_0; // @[Top.scala 38:20]
  wire [7:0] n8_O_1; // @[Top.scala 38:20]
  wire [7:0] n8_O_2; // @[Top.scala 38:20]
  wire [7:0] n8_O_3; // @[Top.scala 38:20]
  wire [7:0] n8_O_4; // @[Top.scala 38:20]
  wire [7:0] n8_O_5; // @[Top.scala 38:20]
  wire [7:0] n8_O_6; // @[Top.scala 38:20]
  wire [7:0] n8_O_7; // @[Top.scala 38:20]
  wire [7:0] n8_O_8; // @[Top.scala 38:20]
  wire [7:0] n8_O_9; // @[Top.scala 38:20]
  wire [7:0] n8_O_10; // @[Top.scala 38:20]
  wire [7:0] n8_O_11; // @[Top.scala 38:20]
  wire [7:0] n8_O_12; // @[Top.scala 38:20]
  wire [7:0] n8_O_13; // @[Top.scala 38:20]
  wire [7:0] n8_O_14; // @[Top.scala 38:20]
  wire [7:0] n8_O_15; // @[Top.scala 38:20]
  wire [7:0] n8_O_16; // @[Top.scala 38:20]
  wire [7:0] n8_O_17; // @[Top.scala 38:20]
  wire [7:0] n8_O_18; // @[Top.scala 38:20]
  wire [7:0] n8_O_19; // @[Top.scala 38:20]
  wire [7:0] n8_O_20; // @[Top.scala 38:20]
  wire [7:0] n8_O_21; // @[Top.scala 38:20]
  wire [7:0] n8_O_22; // @[Top.scala 38:20]
  wire [7:0] n8_O_23; // @[Top.scala 38:20]
  wire [7:0] n8_O_24; // @[Top.scala 38:20]
  wire [7:0] n8_O_25; // @[Top.scala 38:20]
  wire [7:0] n8_O_26; // @[Top.scala 38:20]
  wire [7:0] n8_O_27; // @[Top.scala 38:20]
  wire [7:0] n8_O_28; // @[Top.scala 38:20]
  wire [7:0] n8_O_29; // @[Top.scala 38:20]
  wire [7:0] n8_O_30; // @[Top.scala 38:20]
  wire [7:0] n8_O_31; // @[Top.scala 38:20]
  wire [7:0] n8_O_32; // @[Top.scala 38:20]
  wire [7:0] n8_O_33; // @[Top.scala 38:20]
  wire [7:0] n8_O_34; // @[Top.scala 38:20]
  wire [7:0] n8_O_35; // @[Top.scala 38:20]
  wire [7:0] n8_O_36; // @[Top.scala 38:20]
  wire [7:0] n8_O_37; // @[Top.scala 38:20]
  wire [7:0] n8_O_38; // @[Top.scala 38:20]
  wire [7:0] n8_O_39; // @[Top.scala 38:20]
  wire [7:0] n8_O_40; // @[Top.scala 38:20]
  wire [7:0] n8_O_41; // @[Top.scala 38:20]
  wire [7:0] n8_O_42; // @[Top.scala 38:20]
  wire [7:0] n8_O_43; // @[Top.scala 38:20]
  wire [7:0] n8_O_44; // @[Top.scala 38:20]
  wire [7:0] n8_O_45; // @[Top.scala 38:20]
  wire [7:0] n8_O_46; // @[Top.scala 38:20]
  wire [7:0] n8_O_47; // @[Top.scala 38:20]
  wire [7:0] n8_O_48; // @[Top.scala 38:20]
  wire [7:0] n8_O_49; // @[Top.scala 38:20]
  wire [7:0] n8_O_50; // @[Top.scala 38:20]
  wire [7:0] n8_O_51; // @[Top.scala 38:20]
  wire [7:0] n8_O_52; // @[Top.scala 38:20]
  wire [7:0] n8_O_53; // @[Top.scala 38:20]
  wire [7:0] n8_O_54; // @[Top.scala 38:20]
  wire [7:0] n8_O_55; // @[Top.scala 38:20]
  wire [7:0] n8_O_56; // @[Top.scala 38:20]
  wire [7:0] n8_O_57; // @[Top.scala 38:20]
  wire [7:0] n8_O_58; // @[Top.scala 38:20]
  wire [7:0] n8_O_59; // @[Top.scala 38:20]
  wire [7:0] n8_O_60; // @[Top.scala 38:20]
  wire [7:0] n8_O_61; // @[Top.scala 38:20]
  wire [7:0] n8_O_62; // @[Top.scala 38:20]
  wire [7:0] n8_O_63; // @[Top.scala 38:20]
  wire [7:0] n8_O_64; // @[Top.scala 38:20]
  wire [7:0] n8_O_65; // @[Top.scala 38:20]
  wire [7:0] n8_O_66; // @[Top.scala 38:20]
  wire [7:0] n8_O_67; // @[Top.scala 38:20]
  wire [7:0] n8_O_68; // @[Top.scala 38:20]
  wire [7:0] n8_O_69; // @[Top.scala 38:20]
  wire [7:0] n8_O_70; // @[Top.scala 38:20]
  wire [7:0] n8_O_71; // @[Top.scala 38:20]
  wire [7:0] n8_O_72; // @[Top.scala 38:20]
  wire [7:0] n8_O_73; // @[Top.scala 38:20]
  wire [7:0] n8_O_74; // @[Top.scala 38:20]
  wire [7:0] n8_O_75; // @[Top.scala 38:20]
  wire [7:0] n8_O_76; // @[Top.scala 38:20]
  wire [7:0] n8_O_77; // @[Top.scala 38:20]
  wire [7:0] n8_O_78; // @[Top.scala 38:20]
  wire [7:0] n8_O_79; // @[Top.scala 38:20]
  wire [7:0] n8_O_80; // @[Top.scala 38:20]
  wire [7:0] n8_O_81; // @[Top.scala 38:20]
  wire [7:0] n8_O_82; // @[Top.scala 38:20]
  wire [7:0] n8_O_83; // @[Top.scala 38:20]
  wire [7:0] n8_O_84; // @[Top.scala 38:20]
  wire [7:0] n8_O_85; // @[Top.scala 38:20]
  wire [7:0] n8_O_86; // @[Top.scala 38:20]
  wire [7:0] n8_O_87; // @[Top.scala 38:20]
  wire [7:0] n8_O_88; // @[Top.scala 38:20]
  wire [7:0] n8_O_89; // @[Top.scala 38:20]
  wire [7:0] n8_O_90; // @[Top.scala 38:20]
  wire [7:0] n8_O_91; // @[Top.scala 38:20]
  wire [7:0] n8_O_92; // @[Top.scala 38:20]
  wire [7:0] n8_O_93; // @[Top.scala 38:20]
  wire [7:0] n8_O_94; // @[Top.scala 38:20]
  wire [7:0] n8_O_95; // @[Top.scala 38:20]
  wire [7:0] n8_O_96; // @[Top.scala 38:20]
  wire [7:0] n8_O_97; // @[Top.scala 38:20]
  wire [7:0] n8_O_98; // @[Top.scala 38:20]
  wire [7:0] n8_O_99; // @[Top.scala 38:20]
  wire [7:0] n8_O_100; // @[Top.scala 38:20]
  wire [7:0] n8_O_101; // @[Top.scala 38:20]
  wire [7:0] n8_O_102; // @[Top.scala 38:20]
  wire [7:0] n8_O_103; // @[Top.scala 38:20]
  wire [7:0] n8_O_104; // @[Top.scala 38:20]
  wire [7:0] n8_O_105; // @[Top.scala 38:20]
  wire [7:0] n8_O_106; // @[Top.scala 38:20]
  wire [7:0] n8_O_107; // @[Top.scala 38:20]
  wire [7:0] n8_O_108; // @[Top.scala 38:20]
  wire [7:0] n8_O_109; // @[Top.scala 38:20]
  wire [7:0] n8_O_110; // @[Top.scala 38:20]
  wire [7:0] n8_O_111; // @[Top.scala 38:20]
  wire [7:0] n8_O_112; // @[Top.scala 38:20]
  wire [7:0] n8_O_113; // @[Top.scala 38:20]
  wire [7:0] n8_O_114; // @[Top.scala 38:20]
  wire [7:0] n8_O_115; // @[Top.scala 38:20]
  wire [7:0] n8_O_116; // @[Top.scala 38:20]
  wire [7:0] n8_O_117; // @[Top.scala 38:20]
  wire [7:0] n8_O_118; // @[Top.scala 38:20]
  wire [7:0] n8_O_119; // @[Top.scala 38:20]
  wire [7:0] n8_O_120; // @[Top.scala 38:20]
  wire [7:0] n8_O_121; // @[Top.scala 38:20]
  wire [7:0] n8_O_122; // @[Top.scala 38:20]
  wire [7:0] n8_O_123; // @[Top.scala 38:20]
  wire [7:0] n8_O_124; // @[Top.scala 38:20]
  wire [7:0] n8_O_125; // @[Top.scala 38:20]
  wire [7:0] n8_O_126; // @[Top.scala 38:20]
  wire [7:0] n8_O_127; // @[Top.scala 38:20]
  wire [7:0] n8_O_128; // @[Top.scala 38:20]
  wire [7:0] n8_O_129; // @[Top.scala 38:20]
  wire [7:0] n8_O_130; // @[Top.scala 38:20]
  wire [7:0] n8_O_131; // @[Top.scala 38:20]
  wire [7:0] n8_O_132; // @[Top.scala 38:20]
  wire [7:0] n8_O_133; // @[Top.scala 38:20]
  wire [7:0] n8_O_134; // @[Top.scala 38:20]
  wire [7:0] n8_O_135; // @[Top.scala 38:20]
  wire [7:0] n8_O_136; // @[Top.scala 38:20]
  wire [7:0] n8_O_137; // @[Top.scala 38:20]
  wire [7:0] n8_O_138; // @[Top.scala 38:20]
  wire [7:0] n8_O_139; // @[Top.scala 38:20]
  wire [7:0] n8_O_140; // @[Top.scala 38:20]
  wire [7:0] n8_O_141; // @[Top.scala 38:20]
  wire [7:0] n8_O_142; // @[Top.scala 38:20]
  wire [7:0] n8_O_143; // @[Top.scala 38:20]
  wire [7:0] n8_O_144; // @[Top.scala 38:20]
  wire [7:0] n8_O_145; // @[Top.scala 38:20]
  wire [7:0] n8_O_146; // @[Top.scala 38:20]
  wire [7:0] n8_O_147; // @[Top.scala 38:20]
  wire [7:0] n8_O_148; // @[Top.scala 38:20]
  wire [7:0] n8_O_149; // @[Top.scala 38:20]
  wire [7:0] n8_O_150; // @[Top.scala 38:20]
  wire [7:0] n8_O_151; // @[Top.scala 38:20]
  wire [7:0] n8_O_152; // @[Top.scala 38:20]
  wire [7:0] n8_O_153; // @[Top.scala 38:20]
  wire [7:0] n8_O_154; // @[Top.scala 38:20]
  wire [7:0] n8_O_155; // @[Top.scala 38:20]
  wire [7:0] n8_O_156; // @[Top.scala 38:20]
  wire [7:0] n8_O_157; // @[Top.scala 38:20]
  wire [7:0] n8_O_158; // @[Top.scala 38:20]
  wire [7:0] n8_O_159; // @[Top.scala 38:20]
  wire [7:0] n8_O_160; // @[Top.scala 38:20]
  wire [7:0] n8_O_161; // @[Top.scala 38:20]
  wire [7:0] n8_O_162; // @[Top.scala 38:20]
  wire [7:0] n8_O_163; // @[Top.scala 38:20]
  wire [7:0] n8_O_164; // @[Top.scala 38:20]
  wire [7:0] n8_O_165; // @[Top.scala 38:20]
  wire [7:0] n8_O_166; // @[Top.scala 38:20]
  wire [7:0] n8_O_167; // @[Top.scala 38:20]
  wire [7:0] n8_O_168; // @[Top.scala 38:20]
  wire [7:0] n8_O_169; // @[Top.scala 38:20]
  wire [7:0] n8_O_170; // @[Top.scala 38:20]
  wire [7:0] n8_O_171; // @[Top.scala 38:20]
  wire [7:0] n8_O_172; // @[Top.scala 38:20]
  wire [7:0] n8_O_173; // @[Top.scala 38:20]
  wire [7:0] n8_O_174; // @[Top.scala 38:20]
  wire [7:0] n8_O_175; // @[Top.scala 38:20]
  wire [7:0] n8_O_176; // @[Top.scala 38:20]
  wire [7:0] n8_O_177; // @[Top.scala 38:20]
  wire [7:0] n8_O_178; // @[Top.scala 38:20]
  wire [7:0] n8_O_179; // @[Top.scala 38:20]
  wire [7:0] n8_O_180; // @[Top.scala 38:20]
  wire [7:0] n8_O_181; // @[Top.scala 38:20]
  wire [7:0] n8_O_182; // @[Top.scala 38:20]
  wire [7:0] n8_O_183; // @[Top.scala 38:20]
  wire [7:0] n8_O_184; // @[Top.scala 38:20]
  wire [7:0] n8_O_185; // @[Top.scala 38:20]
  wire [7:0] n8_O_186; // @[Top.scala 38:20]
  wire [7:0] n8_O_187; // @[Top.scala 38:20]
  wire [7:0] n8_O_188; // @[Top.scala 38:20]
  wire [7:0] n8_O_189; // @[Top.scala 38:20]
  wire [7:0] n8_O_190; // @[Top.scala 38:20]
  wire [7:0] n8_O_191; // @[Top.scala 38:20]
  wire [7:0] n8_O_192; // @[Top.scala 38:20]
  wire [7:0] n8_O_193; // @[Top.scala 38:20]
  wire [7:0] n8_O_194; // @[Top.scala 38:20]
  wire [7:0] n8_O_195; // @[Top.scala 38:20]
  wire [7:0] n8_O_196; // @[Top.scala 38:20]
  wire [7:0] n8_O_197; // @[Top.scala 38:20]
  wire [7:0] n8_O_198; // @[Top.scala 38:20]
  wire [7:0] n8_O_199; // @[Top.scala 38:20]
  wire  n9_clock; // @[Top.scala 41:20]
  wire  n9_reset; // @[Top.scala 41:20]
  wire  n9_valid_up; // @[Top.scala 41:20]
  wire  n9_valid_down; // @[Top.scala 41:20]
  wire [7:0] n9_I_0; // @[Top.scala 41:20]
  wire [7:0] n9_I_1; // @[Top.scala 41:20]
  wire [7:0] n9_I_2; // @[Top.scala 41:20]
  wire [7:0] n9_I_3; // @[Top.scala 41:20]
  wire [7:0] n9_I_4; // @[Top.scala 41:20]
  wire [7:0] n9_I_5; // @[Top.scala 41:20]
  wire [7:0] n9_I_6; // @[Top.scala 41:20]
  wire [7:0] n9_I_7; // @[Top.scala 41:20]
  wire [7:0] n9_I_8; // @[Top.scala 41:20]
  wire [7:0] n9_I_9; // @[Top.scala 41:20]
  wire [7:0] n9_I_10; // @[Top.scala 41:20]
  wire [7:0] n9_I_11; // @[Top.scala 41:20]
  wire [7:0] n9_I_12; // @[Top.scala 41:20]
  wire [7:0] n9_I_13; // @[Top.scala 41:20]
  wire [7:0] n9_I_14; // @[Top.scala 41:20]
  wire [7:0] n9_I_15; // @[Top.scala 41:20]
  wire [7:0] n9_I_16; // @[Top.scala 41:20]
  wire [7:0] n9_I_17; // @[Top.scala 41:20]
  wire [7:0] n9_I_18; // @[Top.scala 41:20]
  wire [7:0] n9_I_19; // @[Top.scala 41:20]
  wire [7:0] n9_I_20; // @[Top.scala 41:20]
  wire [7:0] n9_I_21; // @[Top.scala 41:20]
  wire [7:0] n9_I_22; // @[Top.scala 41:20]
  wire [7:0] n9_I_23; // @[Top.scala 41:20]
  wire [7:0] n9_I_24; // @[Top.scala 41:20]
  wire [7:0] n9_I_25; // @[Top.scala 41:20]
  wire [7:0] n9_I_26; // @[Top.scala 41:20]
  wire [7:0] n9_I_27; // @[Top.scala 41:20]
  wire [7:0] n9_I_28; // @[Top.scala 41:20]
  wire [7:0] n9_I_29; // @[Top.scala 41:20]
  wire [7:0] n9_I_30; // @[Top.scala 41:20]
  wire [7:0] n9_I_31; // @[Top.scala 41:20]
  wire [7:0] n9_I_32; // @[Top.scala 41:20]
  wire [7:0] n9_I_33; // @[Top.scala 41:20]
  wire [7:0] n9_I_34; // @[Top.scala 41:20]
  wire [7:0] n9_I_35; // @[Top.scala 41:20]
  wire [7:0] n9_I_36; // @[Top.scala 41:20]
  wire [7:0] n9_I_37; // @[Top.scala 41:20]
  wire [7:0] n9_I_38; // @[Top.scala 41:20]
  wire [7:0] n9_I_39; // @[Top.scala 41:20]
  wire [7:0] n9_I_40; // @[Top.scala 41:20]
  wire [7:0] n9_I_41; // @[Top.scala 41:20]
  wire [7:0] n9_I_42; // @[Top.scala 41:20]
  wire [7:0] n9_I_43; // @[Top.scala 41:20]
  wire [7:0] n9_I_44; // @[Top.scala 41:20]
  wire [7:0] n9_I_45; // @[Top.scala 41:20]
  wire [7:0] n9_I_46; // @[Top.scala 41:20]
  wire [7:0] n9_I_47; // @[Top.scala 41:20]
  wire [7:0] n9_I_48; // @[Top.scala 41:20]
  wire [7:0] n9_I_49; // @[Top.scala 41:20]
  wire [7:0] n9_I_50; // @[Top.scala 41:20]
  wire [7:0] n9_I_51; // @[Top.scala 41:20]
  wire [7:0] n9_I_52; // @[Top.scala 41:20]
  wire [7:0] n9_I_53; // @[Top.scala 41:20]
  wire [7:0] n9_I_54; // @[Top.scala 41:20]
  wire [7:0] n9_I_55; // @[Top.scala 41:20]
  wire [7:0] n9_I_56; // @[Top.scala 41:20]
  wire [7:0] n9_I_57; // @[Top.scala 41:20]
  wire [7:0] n9_I_58; // @[Top.scala 41:20]
  wire [7:0] n9_I_59; // @[Top.scala 41:20]
  wire [7:0] n9_I_60; // @[Top.scala 41:20]
  wire [7:0] n9_I_61; // @[Top.scala 41:20]
  wire [7:0] n9_I_62; // @[Top.scala 41:20]
  wire [7:0] n9_I_63; // @[Top.scala 41:20]
  wire [7:0] n9_I_64; // @[Top.scala 41:20]
  wire [7:0] n9_I_65; // @[Top.scala 41:20]
  wire [7:0] n9_I_66; // @[Top.scala 41:20]
  wire [7:0] n9_I_67; // @[Top.scala 41:20]
  wire [7:0] n9_I_68; // @[Top.scala 41:20]
  wire [7:0] n9_I_69; // @[Top.scala 41:20]
  wire [7:0] n9_I_70; // @[Top.scala 41:20]
  wire [7:0] n9_I_71; // @[Top.scala 41:20]
  wire [7:0] n9_I_72; // @[Top.scala 41:20]
  wire [7:0] n9_I_73; // @[Top.scala 41:20]
  wire [7:0] n9_I_74; // @[Top.scala 41:20]
  wire [7:0] n9_I_75; // @[Top.scala 41:20]
  wire [7:0] n9_I_76; // @[Top.scala 41:20]
  wire [7:0] n9_I_77; // @[Top.scala 41:20]
  wire [7:0] n9_I_78; // @[Top.scala 41:20]
  wire [7:0] n9_I_79; // @[Top.scala 41:20]
  wire [7:0] n9_I_80; // @[Top.scala 41:20]
  wire [7:0] n9_I_81; // @[Top.scala 41:20]
  wire [7:0] n9_I_82; // @[Top.scala 41:20]
  wire [7:0] n9_I_83; // @[Top.scala 41:20]
  wire [7:0] n9_I_84; // @[Top.scala 41:20]
  wire [7:0] n9_I_85; // @[Top.scala 41:20]
  wire [7:0] n9_I_86; // @[Top.scala 41:20]
  wire [7:0] n9_I_87; // @[Top.scala 41:20]
  wire [7:0] n9_I_88; // @[Top.scala 41:20]
  wire [7:0] n9_I_89; // @[Top.scala 41:20]
  wire [7:0] n9_I_90; // @[Top.scala 41:20]
  wire [7:0] n9_I_91; // @[Top.scala 41:20]
  wire [7:0] n9_I_92; // @[Top.scala 41:20]
  wire [7:0] n9_I_93; // @[Top.scala 41:20]
  wire [7:0] n9_I_94; // @[Top.scala 41:20]
  wire [7:0] n9_I_95; // @[Top.scala 41:20]
  wire [7:0] n9_I_96; // @[Top.scala 41:20]
  wire [7:0] n9_I_97; // @[Top.scala 41:20]
  wire [7:0] n9_I_98; // @[Top.scala 41:20]
  wire [7:0] n9_I_99; // @[Top.scala 41:20]
  wire [7:0] n9_I_100; // @[Top.scala 41:20]
  wire [7:0] n9_I_101; // @[Top.scala 41:20]
  wire [7:0] n9_I_102; // @[Top.scala 41:20]
  wire [7:0] n9_I_103; // @[Top.scala 41:20]
  wire [7:0] n9_I_104; // @[Top.scala 41:20]
  wire [7:0] n9_I_105; // @[Top.scala 41:20]
  wire [7:0] n9_I_106; // @[Top.scala 41:20]
  wire [7:0] n9_I_107; // @[Top.scala 41:20]
  wire [7:0] n9_I_108; // @[Top.scala 41:20]
  wire [7:0] n9_I_109; // @[Top.scala 41:20]
  wire [7:0] n9_I_110; // @[Top.scala 41:20]
  wire [7:0] n9_I_111; // @[Top.scala 41:20]
  wire [7:0] n9_I_112; // @[Top.scala 41:20]
  wire [7:0] n9_I_113; // @[Top.scala 41:20]
  wire [7:0] n9_I_114; // @[Top.scala 41:20]
  wire [7:0] n9_I_115; // @[Top.scala 41:20]
  wire [7:0] n9_I_116; // @[Top.scala 41:20]
  wire [7:0] n9_I_117; // @[Top.scala 41:20]
  wire [7:0] n9_I_118; // @[Top.scala 41:20]
  wire [7:0] n9_I_119; // @[Top.scala 41:20]
  wire [7:0] n9_I_120; // @[Top.scala 41:20]
  wire [7:0] n9_I_121; // @[Top.scala 41:20]
  wire [7:0] n9_I_122; // @[Top.scala 41:20]
  wire [7:0] n9_I_123; // @[Top.scala 41:20]
  wire [7:0] n9_I_124; // @[Top.scala 41:20]
  wire [7:0] n9_I_125; // @[Top.scala 41:20]
  wire [7:0] n9_I_126; // @[Top.scala 41:20]
  wire [7:0] n9_I_127; // @[Top.scala 41:20]
  wire [7:0] n9_I_128; // @[Top.scala 41:20]
  wire [7:0] n9_I_129; // @[Top.scala 41:20]
  wire [7:0] n9_I_130; // @[Top.scala 41:20]
  wire [7:0] n9_I_131; // @[Top.scala 41:20]
  wire [7:0] n9_I_132; // @[Top.scala 41:20]
  wire [7:0] n9_I_133; // @[Top.scala 41:20]
  wire [7:0] n9_I_134; // @[Top.scala 41:20]
  wire [7:0] n9_I_135; // @[Top.scala 41:20]
  wire [7:0] n9_I_136; // @[Top.scala 41:20]
  wire [7:0] n9_I_137; // @[Top.scala 41:20]
  wire [7:0] n9_I_138; // @[Top.scala 41:20]
  wire [7:0] n9_I_139; // @[Top.scala 41:20]
  wire [7:0] n9_I_140; // @[Top.scala 41:20]
  wire [7:0] n9_I_141; // @[Top.scala 41:20]
  wire [7:0] n9_I_142; // @[Top.scala 41:20]
  wire [7:0] n9_I_143; // @[Top.scala 41:20]
  wire [7:0] n9_I_144; // @[Top.scala 41:20]
  wire [7:0] n9_I_145; // @[Top.scala 41:20]
  wire [7:0] n9_I_146; // @[Top.scala 41:20]
  wire [7:0] n9_I_147; // @[Top.scala 41:20]
  wire [7:0] n9_I_148; // @[Top.scala 41:20]
  wire [7:0] n9_I_149; // @[Top.scala 41:20]
  wire [7:0] n9_I_150; // @[Top.scala 41:20]
  wire [7:0] n9_I_151; // @[Top.scala 41:20]
  wire [7:0] n9_I_152; // @[Top.scala 41:20]
  wire [7:0] n9_I_153; // @[Top.scala 41:20]
  wire [7:0] n9_I_154; // @[Top.scala 41:20]
  wire [7:0] n9_I_155; // @[Top.scala 41:20]
  wire [7:0] n9_I_156; // @[Top.scala 41:20]
  wire [7:0] n9_I_157; // @[Top.scala 41:20]
  wire [7:0] n9_I_158; // @[Top.scala 41:20]
  wire [7:0] n9_I_159; // @[Top.scala 41:20]
  wire [7:0] n9_I_160; // @[Top.scala 41:20]
  wire [7:0] n9_I_161; // @[Top.scala 41:20]
  wire [7:0] n9_I_162; // @[Top.scala 41:20]
  wire [7:0] n9_I_163; // @[Top.scala 41:20]
  wire [7:0] n9_I_164; // @[Top.scala 41:20]
  wire [7:0] n9_I_165; // @[Top.scala 41:20]
  wire [7:0] n9_I_166; // @[Top.scala 41:20]
  wire [7:0] n9_I_167; // @[Top.scala 41:20]
  wire [7:0] n9_I_168; // @[Top.scala 41:20]
  wire [7:0] n9_I_169; // @[Top.scala 41:20]
  wire [7:0] n9_I_170; // @[Top.scala 41:20]
  wire [7:0] n9_I_171; // @[Top.scala 41:20]
  wire [7:0] n9_I_172; // @[Top.scala 41:20]
  wire [7:0] n9_I_173; // @[Top.scala 41:20]
  wire [7:0] n9_I_174; // @[Top.scala 41:20]
  wire [7:0] n9_I_175; // @[Top.scala 41:20]
  wire [7:0] n9_I_176; // @[Top.scala 41:20]
  wire [7:0] n9_I_177; // @[Top.scala 41:20]
  wire [7:0] n9_I_178; // @[Top.scala 41:20]
  wire [7:0] n9_I_179; // @[Top.scala 41:20]
  wire [7:0] n9_I_180; // @[Top.scala 41:20]
  wire [7:0] n9_I_181; // @[Top.scala 41:20]
  wire [7:0] n9_I_182; // @[Top.scala 41:20]
  wire [7:0] n9_I_183; // @[Top.scala 41:20]
  wire [7:0] n9_I_184; // @[Top.scala 41:20]
  wire [7:0] n9_I_185; // @[Top.scala 41:20]
  wire [7:0] n9_I_186; // @[Top.scala 41:20]
  wire [7:0] n9_I_187; // @[Top.scala 41:20]
  wire [7:0] n9_I_188; // @[Top.scala 41:20]
  wire [7:0] n9_I_189; // @[Top.scala 41:20]
  wire [7:0] n9_I_190; // @[Top.scala 41:20]
  wire [7:0] n9_I_191; // @[Top.scala 41:20]
  wire [7:0] n9_I_192; // @[Top.scala 41:20]
  wire [7:0] n9_I_193; // @[Top.scala 41:20]
  wire [7:0] n9_I_194; // @[Top.scala 41:20]
  wire [7:0] n9_I_195; // @[Top.scala 41:20]
  wire [7:0] n9_I_196; // @[Top.scala 41:20]
  wire [7:0] n9_I_197; // @[Top.scala 41:20]
  wire [7:0] n9_I_198; // @[Top.scala 41:20]
  wire [7:0] n9_I_199; // @[Top.scala 41:20]
  wire [7:0] n9_O_0; // @[Top.scala 41:20]
  wire [7:0] n9_O_1; // @[Top.scala 41:20]
  wire [7:0] n9_O_2; // @[Top.scala 41:20]
  wire [7:0] n9_O_3; // @[Top.scala 41:20]
  wire [7:0] n9_O_4; // @[Top.scala 41:20]
  wire [7:0] n9_O_5; // @[Top.scala 41:20]
  wire [7:0] n9_O_6; // @[Top.scala 41:20]
  wire [7:0] n9_O_7; // @[Top.scala 41:20]
  wire [7:0] n9_O_8; // @[Top.scala 41:20]
  wire [7:0] n9_O_9; // @[Top.scala 41:20]
  wire [7:0] n9_O_10; // @[Top.scala 41:20]
  wire [7:0] n9_O_11; // @[Top.scala 41:20]
  wire [7:0] n9_O_12; // @[Top.scala 41:20]
  wire [7:0] n9_O_13; // @[Top.scala 41:20]
  wire [7:0] n9_O_14; // @[Top.scala 41:20]
  wire [7:0] n9_O_15; // @[Top.scala 41:20]
  wire [7:0] n9_O_16; // @[Top.scala 41:20]
  wire [7:0] n9_O_17; // @[Top.scala 41:20]
  wire [7:0] n9_O_18; // @[Top.scala 41:20]
  wire [7:0] n9_O_19; // @[Top.scala 41:20]
  wire [7:0] n9_O_20; // @[Top.scala 41:20]
  wire [7:0] n9_O_21; // @[Top.scala 41:20]
  wire [7:0] n9_O_22; // @[Top.scala 41:20]
  wire [7:0] n9_O_23; // @[Top.scala 41:20]
  wire [7:0] n9_O_24; // @[Top.scala 41:20]
  wire [7:0] n9_O_25; // @[Top.scala 41:20]
  wire [7:0] n9_O_26; // @[Top.scala 41:20]
  wire [7:0] n9_O_27; // @[Top.scala 41:20]
  wire [7:0] n9_O_28; // @[Top.scala 41:20]
  wire [7:0] n9_O_29; // @[Top.scala 41:20]
  wire [7:0] n9_O_30; // @[Top.scala 41:20]
  wire [7:0] n9_O_31; // @[Top.scala 41:20]
  wire [7:0] n9_O_32; // @[Top.scala 41:20]
  wire [7:0] n9_O_33; // @[Top.scala 41:20]
  wire [7:0] n9_O_34; // @[Top.scala 41:20]
  wire [7:0] n9_O_35; // @[Top.scala 41:20]
  wire [7:0] n9_O_36; // @[Top.scala 41:20]
  wire [7:0] n9_O_37; // @[Top.scala 41:20]
  wire [7:0] n9_O_38; // @[Top.scala 41:20]
  wire [7:0] n9_O_39; // @[Top.scala 41:20]
  wire [7:0] n9_O_40; // @[Top.scala 41:20]
  wire [7:0] n9_O_41; // @[Top.scala 41:20]
  wire [7:0] n9_O_42; // @[Top.scala 41:20]
  wire [7:0] n9_O_43; // @[Top.scala 41:20]
  wire [7:0] n9_O_44; // @[Top.scala 41:20]
  wire [7:0] n9_O_45; // @[Top.scala 41:20]
  wire [7:0] n9_O_46; // @[Top.scala 41:20]
  wire [7:0] n9_O_47; // @[Top.scala 41:20]
  wire [7:0] n9_O_48; // @[Top.scala 41:20]
  wire [7:0] n9_O_49; // @[Top.scala 41:20]
  wire [7:0] n9_O_50; // @[Top.scala 41:20]
  wire [7:0] n9_O_51; // @[Top.scala 41:20]
  wire [7:0] n9_O_52; // @[Top.scala 41:20]
  wire [7:0] n9_O_53; // @[Top.scala 41:20]
  wire [7:0] n9_O_54; // @[Top.scala 41:20]
  wire [7:0] n9_O_55; // @[Top.scala 41:20]
  wire [7:0] n9_O_56; // @[Top.scala 41:20]
  wire [7:0] n9_O_57; // @[Top.scala 41:20]
  wire [7:0] n9_O_58; // @[Top.scala 41:20]
  wire [7:0] n9_O_59; // @[Top.scala 41:20]
  wire [7:0] n9_O_60; // @[Top.scala 41:20]
  wire [7:0] n9_O_61; // @[Top.scala 41:20]
  wire [7:0] n9_O_62; // @[Top.scala 41:20]
  wire [7:0] n9_O_63; // @[Top.scala 41:20]
  wire [7:0] n9_O_64; // @[Top.scala 41:20]
  wire [7:0] n9_O_65; // @[Top.scala 41:20]
  wire [7:0] n9_O_66; // @[Top.scala 41:20]
  wire [7:0] n9_O_67; // @[Top.scala 41:20]
  wire [7:0] n9_O_68; // @[Top.scala 41:20]
  wire [7:0] n9_O_69; // @[Top.scala 41:20]
  wire [7:0] n9_O_70; // @[Top.scala 41:20]
  wire [7:0] n9_O_71; // @[Top.scala 41:20]
  wire [7:0] n9_O_72; // @[Top.scala 41:20]
  wire [7:0] n9_O_73; // @[Top.scala 41:20]
  wire [7:0] n9_O_74; // @[Top.scala 41:20]
  wire [7:0] n9_O_75; // @[Top.scala 41:20]
  wire [7:0] n9_O_76; // @[Top.scala 41:20]
  wire [7:0] n9_O_77; // @[Top.scala 41:20]
  wire [7:0] n9_O_78; // @[Top.scala 41:20]
  wire [7:0] n9_O_79; // @[Top.scala 41:20]
  wire [7:0] n9_O_80; // @[Top.scala 41:20]
  wire [7:0] n9_O_81; // @[Top.scala 41:20]
  wire [7:0] n9_O_82; // @[Top.scala 41:20]
  wire [7:0] n9_O_83; // @[Top.scala 41:20]
  wire [7:0] n9_O_84; // @[Top.scala 41:20]
  wire [7:0] n9_O_85; // @[Top.scala 41:20]
  wire [7:0] n9_O_86; // @[Top.scala 41:20]
  wire [7:0] n9_O_87; // @[Top.scala 41:20]
  wire [7:0] n9_O_88; // @[Top.scala 41:20]
  wire [7:0] n9_O_89; // @[Top.scala 41:20]
  wire [7:0] n9_O_90; // @[Top.scala 41:20]
  wire [7:0] n9_O_91; // @[Top.scala 41:20]
  wire [7:0] n9_O_92; // @[Top.scala 41:20]
  wire [7:0] n9_O_93; // @[Top.scala 41:20]
  wire [7:0] n9_O_94; // @[Top.scala 41:20]
  wire [7:0] n9_O_95; // @[Top.scala 41:20]
  wire [7:0] n9_O_96; // @[Top.scala 41:20]
  wire [7:0] n9_O_97; // @[Top.scala 41:20]
  wire [7:0] n9_O_98; // @[Top.scala 41:20]
  wire [7:0] n9_O_99; // @[Top.scala 41:20]
  wire [7:0] n9_O_100; // @[Top.scala 41:20]
  wire [7:0] n9_O_101; // @[Top.scala 41:20]
  wire [7:0] n9_O_102; // @[Top.scala 41:20]
  wire [7:0] n9_O_103; // @[Top.scala 41:20]
  wire [7:0] n9_O_104; // @[Top.scala 41:20]
  wire [7:0] n9_O_105; // @[Top.scala 41:20]
  wire [7:0] n9_O_106; // @[Top.scala 41:20]
  wire [7:0] n9_O_107; // @[Top.scala 41:20]
  wire [7:0] n9_O_108; // @[Top.scala 41:20]
  wire [7:0] n9_O_109; // @[Top.scala 41:20]
  wire [7:0] n9_O_110; // @[Top.scala 41:20]
  wire [7:0] n9_O_111; // @[Top.scala 41:20]
  wire [7:0] n9_O_112; // @[Top.scala 41:20]
  wire [7:0] n9_O_113; // @[Top.scala 41:20]
  wire [7:0] n9_O_114; // @[Top.scala 41:20]
  wire [7:0] n9_O_115; // @[Top.scala 41:20]
  wire [7:0] n9_O_116; // @[Top.scala 41:20]
  wire [7:0] n9_O_117; // @[Top.scala 41:20]
  wire [7:0] n9_O_118; // @[Top.scala 41:20]
  wire [7:0] n9_O_119; // @[Top.scala 41:20]
  wire [7:0] n9_O_120; // @[Top.scala 41:20]
  wire [7:0] n9_O_121; // @[Top.scala 41:20]
  wire [7:0] n9_O_122; // @[Top.scala 41:20]
  wire [7:0] n9_O_123; // @[Top.scala 41:20]
  wire [7:0] n9_O_124; // @[Top.scala 41:20]
  wire [7:0] n9_O_125; // @[Top.scala 41:20]
  wire [7:0] n9_O_126; // @[Top.scala 41:20]
  wire [7:0] n9_O_127; // @[Top.scala 41:20]
  wire [7:0] n9_O_128; // @[Top.scala 41:20]
  wire [7:0] n9_O_129; // @[Top.scala 41:20]
  wire [7:0] n9_O_130; // @[Top.scala 41:20]
  wire [7:0] n9_O_131; // @[Top.scala 41:20]
  wire [7:0] n9_O_132; // @[Top.scala 41:20]
  wire [7:0] n9_O_133; // @[Top.scala 41:20]
  wire [7:0] n9_O_134; // @[Top.scala 41:20]
  wire [7:0] n9_O_135; // @[Top.scala 41:20]
  wire [7:0] n9_O_136; // @[Top.scala 41:20]
  wire [7:0] n9_O_137; // @[Top.scala 41:20]
  wire [7:0] n9_O_138; // @[Top.scala 41:20]
  wire [7:0] n9_O_139; // @[Top.scala 41:20]
  wire [7:0] n9_O_140; // @[Top.scala 41:20]
  wire [7:0] n9_O_141; // @[Top.scala 41:20]
  wire [7:0] n9_O_142; // @[Top.scala 41:20]
  wire [7:0] n9_O_143; // @[Top.scala 41:20]
  wire [7:0] n9_O_144; // @[Top.scala 41:20]
  wire [7:0] n9_O_145; // @[Top.scala 41:20]
  wire [7:0] n9_O_146; // @[Top.scala 41:20]
  wire [7:0] n9_O_147; // @[Top.scala 41:20]
  wire [7:0] n9_O_148; // @[Top.scala 41:20]
  wire [7:0] n9_O_149; // @[Top.scala 41:20]
  wire [7:0] n9_O_150; // @[Top.scala 41:20]
  wire [7:0] n9_O_151; // @[Top.scala 41:20]
  wire [7:0] n9_O_152; // @[Top.scala 41:20]
  wire [7:0] n9_O_153; // @[Top.scala 41:20]
  wire [7:0] n9_O_154; // @[Top.scala 41:20]
  wire [7:0] n9_O_155; // @[Top.scala 41:20]
  wire [7:0] n9_O_156; // @[Top.scala 41:20]
  wire [7:0] n9_O_157; // @[Top.scala 41:20]
  wire [7:0] n9_O_158; // @[Top.scala 41:20]
  wire [7:0] n9_O_159; // @[Top.scala 41:20]
  wire [7:0] n9_O_160; // @[Top.scala 41:20]
  wire [7:0] n9_O_161; // @[Top.scala 41:20]
  wire [7:0] n9_O_162; // @[Top.scala 41:20]
  wire [7:0] n9_O_163; // @[Top.scala 41:20]
  wire [7:0] n9_O_164; // @[Top.scala 41:20]
  wire [7:0] n9_O_165; // @[Top.scala 41:20]
  wire [7:0] n9_O_166; // @[Top.scala 41:20]
  wire [7:0] n9_O_167; // @[Top.scala 41:20]
  wire [7:0] n9_O_168; // @[Top.scala 41:20]
  wire [7:0] n9_O_169; // @[Top.scala 41:20]
  wire [7:0] n9_O_170; // @[Top.scala 41:20]
  wire [7:0] n9_O_171; // @[Top.scala 41:20]
  wire [7:0] n9_O_172; // @[Top.scala 41:20]
  wire [7:0] n9_O_173; // @[Top.scala 41:20]
  wire [7:0] n9_O_174; // @[Top.scala 41:20]
  wire [7:0] n9_O_175; // @[Top.scala 41:20]
  wire [7:0] n9_O_176; // @[Top.scala 41:20]
  wire [7:0] n9_O_177; // @[Top.scala 41:20]
  wire [7:0] n9_O_178; // @[Top.scala 41:20]
  wire [7:0] n9_O_179; // @[Top.scala 41:20]
  wire [7:0] n9_O_180; // @[Top.scala 41:20]
  wire [7:0] n9_O_181; // @[Top.scala 41:20]
  wire [7:0] n9_O_182; // @[Top.scala 41:20]
  wire [7:0] n9_O_183; // @[Top.scala 41:20]
  wire [7:0] n9_O_184; // @[Top.scala 41:20]
  wire [7:0] n9_O_185; // @[Top.scala 41:20]
  wire [7:0] n9_O_186; // @[Top.scala 41:20]
  wire [7:0] n9_O_187; // @[Top.scala 41:20]
  wire [7:0] n9_O_188; // @[Top.scala 41:20]
  wire [7:0] n9_O_189; // @[Top.scala 41:20]
  wire [7:0] n9_O_190; // @[Top.scala 41:20]
  wire [7:0] n9_O_191; // @[Top.scala 41:20]
  wire [7:0] n9_O_192; // @[Top.scala 41:20]
  wire [7:0] n9_O_193; // @[Top.scala 41:20]
  wire [7:0] n9_O_194; // @[Top.scala 41:20]
  wire [7:0] n9_O_195; // @[Top.scala 41:20]
  wire [7:0] n9_O_196; // @[Top.scala 41:20]
  wire [7:0] n9_O_197; // @[Top.scala 41:20]
  wire [7:0] n9_O_198; // @[Top.scala 41:20]
  wire [7:0] n9_O_199; // @[Top.scala 41:20]
  wire  n10_clock; // @[Top.scala 44:21]
  wire  n10_reset; // @[Top.scala 44:21]
  wire  n10_valid_up; // @[Top.scala 44:21]
  wire  n10_valid_down; // @[Top.scala 44:21]
  wire [7:0] n10_I_0; // @[Top.scala 44:21]
  wire [7:0] n10_I_1; // @[Top.scala 44:21]
  wire [7:0] n10_I_2; // @[Top.scala 44:21]
  wire [7:0] n10_I_3; // @[Top.scala 44:21]
  wire [7:0] n10_I_4; // @[Top.scala 44:21]
  wire [7:0] n10_I_5; // @[Top.scala 44:21]
  wire [7:0] n10_I_6; // @[Top.scala 44:21]
  wire [7:0] n10_I_7; // @[Top.scala 44:21]
  wire [7:0] n10_I_8; // @[Top.scala 44:21]
  wire [7:0] n10_I_9; // @[Top.scala 44:21]
  wire [7:0] n10_I_10; // @[Top.scala 44:21]
  wire [7:0] n10_I_11; // @[Top.scala 44:21]
  wire [7:0] n10_I_12; // @[Top.scala 44:21]
  wire [7:0] n10_I_13; // @[Top.scala 44:21]
  wire [7:0] n10_I_14; // @[Top.scala 44:21]
  wire [7:0] n10_I_15; // @[Top.scala 44:21]
  wire [7:0] n10_I_16; // @[Top.scala 44:21]
  wire [7:0] n10_I_17; // @[Top.scala 44:21]
  wire [7:0] n10_I_18; // @[Top.scala 44:21]
  wire [7:0] n10_I_19; // @[Top.scala 44:21]
  wire [7:0] n10_I_20; // @[Top.scala 44:21]
  wire [7:0] n10_I_21; // @[Top.scala 44:21]
  wire [7:0] n10_I_22; // @[Top.scala 44:21]
  wire [7:0] n10_I_23; // @[Top.scala 44:21]
  wire [7:0] n10_I_24; // @[Top.scala 44:21]
  wire [7:0] n10_I_25; // @[Top.scala 44:21]
  wire [7:0] n10_I_26; // @[Top.scala 44:21]
  wire [7:0] n10_I_27; // @[Top.scala 44:21]
  wire [7:0] n10_I_28; // @[Top.scala 44:21]
  wire [7:0] n10_I_29; // @[Top.scala 44:21]
  wire [7:0] n10_I_30; // @[Top.scala 44:21]
  wire [7:0] n10_I_31; // @[Top.scala 44:21]
  wire [7:0] n10_I_32; // @[Top.scala 44:21]
  wire [7:0] n10_I_33; // @[Top.scala 44:21]
  wire [7:0] n10_I_34; // @[Top.scala 44:21]
  wire [7:0] n10_I_35; // @[Top.scala 44:21]
  wire [7:0] n10_I_36; // @[Top.scala 44:21]
  wire [7:0] n10_I_37; // @[Top.scala 44:21]
  wire [7:0] n10_I_38; // @[Top.scala 44:21]
  wire [7:0] n10_I_39; // @[Top.scala 44:21]
  wire [7:0] n10_I_40; // @[Top.scala 44:21]
  wire [7:0] n10_I_41; // @[Top.scala 44:21]
  wire [7:0] n10_I_42; // @[Top.scala 44:21]
  wire [7:0] n10_I_43; // @[Top.scala 44:21]
  wire [7:0] n10_I_44; // @[Top.scala 44:21]
  wire [7:0] n10_I_45; // @[Top.scala 44:21]
  wire [7:0] n10_I_46; // @[Top.scala 44:21]
  wire [7:0] n10_I_47; // @[Top.scala 44:21]
  wire [7:0] n10_I_48; // @[Top.scala 44:21]
  wire [7:0] n10_I_49; // @[Top.scala 44:21]
  wire [7:0] n10_I_50; // @[Top.scala 44:21]
  wire [7:0] n10_I_51; // @[Top.scala 44:21]
  wire [7:0] n10_I_52; // @[Top.scala 44:21]
  wire [7:0] n10_I_53; // @[Top.scala 44:21]
  wire [7:0] n10_I_54; // @[Top.scala 44:21]
  wire [7:0] n10_I_55; // @[Top.scala 44:21]
  wire [7:0] n10_I_56; // @[Top.scala 44:21]
  wire [7:0] n10_I_57; // @[Top.scala 44:21]
  wire [7:0] n10_I_58; // @[Top.scala 44:21]
  wire [7:0] n10_I_59; // @[Top.scala 44:21]
  wire [7:0] n10_I_60; // @[Top.scala 44:21]
  wire [7:0] n10_I_61; // @[Top.scala 44:21]
  wire [7:0] n10_I_62; // @[Top.scala 44:21]
  wire [7:0] n10_I_63; // @[Top.scala 44:21]
  wire [7:0] n10_I_64; // @[Top.scala 44:21]
  wire [7:0] n10_I_65; // @[Top.scala 44:21]
  wire [7:0] n10_I_66; // @[Top.scala 44:21]
  wire [7:0] n10_I_67; // @[Top.scala 44:21]
  wire [7:0] n10_I_68; // @[Top.scala 44:21]
  wire [7:0] n10_I_69; // @[Top.scala 44:21]
  wire [7:0] n10_I_70; // @[Top.scala 44:21]
  wire [7:0] n10_I_71; // @[Top.scala 44:21]
  wire [7:0] n10_I_72; // @[Top.scala 44:21]
  wire [7:0] n10_I_73; // @[Top.scala 44:21]
  wire [7:0] n10_I_74; // @[Top.scala 44:21]
  wire [7:0] n10_I_75; // @[Top.scala 44:21]
  wire [7:0] n10_I_76; // @[Top.scala 44:21]
  wire [7:0] n10_I_77; // @[Top.scala 44:21]
  wire [7:0] n10_I_78; // @[Top.scala 44:21]
  wire [7:0] n10_I_79; // @[Top.scala 44:21]
  wire [7:0] n10_I_80; // @[Top.scala 44:21]
  wire [7:0] n10_I_81; // @[Top.scala 44:21]
  wire [7:0] n10_I_82; // @[Top.scala 44:21]
  wire [7:0] n10_I_83; // @[Top.scala 44:21]
  wire [7:0] n10_I_84; // @[Top.scala 44:21]
  wire [7:0] n10_I_85; // @[Top.scala 44:21]
  wire [7:0] n10_I_86; // @[Top.scala 44:21]
  wire [7:0] n10_I_87; // @[Top.scala 44:21]
  wire [7:0] n10_I_88; // @[Top.scala 44:21]
  wire [7:0] n10_I_89; // @[Top.scala 44:21]
  wire [7:0] n10_I_90; // @[Top.scala 44:21]
  wire [7:0] n10_I_91; // @[Top.scala 44:21]
  wire [7:0] n10_I_92; // @[Top.scala 44:21]
  wire [7:0] n10_I_93; // @[Top.scala 44:21]
  wire [7:0] n10_I_94; // @[Top.scala 44:21]
  wire [7:0] n10_I_95; // @[Top.scala 44:21]
  wire [7:0] n10_I_96; // @[Top.scala 44:21]
  wire [7:0] n10_I_97; // @[Top.scala 44:21]
  wire [7:0] n10_I_98; // @[Top.scala 44:21]
  wire [7:0] n10_I_99; // @[Top.scala 44:21]
  wire [7:0] n10_I_100; // @[Top.scala 44:21]
  wire [7:0] n10_I_101; // @[Top.scala 44:21]
  wire [7:0] n10_I_102; // @[Top.scala 44:21]
  wire [7:0] n10_I_103; // @[Top.scala 44:21]
  wire [7:0] n10_I_104; // @[Top.scala 44:21]
  wire [7:0] n10_I_105; // @[Top.scala 44:21]
  wire [7:0] n10_I_106; // @[Top.scala 44:21]
  wire [7:0] n10_I_107; // @[Top.scala 44:21]
  wire [7:0] n10_I_108; // @[Top.scala 44:21]
  wire [7:0] n10_I_109; // @[Top.scala 44:21]
  wire [7:0] n10_I_110; // @[Top.scala 44:21]
  wire [7:0] n10_I_111; // @[Top.scala 44:21]
  wire [7:0] n10_I_112; // @[Top.scala 44:21]
  wire [7:0] n10_I_113; // @[Top.scala 44:21]
  wire [7:0] n10_I_114; // @[Top.scala 44:21]
  wire [7:0] n10_I_115; // @[Top.scala 44:21]
  wire [7:0] n10_I_116; // @[Top.scala 44:21]
  wire [7:0] n10_I_117; // @[Top.scala 44:21]
  wire [7:0] n10_I_118; // @[Top.scala 44:21]
  wire [7:0] n10_I_119; // @[Top.scala 44:21]
  wire [7:0] n10_I_120; // @[Top.scala 44:21]
  wire [7:0] n10_I_121; // @[Top.scala 44:21]
  wire [7:0] n10_I_122; // @[Top.scala 44:21]
  wire [7:0] n10_I_123; // @[Top.scala 44:21]
  wire [7:0] n10_I_124; // @[Top.scala 44:21]
  wire [7:0] n10_I_125; // @[Top.scala 44:21]
  wire [7:0] n10_I_126; // @[Top.scala 44:21]
  wire [7:0] n10_I_127; // @[Top.scala 44:21]
  wire [7:0] n10_I_128; // @[Top.scala 44:21]
  wire [7:0] n10_I_129; // @[Top.scala 44:21]
  wire [7:0] n10_I_130; // @[Top.scala 44:21]
  wire [7:0] n10_I_131; // @[Top.scala 44:21]
  wire [7:0] n10_I_132; // @[Top.scala 44:21]
  wire [7:0] n10_I_133; // @[Top.scala 44:21]
  wire [7:0] n10_I_134; // @[Top.scala 44:21]
  wire [7:0] n10_I_135; // @[Top.scala 44:21]
  wire [7:0] n10_I_136; // @[Top.scala 44:21]
  wire [7:0] n10_I_137; // @[Top.scala 44:21]
  wire [7:0] n10_I_138; // @[Top.scala 44:21]
  wire [7:0] n10_I_139; // @[Top.scala 44:21]
  wire [7:0] n10_I_140; // @[Top.scala 44:21]
  wire [7:0] n10_I_141; // @[Top.scala 44:21]
  wire [7:0] n10_I_142; // @[Top.scala 44:21]
  wire [7:0] n10_I_143; // @[Top.scala 44:21]
  wire [7:0] n10_I_144; // @[Top.scala 44:21]
  wire [7:0] n10_I_145; // @[Top.scala 44:21]
  wire [7:0] n10_I_146; // @[Top.scala 44:21]
  wire [7:0] n10_I_147; // @[Top.scala 44:21]
  wire [7:0] n10_I_148; // @[Top.scala 44:21]
  wire [7:0] n10_I_149; // @[Top.scala 44:21]
  wire [7:0] n10_I_150; // @[Top.scala 44:21]
  wire [7:0] n10_I_151; // @[Top.scala 44:21]
  wire [7:0] n10_I_152; // @[Top.scala 44:21]
  wire [7:0] n10_I_153; // @[Top.scala 44:21]
  wire [7:0] n10_I_154; // @[Top.scala 44:21]
  wire [7:0] n10_I_155; // @[Top.scala 44:21]
  wire [7:0] n10_I_156; // @[Top.scala 44:21]
  wire [7:0] n10_I_157; // @[Top.scala 44:21]
  wire [7:0] n10_I_158; // @[Top.scala 44:21]
  wire [7:0] n10_I_159; // @[Top.scala 44:21]
  wire [7:0] n10_I_160; // @[Top.scala 44:21]
  wire [7:0] n10_I_161; // @[Top.scala 44:21]
  wire [7:0] n10_I_162; // @[Top.scala 44:21]
  wire [7:0] n10_I_163; // @[Top.scala 44:21]
  wire [7:0] n10_I_164; // @[Top.scala 44:21]
  wire [7:0] n10_I_165; // @[Top.scala 44:21]
  wire [7:0] n10_I_166; // @[Top.scala 44:21]
  wire [7:0] n10_I_167; // @[Top.scala 44:21]
  wire [7:0] n10_I_168; // @[Top.scala 44:21]
  wire [7:0] n10_I_169; // @[Top.scala 44:21]
  wire [7:0] n10_I_170; // @[Top.scala 44:21]
  wire [7:0] n10_I_171; // @[Top.scala 44:21]
  wire [7:0] n10_I_172; // @[Top.scala 44:21]
  wire [7:0] n10_I_173; // @[Top.scala 44:21]
  wire [7:0] n10_I_174; // @[Top.scala 44:21]
  wire [7:0] n10_I_175; // @[Top.scala 44:21]
  wire [7:0] n10_I_176; // @[Top.scala 44:21]
  wire [7:0] n10_I_177; // @[Top.scala 44:21]
  wire [7:0] n10_I_178; // @[Top.scala 44:21]
  wire [7:0] n10_I_179; // @[Top.scala 44:21]
  wire [7:0] n10_I_180; // @[Top.scala 44:21]
  wire [7:0] n10_I_181; // @[Top.scala 44:21]
  wire [7:0] n10_I_182; // @[Top.scala 44:21]
  wire [7:0] n10_I_183; // @[Top.scala 44:21]
  wire [7:0] n10_I_184; // @[Top.scala 44:21]
  wire [7:0] n10_I_185; // @[Top.scala 44:21]
  wire [7:0] n10_I_186; // @[Top.scala 44:21]
  wire [7:0] n10_I_187; // @[Top.scala 44:21]
  wire [7:0] n10_I_188; // @[Top.scala 44:21]
  wire [7:0] n10_I_189; // @[Top.scala 44:21]
  wire [7:0] n10_I_190; // @[Top.scala 44:21]
  wire [7:0] n10_I_191; // @[Top.scala 44:21]
  wire [7:0] n10_I_192; // @[Top.scala 44:21]
  wire [7:0] n10_I_193; // @[Top.scala 44:21]
  wire [7:0] n10_I_194; // @[Top.scala 44:21]
  wire [7:0] n10_I_195; // @[Top.scala 44:21]
  wire [7:0] n10_I_196; // @[Top.scala 44:21]
  wire [7:0] n10_I_197; // @[Top.scala 44:21]
  wire [7:0] n10_I_198; // @[Top.scala 44:21]
  wire [7:0] n10_I_199; // @[Top.scala 44:21]
  wire [7:0] n10_O_0; // @[Top.scala 44:21]
  wire [7:0] n10_O_1; // @[Top.scala 44:21]
  wire [7:0] n10_O_2; // @[Top.scala 44:21]
  wire [7:0] n10_O_3; // @[Top.scala 44:21]
  wire [7:0] n10_O_4; // @[Top.scala 44:21]
  wire [7:0] n10_O_5; // @[Top.scala 44:21]
  wire [7:0] n10_O_6; // @[Top.scala 44:21]
  wire [7:0] n10_O_7; // @[Top.scala 44:21]
  wire [7:0] n10_O_8; // @[Top.scala 44:21]
  wire [7:0] n10_O_9; // @[Top.scala 44:21]
  wire [7:0] n10_O_10; // @[Top.scala 44:21]
  wire [7:0] n10_O_11; // @[Top.scala 44:21]
  wire [7:0] n10_O_12; // @[Top.scala 44:21]
  wire [7:0] n10_O_13; // @[Top.scala 44:21]
  wire [7:0] n10_O_14; // @[Top.scala 44:21]
  wire [7:0] n10_O_15; // @[Top.scala 44:21]
  wire [7:0] n10_O_16; // @[Top.scala 44:21]
  wire [7:0] n10_O_17; // @[Top.scala 44:21]
  wire [7:0] n10_O_18; // @[Top.scala 44:21]
  wire [7:0] n10_O_19; // @[Top.scala 44:21]
  wire [7:0] n10_O_20; // @[Top.scala 44:21]
  wire [7:0] n10_O_21; // @[Top.scala 44:21]
  wire [7:0] n10_O_22; // @[Top.scala 44:21]
  wire [7:0] n10_O_23; // @[Top.scala 44:21]
  wire [7:0] n10_O_24; // @[Top.scala 44:21]
  wire [7:0] n10_O_25; // @[Top.scala 44:21]
  wire [7:0] n10_O_26; // @[Top.scala 44:21]
  wire [7:0] n10_O_27; // @[Top.scala 44:21]
  wire [7:0] n10_O_28; // @[Top.scala 44:21]
  wire [7:0] n10_O_29; // @[Top.scala 44:21]
  wire [7:0] n10_O_30; // @[Top.scala 44:21]
  wire [7:0] n10_O_31; // @[Top.scala 44:21]
  wire [7:0] n10_O_32; // @[Top.scala 44:21]
  wire [7:0] n10_O_33; // @[Top.scala 44:21]
  wire [7:0] n10_O_34; // @[Top.scala 44:21]
  wire [7:0] n10_O_35; // @[Top.scala 44:21]
  wire [7:0] n10_O_36; // @[Top.scala 44:21]
  wire [7:0] n10_O_37; // @[Top.scala 44:21]
  wire [7:0] n10_O_38; // @[Top.scala 44:21]
  wire [7:0] n10_O_39; // @[Top.scala 44:21]
  wire [7:0] n10_O_40; // @[Top.scala 44:21]
  wire [7:0] n10_O_41; // @[Top.scala 44:21]
  wire [7:0] n10_O_42; // @[Top.scala 44:21]
  wire [7:0] n10_O_43; // @[Top.scala 44:21]
  wire [7:0] n10_O_44; // @[Top.scala 44:21]
  wire [7:0] n10_O_45; // @[Top.scala 44:21]
  wire [7:0] n10_O_46; // @[Top.scala 44:21]
  wire [7:0] n10_O_47; // @[Top.scala 44:21]
  wire [7:0] n10_O_48; // @[Top.scala 44:21]
  wire [7:0] n10_O_49; // @[Top.scala 44:21]
  wire [7:0] n10_O_50; // @[Top.scala 44:21]
  wire [7:0] n10_O_51; // @[Top.scala 44:21]
  wire [7:0] n10_O_52; // @[Top.scala 44:21]
  wire [7:0] n10_O_53; // @[Top.scala 44:21]
  wire [7:0] n10_O_54; // @[Top.scala 44:21]
  wire [7:0] n10_O_55; // @[Top.scala 44:21]
  wire [7:0] n10_O_56; // @[Top.scala 44:21]
  wire [7:0] n10_O_57; // @[Top.scala 44:21]
  wire [7:0] n10_O_58; // @[Top.scala 44:21]
  wire [7:0] n10_O_59; // @[Top.scala 44:21]
  wire [7:0] n10_O_60; // @[Top.scala 44:21]
  wire [7:0] n10_O_61; // @[Top.scala 44:21]
  wire [7:0] n10_O_62; // @[Top.scala 44:21]
  wire [7:0] n10_O_63; // @[Top.scala 44:21]
  wire [7:0] n10_O_64; // @[Top.scala 44:21]
  wire [7:0] n10_O_65; // @[Top.scala 44:21]
  wire [7:0] n10_O_66; // @[Top.scala 44:21]
  wire [7:0] n10_O_67; // @[Top.scala 44:21]
  wire [7:0] n10_O_68; // @[Top.scala 44:21]
  wire [7:0] n10_O_69; // @[Top.scala 44:21]
  wire [7:0] n10_O_70; // @[Top.scala 44:21]
  wire [7:0] n10_O_71; // @[Top.scala 44:21]
  wire [7:0] n10_O_72; // @[Top.scala 44:21]
  wire [7:0] n10_O_73; // @[Top.scala 44:21]
  wire [7:0] n10_O_74; // @[Top.scala 44:21]
  wire [7:0] n10_O_75; // @[Top.scala 44:21]
  wire [7:0] n10_O_76; // @[Top.scala 44:21]
  wire [7:0] n10_O_77; // @[Top.scala 44:21]
  wire [7:0] n10_O_78; // @[Top.scala 44:21]
  wire [7:0] n10_O_79; // @[Top.scala 44:21]
  wire [7:0] n10_O_80; // @[Top.scala 44:21]
  wire [7:0] n10_O_81; // @[Top.scala 44:21]
  wire [7:0] n10_O_82; // @[Top.scala 44:21]
  wire [7:0] n10_O_83; // @[Top.scala 44:21]
  wire [7:0] n10_O_84; // @[Top.scala 44:21]
  wire [7:0] n10_O_85; // @[Top.scala 44:21]
  wire [7:0] n10_O_86; // @[Top.scala 44:21]
  wire [7:0] n10_O_87; // @[Top.scala 44:21]
  wire [7:0] n10_O_88; // @[Top.scala 44:21]
  wire [7:0] n10_O_89; // @[Top.scala 44:21]
  wire [7:0] n10_O_90; // @[Top.scala 44:21]
  wire [7:0] n10_O_91; // @[Top.scala 44:21]
  wire [7:0] n10_O_92; // @[Top.scala 44:21]
  wire [7:0] n10_O_93; // @[Top.scala 44:21]
  wire [7:0] n10_O_94; // @[Top.scala 44:21]
  wire [7:0] n10_O_95; // @[Top.scala 44:21]
  wire [7:0] n10_O_96; // @[Top.scala 44:21]
  wire [7:0] n10_O_97; // @[Top.scala 44:21]
  wire [7:0] n10_O_98; // @[Top.scala 44:21]
  wire [7:0] n10_O_99; // @[Top.scala 44:21]
  wire [7:0] n10_O_100; // @[Top.scala 44:21]
  wire [7:0] n10_O_101; // @[Top.scala 44:21]
  wire [7:0] n10_O_102; // @[Top.scala 44:21]
  wire [7:0] n10_O_103; // @[Top.scala 44:21]
  wire [7:0] n10_O_104; // @[Top.scala 44:21]
  wire [7:0] n10_O_105; // @[Top.scala 44:21]
  wire [7:0] n10_O_106; // @[Top.scala 44:21]
  wire [7:0] n10_O_107; // @[Top.scala 44:21]
  wire [7:0] n10_O_108; // @[Top.scala 44:21]
  wire [7:0] n10_O_109; // @[Top.scala 44:21]
  wire [7:0] n10_O_110; // @[Top.scala 44:21]
  wire [7:0] n10_O_111; // @[Top.scala 44:21]
  wire [7:0] n10_O_112; // @[Top.scala 44:21]
  wire [7:0] n10_O_113; // @[Top.scala 44:21]
  wire [7:0] n10_O_114; // @[Top.scala 44:21]
  wire [7:0] n10_O_115; // @[Top.scala 44:21]
  wire [7:0] n10_O_116; // @[Top.scala 44:21]
  wire [7:0] n10_O_117; // @[Top.scala 44:21]
  wire [7:0] n10_O_118; // @[Top.scala 44:21]
  wire [7:0] n10_O_119; // @[Top.scala 44:21]
  wire [7:0] n10_O_120; // @[Top.scala 44:21]
  wire [7:0] n10_O_121; // @[Top.scala 44:21]
  wire [7:0] n10_O_122; // @[Top.scala 44:21]
  wire [7:0] n10_O_123; // @[Top.scala 44:21]
  wire [7:0] n10_O_124; // @[Top.scala 44:21]
  wire [7:0] n10_O_125; // @[Top.scala 44:21]
  wire [7:0] n10_O_126; // @[Top.scala 44:21]
  wire [7:0] n10_O_127; // @[Top.scala 44:21]
  wire [7:0] n10_O_128; // @[Top.scala 44:21]
  wire [7:0] n10_O_129; // @[Top.scala 44:21]
  wire [7:0] n10_O_130; // @[Top.scala 44:21]
  wire [7:0] n10_O_131; // @[Top.scala 44:21]
  wire [7:0] n10_O_132; // @[Top.scala 44:21]
  wire [7:0] n10_O_133; // @[Top.scala 44:21]
  wire [7:0] n10_O_134; // @[Top.scala 44:21]
  wire [7:0] n10_O_135; // @[Top.scala 44:21]
  wire [7:0] n10_O_136; // @[Top.scala 44:21]
  wire [7:0] n10_O_137; // @[Top.scala 44:21]
  wire [7:0] n10_O_138; // @[Top.scala 44:21]
  wire [7:0] n10_O_139; // @[Top.scala 44:21]
  wire [7:0] n10_O_140; // @[Top.scala 44:21]
  wire [7:0] n10_O_141; // @[Top.scala 44:21]
  wire [7:0] n10_O_142; // @[Top.scala 44:21]
  wire [7:0] n10_O_143; // @[Top.scala 44:21]
  wire [7:0] n10_O_144; // @[Top.scala 44:21]
  wire [7:0] n10_O_145; // @[Top.scala 44:21]
  wire [7:0] n10_O_146; // @[Top.scala 44:21]
  wire [7:0] n10_O_147; // @[Top.scala 44:21]
  wire [7:0] n10_O_148; // @[Top.scala 44:21]
  wire [7:0] n10_O_149; // @[Top.scala 44:21]
  wire [7:0] n10_O_150; // @[Top.scala 44:21]
  wire [7:0] n10_O_151; // @[Top.scala 44:21]
  wire [7:0] n10_O_152; // @[Top.scala 44:21]
  wire [7:0] n10_O_153; // @[Top.scala 44:21]
  wire [7:0] n10_O_154; // @[Top.scala 44:21]
  wire [7:0] n10_O_155; // @[Top.scala 44:21]
  wire [7:0] n10_O_156; // @[Top.scala 44:21]
  wire [7:0] n10_O_157; // @[Top.scala 44:21]
  wire [7:0] n10_O_158; // @[Top.scala 44:21]
  wire [7:0] n10_O_159; // @[Top.scala 44:21]
  wire [7:0] n10_O_160; // @[Top.scala 44:21]
  wire [7:0] n10_O_161; // @[Top.scala 44:21]
  wire [7:0] n10_O_162; // @[Top.scala 44:21]
  wire [7:0] n10_O_163; // @[Top.scala 44:21]
  wire [7:0] n10_O_164; // @[Top.scala 44:21]
  wire [7:0] n10_O_165; // @[Top.scala 44:21]
  wire [7:0] n10_O_166; // @[Top.scala 44:21]
  wire [7:0] n10_O_167; // @[Top.scala 44:21]
  wire [7:0] n10_O_168; // @[Top.scala 44:21]
  wire [7:0] n10_O_169; // @[Top.scala 44:21]
  wire [7:0] n10_O_170; // @[Top.scala 44:21]
  wire [7:0] n10_O_171; // @[Top.scala 44:21]
  wire [7:0] n10_O_172; // @[Top.scala 44:21]
  wire [7:0] n10_O_173; // @[Top.scala 44:21]
  wire [7:0] n10_O_174; // @[Top.scala 44:21]
  wire [7:0] n10_O_175; // @[Top.scala 44:21]
  wire [7:0] n10_O_176; // @[Top.scala 44:21]
  wire [7:0] n10_O_177; // @[Top.scala 44:21]
  wire [7:0] n10_O_178; // @[Top.scala 44:21]
  wire [7:0] n10_O_179; // @[Top.scala 44:21]
  wire [7:0] n10_O_180; // @[Top.scala 44:21]
  wire [7:0] n10_O_181; // @[Top.scala 44:21]
  wire [7:0] n10_O_182; // @[Top.scala 44:21]
  wire [7:0] n10_O_183; // @[Top.scala 44:21]
  wire [7:0] n10_O_184; // @[Top.scala 44:21]
  wire [7:0] n10_O_185; // @[Top.scala 44:21]
  wire [7:0] n10_O_186; // @[Top.scala 44:21]
  wire [7:0] n10_O_187; // @[Top.scala 44:21]
  wire [7:0] n10_O_188; // @[Top.scala 44:21]
  wire [7:0] n10_O_189; // @[Top.scala 44:21]
  wire [7:0] n10_O_190; // @[Top.scala 44:21]
  wire [7:0] n10_O_191; // @[Top.scala 44:21]
  wire [7:0] n10_O_192; // @[Top.scala 44:21]
  wire [7:0] n10_O_193; // @[Top.scala 44:21]
  wire [7:0] n10_O_194; // @[Top.scala 44:21]
  wire [7:0] n10_O_195; // @[Top.scala 44:21]
  wire [7:0] n10_O_196; // @[Top.scala 44:21]
  wire [7:0] n10_O_197; // @[Top.scala 44:21]
  wire [7:0] n10_O_198; // @[Top.scala 44:21]
  wire [7:0] n10_O_199; // @[Top.scala 44:21]
  FIFO n1 ( // @[Top.scala 32:20]
    .clock(n1_clock),
    .reset(n1_reset),
    .valid_up(n1_valid_up),
    .valid_down(n1_valid_down),
    .I_0(n1_I_0),
    .I_1(n1_I_1),
    .I_2(n1_I_2),
    .I_3(n1_I_3),
    .I_4(n1_I_4),
    .I_5(n1_I_5),
    .I_6(n1_I_6),
    .I_7(n1_I_7),
    .I_8(n1_I_8),
    .I_9(n1_I_9),
    .I_10(n1_I_10),
    .I_11(n1_I_11),
    .I_12(n1_I_12),
    .I_13(n1_I_13),
    .I_14(n1_I_14),
    .I_15(n1_I_15),
    .I_16(n1_I_16),
    .I_17(n1_I_17),
    .I_18(n1_I_18),
    .I_19(n1_I_19),
    .I_20(n1_I_20),
    .I_21(n1_I_21),
    .I_22(n1_I_22),
    .I_23(n1_I_23),
    .I_24(n1_I_24),
    .I_25(n1_I_25),
    .I_26(n1_I_26),
    .I_27(n1_I_27),
    .I_28(n1_I_28),
    .I_29(n1_I_29),
    .I_30(n1_I_30),
    .I_31(n1_I_31),
    .I_32(n1_I_32),
    .I_33(n1_I_33),
    .I_34(n1_I_34),
    .I_35(n1_I_35),
    .I_36(n1_I_36),
    .I_37(n1_I_37),
    .I_38(n1_I_38),
    .I_39(n1_I_39),
    .I_40(n1_I_40),
    .I_41(n1_I_41),
    .I_42(n1_I_42),
    .I_43(n1_I_43),
    .I_44(n1_I_44),
    .I_45(n1_I_45),
    .I_46(n1_I_46),
    .I_47(n1_I_47),
    .I_48(n1_I_48),
    .I_49(n1_I_49),
    .I_50(n1_I_50),
    .I_51(n1_I_51),
    .I_52(n1_I_52),
    .I_53(n1_I_53),
    .I_54(n1_I_54),
    .I_55(n1_I_55),
    .I_56(n1_I_56),
    .I_57(n1_I_57),
    .I_58(n1_I_58),
    .I_59(n1_I_59),
    .I_60(n1_I_60),
    .I_61(n1_I_61),
    .I_62(n1_I_62),
    .I_63(n1_I_63),
    .I_64(n1_I_64),
    .I_65(n1_I_65),
    .I_66(n1_I_66),
    .I_67(n1_I_67),
    .I_68(n1_I_68),
    .I_69(n1_I_69),
    .I_70(n1_I_70),
    .I_71(n1_I_71),
    .I_72(n1_I_72),
    .I_73(n1_I_73),
    .I_74(n1_I_74),
    .I_75(n1_I_75),
    .I_76(n1_I_76),
    .I_77(n1_I_77),
    .I_78(n1_I_78),
    .I_79(n1_I_79),
    .I_80(n1_I_80),
    .I_81(n1_I_81),
    .I_82(n1_I_82),
    .I_83(n1_I_83),
    .I_84(n1_I_84),
    .I_85(n1_I_85),
    .I_86(n1_I_86),
    .I_87(n1_I_87),
    .I_88(n1_I_88),
    .I_89(n1_I_89),
    .I_90(n1_I_90),
    .I_91(n1_I_91),
    .I_92(n1_I_92),
    .I_93(n1_I_93),
    .I_94(n1_I_94),
    .I_95(n1_I_95),
    .I_96(n1_I_96),
    .I_97(n1_I_97),
    .I_98(n1_I_98),
    .I_99(n1_I_99),
    .I_100(n1_I_100),
    .I_101(n1_I_101),
    .I_102(n1_I_102),
    .I_103(n1_I_103),
    .I_104(n1_I_104),
    .I_105(n1_I_105),
    .I_106(n1_I_106),
    .I_107(n1_I_107),
    .I_108(n1_I_108),
    .I_109(n1_I_109),
    .I_110(n1_I_110),
    .I_111(n1_I_111),
    .I_112(n1_I_112),
    .I_113(n1_I_113),
    .I_114(n1_I_114),
    .I_115(n1_I_115),
    .I_116(n1_I_116),
    .I_117(n1_I_117),
    .I_118(n1_I_118),
    .I_119(n1_I_119),
    .I_120(n1_I_120),
    .I_121(n1_I_121),
    .I_122(n1_I_122),
    .I_123(n1_I_123),
    .I_124(n1_I_124),
    .I_125(n1_I_125),
    .I_126(n1_I_126),
    .I_127(n1_I_127),
    .I_128(n1_I_128),
    .I_129(n1_I_129),
    .I_130(n1_I_130),
    .I_131(n1_I_131),
    .I_132(n1_I_132),
    .I_133(n1_I_133),
    .I_134(n1_I_134),
    .I_135(n1_I_135),
    .I_136(n1_I_136),
    .I_137(n1_I_137),
    .I_138(n1_I_138),
    .I_139(n1_I_139),
    .I_140(n1_I_140),
    .I_141(n1_I_141),
    .I_142(n1_I_142),
    .I_143(n1_I_143),
    .I_144(n1_I_144),
    .I_145(n1_I_145),
    .I_146(n1_I_146),
    .I_147(n1_I_147),
    .I_148(n1_I_148),
    .I_149(n1_I_149),
    .I_150(n1_I_150),
    .I_151(n1_I_151),
    .I_152(n1_I_152),
    .I_153(n1_I_153),
    .I_154(n1_I_154),
    .I_155(n1_I_155),
    .I_156(n1_I_156),
    .I_157(n1_I_157),
    .I_158(n1_I_158),
    .I_159(n1_I_159),
    .I_160(n1_I_160),
    .I_161(n1_I_161),
    .I_162(n1_I_162),
    .I_163(n1_I_163),
    .I_164(n1_I_164),
    .I_165(n1_I_165),
    .I_166(n1_I_166),
    .I_167(n1_I_167),
    .I_168(n1_I_168),
    .I_169(n1_I_169),
    .I_170(n1_I_170),
    .I_171(n1_I_171),
    .I_172(n1_I_172),
    .I_173(n1_I_173),
    .I_174(n1_I_174),
    .I_175(n1_I_175),
    .I_176(n1_I_176),
    .I_177(n1_I_177),
    .I_178(n1_I_178),
    .I_179(n1_I_179),
    .I_180(n1_I_180),
    .I_181(n1_I_181),
    .I_182(n1_I_182),
    .I_183(n1_I_183),
    .I_184(n1_I_184),
    .I_185(n1_I_185),
    .I_186(n1_I_186),
    .I_187(n1_I_187),
    .I_188(n1_I_188),
    .I_189(n1_I_189),
    .I_190(n1_I_190),
    .I_191(n1_I_191),
    .I_192(n1_I_192),
    .I_193(n1_I_193),
    .I_194(n1_I_194),
    .I_195(n1_I_195),
    .I_196(n1_I_196),
    .I_197(n1_I_197),
    .I_198(n1_I_198),
    .I_199(n1_I_199),
    .O_0(n1_O_0),
    .O_1(n1_O_1),
    .O_2(n1_O_2),
    .O_3(n1_O_3),
    .O_4(n1_O_4),
    .O_5(n1_O_5),
    .O_6(n1_O_6),
    .O_7(n1_O_7),
    .O_8(n1_O_8),
    .O_9(n1_O_9),
    .O_10(n1_O_10),
    .O_11(n1_O_11),
    .O_12(n1_O_12),
    .O_13(n1_O_13),
    .O_14(n1_O_14),
    .O_15(n1_O_15),
    .O_16(n1_O_16),
    .O_17(n1_O_17),
    .O_18(n1_O_18),
    .O_19(n1_O_19),
    .O_20(n1_O_20),
    .O_21(n1_O_21),
    .O_22(n1_O_22),
    .O_23(n1_O_23),
    .O_24(n1_O_24),
    .O_25(n1_O_25),
    .O_26(n1_O_26),
    .O_27(n1_O_27),
    .O_28(n1_O_28),
    .O_29(n1_O_29),
    .O_30(n1_O_30),
    .O_31(n1_O_31),
    .O_32(n1_O_32),
    .O_33(n1_O_33),
    .O_34(n1_O_34),
    .O_35(n1_O_35),
    .O_36(n1_O_36),
    .O_37(n1_O_37),
    .O_38(n1_O_38),
    .O_39(n1_O_39),
    .O_40(n1_O_40),
    .O_41(n1_O_41),
    .O_42(n1_O_42),
    .O_43(n1_O_43),
    .O_44(n1_O_44),
    .O_45(n1_O_45),
    .O_46(n1_O_46),
    .O_47(n1_O_47),
    .O_48(n1_O_48),
    .O_49(n1_O_49),
    .O_50(n1_O_50),
    .O_51(n1_O_51),
    .O_52(n1_O_52),
    .O_53(n1_O_53),
    .O_54(n1_O_54),
    .O_55(n1_O_55),
    .O_56(n1_O_56),
    .O_57(n1_O_57),
    .O_58(n1_O_58),
    .O_59(n1_O_59),
    .O_60(n1_O_60),
    .O_61(n1_O_61),
    .O_62(n1_O_62),
    .O_63(n1_O_63),
    .O_64(n1_O_64),
    .O_65(n1_O_65),
    .O_66(n1_O_66),
    .O_67(n1_O_67),
    .O_68(n1_O_68),
    .O_69(n1_O_69),
    .O_70(n1_O_70),
    .O_71(n1_O_71),
    .O_72(n1_O_72),
    .O_73(n1_O_73),
    .O_74(n1_O_74),
    .O_75(n1_O_75),
    .O_76(n1_O_76),
    .O_77(n1_O_77),
    .O_78(n1_O_78),
    .O_79(n1_O_79),
    .O_80(n1_O_80),
    .O_81(n1_O_81),
    .O_82(n1_O_82),
    .O_83(n1_O_83),
    .O_84(n1_O_84),
    .O_85(n1_O_85),
    .O_86(n1_O_86),
    .O_87(n1_O_87),
    .O_88(n1_O_88),
    .O_89(n1_O_89),
    .O_90(n1_O_90),
    .O_91(n1_O_91),
    .O_92(n1_O_92),
    .O_93(n1_O_93),
    .O_94(n1_O_94),
    .O_95(n1_O_95),
    .O_96(n1_O_96),
    .O_97(n1_O_97),
    .O_98(n1_O_98),
    .O_99(n1_O_99),
    .O_100(n1_O_100),
    .O_101(n1_O_101),
    .O_102(n1_O_102),
    .O_103(n1_O_103),
    .O_104(n1_O_104),
    .O_105(n1_O_105),
    .O_106(n1_O_106),
    .O_107(n1_O_107),
    .O_108(n1_O_108),
    .O_109(n1_O_109),
    .O_110(n1_O_110),
    .O_111(n1_O_111),
    .O_112(n1_O_112),
    .O_113(n1_O_113),
    .O_114(n1_O_114),
    .O_115(n1_O_115),
    .O_116(n1_O_116),
    .O_117(n1_O_117),
    .O_118(n1_O_118),
    .O_119(n1_O_119),
    .O_120(n1_O_120),
    .O_121(n1_O_121),
    .O_122(n1_O_122),
    .O_123(n1_O_123),
    .O_124(n1_O_124),
    .O_125(n1_O_125),
    .O_126(n1_O_126),
    .O_127(n1_O_127),
    .O_128(n1_O_128),
    .O_129(n1_O_129),
    .O_130(n1_O_130),
    .O_131(n1_O_131),
    .O_132(n1_O_132),
    .O_133(n1_O_133),
    .O_134(n1_O_134),
    .O_135(n1_O_135),
    .O_136(n1_O_136),
    .O_137(n1_O_137),
    .O_138(n1_O_138),
    .O_139(n1_O_139),
    .O_140(n1_O_140),
    .O_141(n1_O_141),
    .O_142(n1_O_142),
    .O_143(n1_O_143),
    .O_144(n1_O_144),
    .O_145(n1_O_145),
    .O_146(n1_O_146),
    .O_147(n1_O_147),
    .O_148(n1_O_148),
    .O_149(n1_O_149),
    .O_150(n1_O_150),
    .O_151(n1_O_151),
    .O_152(n1_O_152),
    .O_153(n1_O_153),
    .O_154(n1_O_154),
    .O_155(n1_O_155),
    .O_156(n1_O_156),
    .O_157(n1_O_157),
    .O_158(n1_O_158),
    .O_159(n1_O_159),
    .O_160(n1_O_160),
    .O_161(n1_O_161),
    .O_162(n1_O_162),
    .O_163(n1_O_163),
    .O_164(n1_O_164),
    .O_165(n1_O_165),
    .O_166(n1_O_166),
    .O_167(n1_O_167),
    .O_168(n1_O_168),
    .O_169(n1_O_169),
    .O_170(n1_O_170),
    .O_171(n1_O_171),
    .O_172(n1_O_172),
    .O_173(n1_O_173),
    .O_174(n1_O_174),
    .O_175(n1_O_175),
    .O_176(n1_O_176),
    .O_177(n1_O_177),
    .O_178(n1_O_178),
    .O_179(n1_O_179),
    .O_180(n1_O_180),
    .O_181(n1_O_181),
    .O_182(n1_O_182),
    .O_183(n1_O_183),
    .O_184(n1_O_184),
    .O_185(n1_O_185),
    .O_186(n1_O_186),
    .O_187(n1_O_187),
    .O_188(n1_O_188),
    .O_189(n1_O_189),
    .O_190(n1_O_190),
    .O_191(n1_O_191),
    .O_192(n1_O_192),
    .O_193(n1_O_193),
    .O_194(n1_O_194),
    .O_195(n1_O_195),
    .O_196(n1_O_196),
    .O_197(n1_O_197),
    .O_198(n1_O_198),
    .O_199(n1_O_199)
  );
  MapS n7 ( // @[Top.scala 35:20]
    .clock(n7_clock),
    .reset(n7_reset),
    .valid_up(n7_valid_up),
    .valid_down(n7_valid_down),
    .I_0(n7_I_0),
    .I_1(n7_I_1),
    .I_2(n7_I_2),
    .I_3(n7_I_3),
    .I_4(n7_I_4),
    .I_5(n7_I_5),
    .I_6(n7_I_6),
    .I_7(n7_I_7),
    .I_8(n7_I_8),
    .I_9(n7_I_9),
    .I_10(n7_I_10),
    .I_11(n7_I_11),
    .I_12(n7_I_12),
    .I_13(n7_I_13),
    .I_14(n7_I_14),
    .I_15(n7_I_15),
    .I_16(n7_I_16),
    .I_17(n7_I_17),
    .I_18(n7_I_18),
    .I_19(n7_I_19),
    .I_20(n7_I_20),
    .I_21(n7_I_21),
    .I_22(n7_I_22),
    .I_23(n7_I_23),
    .I_24(n7_I_24),
    .I_25(n7_I_25),
    .I_26(n7_I_26),
    .I_27(n7_I_27),
    .I_28(n7_I_28),
    .I_29(n7_I_29),
    .I_30(n7_I_30),
    .I_31(n7_I_31),
    .I_32(n7_I_32),
    .I_33(n7_I_33),
    .I_34(n7_I_34),
    .I_35(n7_I_35),
    .I_36(n7_I_36),
    .I_37(n7_I_37),
    .I_38(n7_I_38),
    .I_39(n7_I_39),
    .I_40(n7_I_40),
    .I_41(n7_I_41),
    .I_42(n7_I_42),
    .I_43(n7_I_43),
    .I_44(n7_I_44),
    .I_45(n7_I_45),
    .I_46(n7_I_46),
    .I_47(n7_I_47),
    .I_48(n7_I_48),
    .I_49(n7_I_49),
    .I_50(n7_I_50),
    .I_51(n7_I_51),
    .I_52(n7_I_52),
    .I_53(n7_I_53),
    .I_54(n7_I_54),
    .I_55(n7_I_55),
    .I_56(n7_I_56),
    .I_57(n7_I_57),
    .I_58(n7_I_58),
    .I_59(n7_I_59),
    .I_60(n7_I_60),
    .I_61(n7_I_61),
    .I_62(n7_I_62),
    .I_63(n7_I_63),
    .I_64(n7_I_64),
    .I_65(n7_I_65),
    .I_66(n7_I_66),
    .I_67(n7_I_67),
    .I_68(n7_I_68),
    .I_69(n7_I_69),
    .I_70(n7_I_70),
    .I_71(n7_I_71),
    .I_72(n7_I_72),
    .I_73(n7_I_73),
    .I_74(n7_I_74),
    .I_75(n7_I_75),
    .I_76(n7_I_76),
    .I_77(n7_I_77),
    .I_78(n7_I_78),
    .I_79(n7_I_79),
    .I_80(n7_I_80),
    .I_81(n7_I_81),
    .I_82(n7_I_82),
    .I_83(n7_I_83),
    .I_84(n7_I_84),
    .I_85(n7_I_85),
    .I_86(n7_I_86),
    .I_87(n7_I_87),
    .I_88(n7_I_88),
    .I_89(n7_I_89),
    .I_90(n7_I_90),
    .I_91(n7_I_91),
    .I_92(n7_I_92),
    .I_93(n7_I_93),
    .I_94(n7_I_94),
    .I_95(n7_I_95),
    .I_96(n7_I_96),
    .I_97(n7_I_97),
    .I_98(n7_I_98),
    .I_99(n7_I_99),
    .I_100(n7_I_100),
    .I_101(n7_I_101),
    .I_102(n7_I_102),
    .I_103(n7_I_103),
    .I_104(n7_I_104),
    .I_105(n7_I_105),
    .I_106(n7_I_106),
    .I_107(n7_I_107),
    .I_108(n7_I_108),
    .I_109(n7_I_109),
    .I_110(n7_I_110),
    .I_111(n7_I_111),
    .I_112(n7_I_112),
    .I_113(n7_I_113),
    .I_114(n7_I_114),
    .I_115(n7_I_115),
    .I_116(n7_I_116),
    .I_117(n7_I_117),
    .I_118(n7_I_118),
    .I_119(n7_I_119),
    .I_120(n7_I_120),
    .I_121(n7_I_121),
    .I_122(n7_I_122),
    .I_123(n7_I_123),
    .I_124(n7_I_124),
    .I_125(n7_I_125),
    .I_126(n7_I_126),
    .I_127(n7_I_127),
    .I_128(n7_I_128),
    .I_129(n7_I_129),
    .I_130(n7_I_130),
    .I_131(n7_I_131),
    .I_132(n7_I_132),
    .I_133(n7_I_133),
    .I_134(n7_I_134),
    .I_135(n7_I_135),
    .I_136(n7_I_136),
    .I_137(n7_I_137),
    .I_138(n7_I_138),
    .I_139(n7_I_139),
    .I_140(n7_I_140),
    .I_141(n7_I_141),
    .I_142(n7_I_142),
    .I_143(n7_I_143),
    .I_144(n7_I_144),
    .I_145(n7_I_145),
    .I_146(n7_I_146),
    .I_147(n7_I_147),
    .I_148(n7_I_148),
    .I_149(n7_I_149),
    .I_150(n7_I_150),
    .I_151(n7_I_151),
    .I_152(n7_I_152),
    .I_153(n7_I_153),
    .I_154(n7_I_154),
    .I_155(n7_I_155),
    .I_156(n7_I_156),
    .I_157(n7_I_157),
    .I_158(n7_I_158),
    .I_159(n7_I_159),
    .I_160(n7_I_160),
    .I_161(n7_I_161),
    .I_162(n7_I_162),
    .I_163(n7_I_163),
    .I_164(n7_I_164),
    .I_165(n7_I_165),
    .I_166(n7_I_166),
    .I_167(n7_I_167),
    .I_168(n7_I_168),
    .I_169(n7_I_169),
    .I_170(n7_I_170),
    .I_171(n7_I_171),
    .I_172(n7_I_172),
    .I_173(n7_I_173),
    .I_174(n7_I_174),
    .I_175(n7_I_175),
    .I_176(n7_I_176),
    .I_177(n7_I_177),
    .I_178(n7_I_178),
    .I_179(n7_I_179),
    .I_180(n7_I_180),
    .I_181(n7_I_181),
    .I_182(n7_I_182),
    .I_183(n7_I_183),
    .I_184(n7_I_184),
    .I_185(n7_I_185),
    .I_186(n7_I_186),
    .I_187(n7_I_187),
    .I_188(n7_I_188),
    .I_189(n7_I_189),
    .I_190(n7_I_190),
    .I_191(n7_I_191),
    .I_192(n7_I_192),
    .I_193(n7_I_193),
    .I_194(n7_I_194),
    .I_195(n7_I_195),
    .I_196(n7_I_196),
    .I_197(n7_I_197),
    .I_198(n7_I_198),
    .I_199(n7_I_199),
    .O_0(n7_O_0),
    .O_1(n7_O_1),
    .O_2(n7_O_2),
    .O_3(n7_O_3),
    .O_4(n7_O_4),
    .O_5(n7_O_5),
    .O_6(n7_O_6),
    .O_7(n7_O_7),
    .O_8(n7_O_8),
    .O_9(n7_O_9),
    .O_10(n7_O_10),
    .O_11(n7_O_11),
    .O_12(n7_O_12),
    .O_13(n7_O_13),
    .O_14(n7_O_14),
    .O_15(n7_O_15),
    .O_16(n7_O_16),
    .O_17(n7_O_17),
    .O_18(n7_O_18),
    .O_19(n7_O_19),
    .O_20(n7_O_20),
    .O_21(n7_O_21),
    .O_22(n7_O_22),
    .O_23(n7_O_23),
    .O_24(n7_O_24),
    .O_25(n7_O_25),
    .O_26(n7_O_26),
    .O_27(n7_O_27),
    .O_28(n7_O_28),
    .O_29(n7_O_29),
    .O_30(n7_O_30),
    .O_31(n7_O_31),
    .O_32(n7_O_32),
    .O_33(n7_O_33),
    .O_34(n7_O_34),
    .O_35(n7_O_35),
    .O_36(n7_O_36),
    .O_37(n7_O_37),
    .O_38(n7_O_38),
    .O_39(n7_O_39),
    .O_40(n7_O_40),
    .O_41(n7_O_41),
    .O_42(n7_O_42),
    .O_43(n7_O_43),
    .O_44(n7_O_44),
    .O_45(n7_O_45),
    .O_46(n7_O_46),
    .O_47(n7_O_47),
    .O_48(n7_O_48),
    .O_49(n7_O_49),
    .O_50(n7_O_50),
    .O_51(n7_O_51),
    .O_52(n7_O_52),
    .O_53(n7_O_53),
    .O_54(n7_O_54),
    .O_55(n7_O_55),
    .O_56(n7_O_56),
    .O_57(n7_O_57),
    .O_58(n7_O_58),
    .O_59(n7_O_59),
    .O_60(n7_O_60),
    .O_61(n7_O_61),
    .O_62(n7_O_62),
    .O_63(n7_O_63),
    .O_64(n7_O_64),
    .O_65(n7_O_65),
    .O_66(n7_O_66),
    .O_67(n7_O_67),
    .O_68(n7_O_68),
    .O_69(n7_O_69),
    .O_70(n7_O_70),
    .O_71(n7_O_71),
    .O_72(n7_O_72),
    .O_73(n7_O_73),
    .O_74(n7_O_74),
    .O_75(n7_O_75),
    .O_76(n7_O_76),
    .O_77(n7_O_77),
    .O_78(n7_O_78),
    .O_79(n7_O_79),
    .O_80(n7_O_80),
    .O_81(n7_O_81),
    .O_82(n7_O_82),
    .O_83(n7_O_83),
    .O_84(n7_O_84),
    .O_85(n7_O_85),
    .O_86(n7_O_86),
    .O_87(n7_O_87),
    .O_88(n7_O_88),
    .O_89(n7_O_89),
    .O_90(n7_O_90),
    .O_91(n7_O_91),
    .O_92(n7_O_92),
    .O_93(n7_O_93),
    .O_94(n7_O_94),
    .O_95(n7_O_95),
    .O_96(n7_O_96),
    .O_97(n7_O_97),
    .O_98(n7_O_98),
    .O_99(n7_O_99),
    .O_100(n7_O_100),
    .O_101(n7_O_101),
    .O_102(n7_O_102),
    .O_103(n7_O_103),
    .O_104(n7_O_104),
    .O_105(n7_O_105),
    .O_106(n7_O_106),
    .O_107(n7_O_107),
    .O_108(n7_O_108),
    .O_109(n7_O_109),
    .O_110(n7_O_110),
    .O_111(n7_O_111),
    .O_112(n7_O_112),
    .O_113(n7_O_113),
    .O_114(n7_O_114),
    .O_115(n7_O_115),
    .O_116(n7_O_116),
    .O_117(n7_O_117),
    .O_118(n7_O_118),
    .O_119(n7_O_119),
    .O_120(n7_O_120),
    .O_121(n7_O_121),
    .O_122(n7_O_122),
    .O_123(n7_O_123),
    .O_124(n7_O_124),
    .O_125(n7_O_125),
    .O_126(n7_O_126),
    .O_127(n7_O_127),
    .O_128(n7_O_128),
    .O_129(n7_O_129),
    .O_130(n7_O_130),
    .O_131(n7_O_131),
    .O_132(n7_O_132),
    .O_133(n7_O_133),
    .O_134(n7_O_134),
    .O_135(n7_O_135),
    .O_136(n7_O_136),
    .O_137(n7_O_137),
    .O_138(n7_O_138),
    .O_139(n7_O_139),
    .O_140(n7_O_140),
    .O_141(n7_O_141),
    .O_142(n7_O_142),
    .O_143(n7_O_143),
    .O_144(n7_O_144),
    .O_145(n7_O_145),
    .O_146(n7_O_146),
    .O_147(n7_O_147),
    .O_148(n7_O_148),
    .O_149(n7_O_149),
    .O_150(n7_O_150),
    .O_151(n7_O_151),
    .O_152(n7_O_152),
    .O_153(n7_O_153),
    .O_154(n7_O_154),
    .O_155(n7_O_155),
    .O_156(n7_O_156),
    .O_157(n7_O_157),
    .O_158(n7_O_158),
    .O_159(n7_O_159),
    .O_160(n7_O_160),
    .O_161(n7_O_161),
    .O_162(n7_O_162),
    .O_163(n7_O_163),
    .O_164(n7_O_164),
    .O_165(n7_O_165),
    .O_166(n7_O_166),
    .O_167(n7_O_167),
    .O_168(n7_O_168),
    .O_169(n7_O_169),
    .O_170(n7_O_170),
    .O_171(n7_O_171),
    .O_172(n7_O_172),
    .O_173(n7_O_173),
    .O_174(n7_O_174),
    .O_175(n7_O_175),
    .O_176(n7_O_176),
    .O_177(n7_O_177),
    .O_178(n7_O_178),
    .O_179(n7_O_179),
    .O_180(n7_O_180),
    .O_181(n7_O_181),
    .O_182(n7_O_182),
    .O_183(n7_O_183),
    .O_184(n7_O_184),
    .O_185(n7_O_185),
    .O_186(n7_O_186),
    .O_187(n7_O_187),
    .O_188(n7_O_188),
    .O_189(n7_O_189),
    .O_190(n7_O_190),
    .O_191(n7_O_191),
    .O_192(n7_O_192),
    .O_193(n7_O_193),
    .O_194(n7_O_194),
    .O_195(n7_O_195),
    .O_196(n7_O_196),
    .O_197(n7_O_197),
    .O_198(n7_O_198),
    .O_199(n7_O_199)
  );
  FIFO n8 ( // @[Top.scala 38:20]
    .clock(n8_clock),
    .reset(n8_reset),
    .valid_up(n8_valid_up),
    .valid_down(n8_valid_down),
    .I_0(n8_I_0),
    .I_1(n8_I_1),
    .I_2(n8_I_2),
    .I_3(n8_I_3),
    .I_4(n8_I_4),
    .I_5(n8_I_5),
    .I_6(n8_I_6),
    .I_7(n8_I_7),
    .I_8(n8_I_8),
    .I_9(n8_I_9),
    .I_10(n8_I_10),
    .I_11(n8_I_11),
    .I_12(n8_I_12),
    .I_13(n8_I_13),
    .I_14(n8_I_14),
    .I_15(n8_I_15),
    .I_16(n8_I_16),
    .I_17(n8_I_17),
    .I_18(n8_I_18),
    .I_19(n8_I_19),
    .I_20(n8_I_20),
    .I_21(n8_I_21),
    .I_22(n8_I_22),
    .I_23(n8_I_23),
    .I_24(n8_I_24),
    .I_25(n8_I_25),
    .I_26(n8_I_26),
    .I_27(n8_I_27),
    .I_28(n8_I_28),
    .I_29(n8_I_29),
    .I_30(n8_I_30),
    .I_31(n8_I_31),
    .I_32(n8_I_32),
    .I_33(n8_I_33),
    .I_34(n8_I_34),
    .I_35(n8_I_35),
    .I_36(n8_I_36),
    .I_37(n8_I_37),
    .I_38(n8_I_38),
    .I_39(n8_I_39),
    .I_40(n8_I_40),
    .I_41(n8_I_41),
    .I_42(n8_I_42),
    .I_43(n8_I_43),
    .I_44(n8_I_44),
    .I_45(n8_I_45),
    .I_46(n8_I_46),
    .I_47(n8_I_47),
    .I_48(n8_I_48),
    .I_49(n8_I_49),
    .I_50(n8_I_50),
    .I_51(n8_I_51),
    .I_52(n8_I_52),
    .I_53(n8_I_53),
    .I_54(n8_I_54),
    .I_55(n8_I_55),
    .I_56(n8_I_56),
    .I_57(n8_I_57),
    .I_58(n8_I_58),
    .I_59(n8_I_59),
    .I_60(n8_I_60),
    .I_61(n8_I_61),
    .I_62(n8_I_62),
    .I_63(n8_I_63),
    .I_64(n8_I_64),
    .I_65(n8_I_65),
    .I_66(n8_I_66),
    .I_67(n8_I_67),
    .I_68(n8_I_68),
    .I_69(n8_I_69),
    .I_70(n8_I_70),
    .I_71(n8_I_71),
    .I_72(n8_I_72),
    .I_73(n8_I_73),
    .I_74(n8_I_74),
    .I_75(n8_I_75),
    .I_76(n8_I_76),
    .I_77(n8_I_77),
    .I_78(n8_I_78),
    .I_79(n8_I_79),
    .I_80(n8_I_80),
    .I_81(n8_I_81),
    .I_82(n8_I_82),
    .I_83(n8_I_83),
    .I_84(n8_I_84),
    .I_85(n8_I_85),
    .I_86(n8_I_86),
    .I_87(n8_I_87),
    .I_88(n8_I_88),
    .I_89(n8_I_89),
    .I_90(n8_I_90),
    .I_91(n8_I_91),
    .I_92(n8_I_92),
    .I_93(n8_I_93),
    .I_94(n8_I_94),
    .I_95(n8_I_95),
    .I_96(n8_I_96),
    .I_97(n8_I_97),
    .I_98(n8_I_98),
    .I_99(n8_I_99),
    .I_100(n8_I_100),
    .I_101(n8_I_101),
    .I_102(n8_I_102),
    .I_103(n8_I_103),
    .I_104(n8_I_104),
    .I_105(n8_I_105),
    .I_106(n8_I_106),
    .I_107(n8_I_107),
    .I_108(n8_I_108),
    .I_109(n8_I_109),
    .I_110(n8_I_110),
    .I_111(n8_I_111),
    .I_112(n8_I_112),
    .I_113(n8_I_113),
    .I_114(n8_I_114),
    .I_115(n8_I_115),
    .I_116(n8_I_116),
    .I_117(n8_I_117),
    .I_118(n8_I_118),
    .I_119(n8_I_119),
    .I_120(n8_I_120),
    .I_121(n8_I_121),
    .I_122(n8_I_122),
    .I_123(n8_I_123),
    .I_124(n8_I_124),
    .I_125(n8_I_125),
    .I_126(n8_I_126),
    .I_127(n8_I_127),
    .I_128(n8_I_128),
    .I_129(n8_I_129),
    .I_130(n8_I_130),
    .I_131(n8_I_131),
    .I_132(n8_I_132),
    .I_133(n8_I_133),
    .I_134(n8_I_134),
    .I_135(n8_I_135),
    .I_136(n8_I_136),
    .I_137(n8_I_137),
    .I_138(n8_I_138),
    .I_139(n8_I_139),
    .I_140(n8_I_140),
    .I_141(n8_I_141),
    .I_142(n8_I_142),
    .I_143(n8_I_143),
    .I_144(n8_I_144),
    .I_145(n8_I_145),
    .I_146(n8_I_146),
    .I_147(n8_I_147),
    .I_148(n8_I_148),
    .I_149(n8_I_149),
    .I_150(n8_I_150),
    .I_151(n8_I_151),
    .I_152(n8_I_152),
    .I_153(n8_I_153),
    .I_154(n8_I_154),
    .I_155(n8_I_155),
    .I_156(n8_I_156),
    .I_157(n8_I_157),
    .I_158(n8_I_158),
    .I_159(n8_I_159),
    .I_160(n8_I_160),
    .I_161(n8_I_161),
    .I_162(n8_I_162),
    .I_163(n8_I_163),
    .I_164(n8_I_164),
    .I_165(n8_I_165),
    .I_166(n8_I_166),
    .I_167(n8_I_167),
    .I_168(n8_I_168),
    .I_169(n8_I_169),
    .I_170(n8_I_170),
    .I_171(n8_I_171),
    .I_172(n8_I_172),
    .I_173(n8_I_173),
    .I_174(n8_I_174),
    .I_175(n8_I_175),
    .I_176(n8_I_176),
    .I_177(n8_I_177),
    .I_178(n8_I_178),
    .I_179(n8_I_179),
    .I_180(n8_I_180),
    .I_181(n8_I_181),
    .I_182(n8_I_182),
    .I_183(n8_I_183),
    .I_184(n8_I_184),
    .I_185(n8_I_185),
    .I_186(n8_I_186),
    .I_187(n8_I_187),
    .I_188(n8_I_188),
    .I_189(n8_I_189),
    .I_190(n8_I_190),
    .I_191(n8_I_191),
    .I_192(n8_I_192),
    .I_193(n8_I_193),
    .I_194(n8_I_194),
    .I_195(n8_I_195),
    .I_196(n8_I_196),
    .I_197(n8_I_197),
    .I_198(n8_I_198),
    .I_199(n8_I_199),
    .O_0(n8_O_0),
    .O_1(n8_O_1),
    .O_2(n8_O_2),
    .O_3(n8_O_3),
    .O_4(n8_O_4),
    .O_5(n8_O_5),
    .O_6(n8_O_6),
    .O_7(n8_O_7),
    .O_8(n8_O_8),
    .O_9(n8_O_9),
    .O_10(n8_O_10),
    .O_11(n8_O_11),
    .O_12(n8_O_12),
    .O_13(n8_O_13),
    .O_14(n8_O_14),
    .O_15(n8_O_15),
    .O_16(n8_O_16),
    .O_17(n8_O_17),
    .O_18(n8_O_18),
    .O_19(n8_O_19),
    .O_20(n8_O_20),
    .O_21(n8_O_21),
    .O_22(n8_O_22),
    .O_23(n8_O_23),
    .O_24(n8_O_24),
    .O_25(n8_O_25),
    .O_26(n8_O_26),
    .O_27(n8_O_27),
    .O_28(n8_O_28),
    .O_29(n8_O_29),
    .O_30(n8_O_30),
    .O_31(n8_O_31),
    .O_32(n8_O_32),
    .O_33(n8_O_33),
    .O_34(n8_O_34),
    .O_35(n8_O_35),
    .O_36(n8_O_36),
    .O_37(n8_O_37),
    .O_38(n8_O_38),
    .O_39(n8_O_39),
    .O_40(n8_O_40),
    .O_41(n8_O_41),
    .O_42(n8_O_42),
    .O_43(n8_O_43),
    .O_44(n8_O_44),
    .O_45(n8_O_45),
    .O_46(n8_O_46),
    .O_47(n8_O_47),
    .O_48(n8_O_48),
    .O_49(n8_O_49),
    .O_50(n8_O_50),
    .O_51(n8_O_51),
    .O_52(n8_O_52),
    .O_53(n8_O_53),
    .O_54(n8_O_54),
    .O_55(n8_O_55),
    .O_56(n8_O_56),
    .O_57(n8_O_57),
    .O_58(n8_O_58),
    .O_59(n8_O_59),
    .O_60(n8_O_60),
    .O_61(n8_O_61),
    .O_62(n8_O_62),
    .O_63(n8_O_63),
    .O_64(n8_O_64),
    .O_65(n8_O_65),
    .O_66(n8_O_66),
    .O_67(n8_O_67),
    .O_68(n8_O_68),
    .O_69(n8_O_69),
    .O_70(n8_O_70),
    .O_71(n8_O_71),
    .O_72(n8_O_72),
    .O_73(n8_O_73),
    .O_74(n8_O_74),
    .O_75(n8_O_75),
    .O_76(n8_O_76),
    .O_77(n8_O_77),
    .O_78(n8_O_78),
    .O_79(n8_O_79),
    .O_80(n8_O_80),
    .O_81(n8_O_81),
    .O_82(n8_O_82),
    .O_83(n8_O_83),
    .O_84(n8_O_84),
    .O_85(n8_O_85),
    .O_86(n8_O_86),
    .O_87(n8_O_87),
    .O_88(n8_O_88),
    .O_89(n8_O_89),
    .O_90(n8_O_90),
    .O_91(n8_O_91),
    .O_92(n8_O_92),
    .O_93(n8_O_93),
    .O_94(n8_O_94),
    .O_95(n8_O_95),
    .O_96(n8_O_96),
    .O_97(n8_O_97),
    .O_98(n8_O_98),
    .O_99(n8_O_99),
    .O_100(n8_O_100),
    .O_101(n8_O_101),
    .O_102(n8_O_102),
    .O_103(n8_O_103),
    .O_104(n8_O_104),
    .O_105(n8_O_105),
    .O_106(n8_O_106),
    .O_107(n8_O_107),
    .O_108(n8_O_108),
    .O_109(n8_O_109),
    .O_110(n8_O_110),
    .O_111(n8_O_111),
    .O_112(n8_O_112),
    .O_113(n8_O_113),
    .O_114(n8_O_114),
    .O_115(n8_O_115),
    .O_116(n8_O_116),
    .O_117(n8_O_117),
    .O_118(n8_O_118),
    .O_119(n8_O_119),
    .O_120(n8_O_120),
    .O_121(n8_O_121),
    .O_122(n8_O_122),
    .O_123(n8_O_123),
    .O_124(n8_O_124),
    .O_125(n8_O_125),
    .O_126(n8_O_126),
    .O_127(n8_O_127),
    .O_128(n8_O_128),
    .O_129(n8_O_129),
    .O_130(n8_O_130),
    .O_131(n8_O_131),
    .O_132(n8_O_132),
    .O_133(n8_O_133),
    .O_134(n8_O_134),
    .O_135(n8_O_135),
    .O_136(n8_O_136),
    .O_137(n8_O_137),
    .O_138(n8_O_138),
    .O_139(n8_O_139),
    .O_140(n8_O_140),
    .O_141(n8_O_141),
    .O_142(n8_O_142),
    .O_143(n8_O_143),
    .O_144(n8_O_144),
    .O_145(n8_O_145),
    .O_146(n8_O_146),
    .O_147(n8_O_147),
    .O_148(n8_O_148),
    .O_149(n8_O_149),
    .O_150(n8_O_150),
    .O_151(n8_O_151),
    .O_152(n8_O_152),
    .O_153(n8_O_153),
    .O_154(n8_O_154),
    .O_155(n8_O_155),
    .O_156(n8_O_156),
    .O_157(n8_O_157),
    .O_158(n8_O_158),
    .O_159(n8_O_159),
    .O_160(n8_O_160),
    .O_161(n8_O_161),
    .O_162(n8_O_162),
    .O_163(n8_O_163),
    .O_164(n8_O_164),
    .O_165(n8_O_165),
    .O_166(n8_O_166),
    .O_167(n8_O_167),
    .O_168(n8_O_168),
    .O_169(n8_O_169),
    .O_170(n8_O_170),
    .O_171(n8_O_171),
    .O_172(n8_O_172),
    .O_173(n8_O_173),
    .O_174(n8_O_174),
    .O_175(n8_O_175),
    .O_176(n8_O_176),
    .O_177(n8_O_177),
    .O_178(n8_O_178),
    .O_179(n8_O_179),
    .O_180(n8_O_180),
    .O_181(n8_O_181),
    .O_182(n8_O_182),
    .O_183(n8_O_183),
    .O_184(n8_O_184),
    .O_185(n8_O_185),
    .O_186(n8_O_186),
    .O_187(n8_O_187),
    .O_188(n8_O_188),
    .O_189(n8_O_189),
    .O_190(n8_O_190),
    .O_191(n8_O_191),
    .O_192(n8_O_192),
    .O_193(n8_O_193),
    .O_194(n8_O_194),
    .O_195(n8_O_195),
    .O_196(n8_O_196),
    .O_197(n8_O_197),
    .O_198(n8_O_198),
    .O_199(n8_O_199)
  );
  FIFO n9 ( // @[Top.scala 41:20]
    .clock(n9_clock),
    .reset(n9_reset),
    .valid_up(n9_valid_up),
    .valid_down(n9_valid_down),
    .I_0(n9_I_0),
    .I_1(n9_I_1),
    .I_2(n9_I_2),
    .I_3(n9_I_3),
    .I_4(n9_I_4),
    .I_5(n9_I_5),
    .I_6(n9_I_6),
    .I_7(n9_I_7),
    .I_8(n9_I_8),
    .I_9(n9_I_9),
    .I_10(n9_I_10),
    .I_11(n9_I_11),
    .I_12(n9_I_12),
    .I_13(n9_I_13),
    .I_14(n9_I_14),
    .I_15(n9_I_15),
    .I_16(n9_I_16),
    .I_17(n9_I_17),
    .I_18(n9_I_18),
    .I_19(n9_I_19),
    .I_20(n9_I_20),
    .I_21(n9_I_21),
    .I_22(n9_I_22),
    .I_23(n9_I_23),
    .I_24(n9_I_24),
    .I_25(n9_I_25),
    .I_26(n9_I_26),
    .I_27(n9_I_27),
    .I_28(n9_I_28),
    .I_29(n9_I_29),
    .I_30(n9_I_30),
    .I_31(n9_I_31),
    .I_32(n9_I_32),
    .I_33(n9_I_33),
    .I_34(n9_I_34),
    .I_35(n9_I_35),
    .I_36(n9_I_36),
    .I_37(n9_I_37),
    .I_38(n9_I_38),
    .I_39(n9_I_39),
    .I_40(n9_I_40),
    .I_41(n9_I_41),
    .I_42(n9_I_42),
    .I_43(n9_I_43),
    .I_44(n9_I_44),
    .I_45(n9_I_45),
    .I_46(n9_I_46),
    .I_47(n9_I_47),
    .I_48(n9_I_48),
    .I_49(n9_I_49),
    .I_50(n9_I_50),
    .I_51(n9_I_51),
    .I_52(n9_I_52),
    .I_53(n9_I_53),
    .I_54(n9_I_54),
    .I_55(n9_I_55),
    .I_56(n9_I_56),
    .I_57(n9_I_57),
    .I_58(n9_I_58),
    .I_59(n9_I_59),
    .I_60(n9_I_60),
    .I_61(n9_I_61),
    .I_62(n9_I_62),
    .I_63(n9_I_63),
    .I_64(n9_I_64),
    .I_65(n9_I_65),
    .I_66(n9_I_66),
    .I_67(n9_I_67),
    .I_68(n9_I_68),
    .I_69(n9_I_69),
    .I_70(n9_I_70),
    .I_71(n9_I_71),
    .I_72(n9_I_72),
    .I_73(n9_I_73),
    .I_74(n9_I_74),
    .I_75(n9_I_75),
    .I_76(n9_I_76),
    .I_77(n9_I_77),
    .I_78(n9_I_78),
    .I_79(n9_I_79),
    .I_80(n9_I_80),
    .I_81(n9_I_81),
    .I_82(n9_I_82),
    .I_83(n9_I_83),
    .I_84(n9_I_84),
    .I_85(n9_I_85),
    .I_86(n9_I_86),
    .I_87(n9_I_87),
    .I_88(n9_I_88),
    .I_89(n9_I_89),
    .I_90(n9_I_90),
    .I_91(n9_I_91),
    .I_92(n9_I_92),
    .I_93(n9_I_93),
    .I_94(n9_I_94),
    .I_95(n9_I_95),
    .I_96(n9_I_96),
    .I_97(n9_I_97),
    .I_98(n9_I_98),
    .I_99(n9_I_99),
    .I_100(n9_I_100),
    .I_101(n9_I_101),
    .I_102(n9_I_102),
    .I_103(n9_I_103),
    .I_104(n9_I_104),
    .I_105(n9_I_105),
    .I_106(n9_I_106),
    .I_107(n9_I_107),
    .I_108(n9_I_108),
    .I_109(n9_I_109),
    .I_110(n9_I_110),
    .I_111(n9_I_111),
    .I_112(n9_I_112),
    .I_113(n9_I_113),
    .I_114(n9_I_114),
    .I_115(n9_I_115),
    .I_116(n9_I_116),
    .I_117(n9_I_117),
    .I_118(n9_I_118),
    .I_119(n9_I_119),
    .I_120(n9_I_120),
    .I_121(n9_I_121),
    .I_122(n9_I_122),
    .I_123(n9_I_123),
    .I_124(n9_I_124),
    .I_125(n9_I_125),
    .I_126(n9_I_126),
    .I_127(n9_I_127),
    .I_128(n9_I_128),
    .I_129(n9_I_129),
    .I_130(n9_I_130),
    .I_131(n9_I_131),
    .I_132(n9_I_132),
    .I_133(n9_I_133),
    .I_134(n9_I_134),
    .I_135(n9_I_135),
    .I_136(n9_I_136),
    .I_137(n9_I_137),
    .I_138(n9_I_138),
    .I_139(n9_I_139),
    .I_140(n9_I_140),
    .I_141(n9_I_141),
    .I_142(n9_I_142),
    .I_143(n9_I_143),
    .I_144(n9_I_144),
    .I_145(n9_I_145),
    .I_146(n9_I_146),
    .I_147(n9_I_147),
    .I_148(n9_I_148),
    .I_149(n9_I_149),
    .I_150(n9_I_150),
    .I_151(n9_I_151),
    .I_152(n9_I_152),
    .I_153(n9_I_153),
    .I_154(n9_I_154),
    .I_155(n9_I_155),
    .I_156(n9_I_156),
    .I_157(n9_I_157),
    .I_158(n9_I_158),
    .I_159(n9_I_159),
    .I_160(n9_I_160),
    .I_161(n9_I_161),
    .I_162(n9_I_162),
    .I_163(n9_I_163),
    .I_164(n9_I_164),
    .I_165(n9_I_165),
    .I_166(n9_I_166),
    .I_167(n9_I_167),
    .I_168(n9_I_168),
    .I_169(n9_I_169),
    .I_170(n9_I_170),
    .I_171(n9_I_171),
    .I_172(n9_I_172),
    .I_173(n9_I_173),
    .I_174(n9_I_174),
    .I_175(n9_I_175),
    .I_176(n9_I_176),
    .I_177(n9_I_177),
    .I_178(n9_I_178),
    .I_179(n9_I_179),
    .I_180(n9_I_180),
    .I_181(n9_I_181),
    .I_182(n9_I_182),
    .I_183(n9_I_183),
    .I_184(n9_I_184),
    .I_185(n9_I_185),
    .I_186(n9_I_186),
    .I_187(n9_I_187),
    .I_188(n9_I_188),
    .I_189(n9_I_189),
    .I_190(n9_I_190),
    .I_191(n9_I_191),
    .I_192(n9_I_192),
    .I_193(n9_I_193),
    .I_194(n9_I_194),
    .I_195(n9_I_195),
    .I_196(n9_I_196),
    .I_197(n9_I_197),
    .I_198(n9_I_198),
    .I_199(n9_I_199),
    .O_0(n9_O_0),
    .O_1(n9_O_1),
    .O_2(n9_O_2),
    .O_3(n9_O_3),
    .O_4(n9_O_4),
    .O_5(n9_O_5),
    .O_6(n9_O_6),
    .O_7(n9_O_7),
    .O_8(n9_O_8),
    .O_9(n9_O_9),
    .O_10(n9_O_10),
    .O_11(n9_O_11),
    .O_12(n9_O_12),
    .O_13(n9_O_13),
    .O_14(n9_O_14),
    .O_15(n9_O_15),
    .O_16(n9_O_16),
    .O_17(n9_O_17),
    .O_18(n9_O_18),
    .O_19(n9_O_19),
    .O_20(n9_O_20),
    .O_21(n9_O_21),
    .O_22(n9_O_22),
    .O_23(n9_O_23),
    .O_24(n9_O_24),
    .O_25(n9_O_25),
    .O_26(n9_O_26),
    .O_27(n9_O_27),
    .O_28(n9_O_28),
    .O_29(n9_O_29),
    .O_30(n9_O_30),
    .O_31(n9_O_31),
    .O_32(n9_O_32),
    .O_33(n9_O_33),
    .O_34(n9_O_34),
    .O_35(n9_O_35),
    .O_36(n9_O_36),
    .O_37(n9_O_37),
    .O_38(n9_O_38),
    .O_39(n9_O_39),
    .O_40(n9_O_40),
    .O_41(n9_O_41),
    .O_42(n9_O_42),
    .O_43(n9_O_43),
    .O_44(n9_O_44),
    .O_45(n9_O_45),
    .O_46(n9_O_46),
    .O_47(n9_O_47),
    .O_48(n9_O_48),
    .O_49(n9_O_49),
    .O_50(n9_O_50),
    .O_51(n9_O_51),
    .O_52(n9_O_52),
    .O_53(n9_O_53),
    .O_54(n9_O_54),
    .O_55(n9_O_55),
    .O_56(n9_O_56),
    .O_57(n9_O_57),
    .O_58(n9_O_58),
    .O_59(n9_O_59),
    .O_60(n9_O_60),
    .O_61(n9_O_61),
    .O_62(n9_O_62),
    .O_63(n9_O_63),
    .O_64(n9_O_64),
    .O_65(n9_O_65),
    .O_66(n9_O_66),
    .O_67(n9_O_67),
    .O_68(n9_O_68),
    .O_69(n9_O_69),
    .O_70(n9_O_70),
    .O_71(n9_O_71),
    .O_72(n9_O_72),
    .O_73(n9_O_73),
    .O_74(n9_O_74),
    .O_75(n9_O_75),
    .O_76(n9_O_76),
    .O_77(n9_O_77),
    .O_78(n9_O_78),
    .O_79(n9_O_79),
    .O_80(n9_O_80),
    .O_81(n9_O_81),
    .O_82(n9_O_82),
    .O_83(n9_O_83),
    .O_84(n9_O_84),
    .O_85(n9_O_85),
    .O_86(n9_O_86),
    .O_87(n9_O_87),
    .O_88(n9_O_88),
    .O_89(n9_O_89),
    .O_90(n9_O_90),
    .O_91(n9_O_91),
    .O_92(n9_O_92),
    .O_93(n9_O_93),
    .O_94(n9_O_94),
    .O_95(n9_O_95),
    .O_96(n9_O_96),
    .O_97(n9_O_97),
    .O_98(n9_O_98),
    .O_99(n9_O_99),
    .O_100(n9_O_100),
    .O_101(n9_O_101),
    .O_102(n9_O_102),
    .O_103(n9_O_103),
    .O_104(n9_O_104),
    .O_105(n9_O_105),
    .O_106(n9_O_106),
    .O_107(n9_O_107),
    .O_108(n9_O_108),
    .O_109(n9_O_109),
    .O_110(n9_O_110),
    .O_111(n9_O_111),
    .O_112(n9_O_112),
    .O_113(n9_O_113),
    .O_114(n9_O_114),
    .O_115(n9_O_115),
    .O_116(n9_O_116),
    .O_117(n9_O_117),
    .O_118(n9_O_118),
    .O_119(n9_O_119),
    .O_120(n9_O_120),
    .O_121(n9_O_121),
    .O_122(n9_O_122),
    .O_123(n9_O_123),
    .O_124(n9_O_124),
    .O_125(n9_O_125),
    .O_126(n9_O_126),
    .O_127(n9_O_127),
    .O_128(n9_O_128),
    .O_129(n9_O_129),
    .O_130(n9_O_130),
    .O_131(n9_O_131),
    .O_132(n9_O_132),
    .O_133(n9_O_133),
    .O_134(n9_O_134),
    .O_135(n9_O_135),
    .O_136(n9_O_136),
    .O_137(n9_O_137),
    .O_138(n9_O_138),
    .O_139(n9_O_139),
    .O_140(n9_O_140),
    .O_141(n9_O_141),
    .O_142(n9_O_142),
    .O_143(n9_O_143),
    .O_144(n9_O_144),
    .O_145(n9_O_145),
    .O_146(n9_O_146),
    .O_147(n9_O_147),
    .O_148(n9_O_148),
    .O_149(n9_O_149),
    .O_150(n9_O_150),
    .O_151(n9_O_151),
    .O_152(n9_O_152),
    .O_153(n9_O_153),
    .O_154(n9_O_154),
    .O_155(n9_O_155),
    .O_156(n9_O_156),
    .O_157(n9_O_157),
    .O_158(n9_O_158),
    .O_159(n9_O_159),
    .O_160(n9_O_160),
    .O_161(n9_O_161),
    .O_162(n9_O_162),
    .O_163(n9_O_163),
    .O_164(n9_O_164),
    .O_165(n9_O_165),
    .O_166(n9_O_166),
    .O_167(n9_O_167),
    .O_168(n9_O_168),
    .O_169(n9_O_169),
    .O_170(n9_O_170),
    .O_171(n9_O_171),
    .O_172(n9_O_172),
    .O_173(n9_O_173),
    .O_174(n9_O_174),
    .O_175(n9_O_175),
    .O_176(n9_O_176),
    .O_177(n9_O_177),
    .O_178(n9_O_178),
    .O_179(n9_O_179),
    .O_180(n9_O_180),
    .O_181(n9_O_181),
    .O_182(n9_O_182),
    .O_183(n9_O_183),
    .O_184(n9_O_184),
    .O_185(n9_O_185),
    .O_186(n9_O_186),
    .O_187(n9_O_187),
    .O_188(n9_O_188),
    .O_189(n9_O_189),
    .O_190(n9_O_190),
    .O_191(n9_O_191),
    .O_192(n9_O_192),
    .O_193(n9_O_193),
    .O_194(n9_O_194),
    .O_195(n9_O_195),
    .O_196(n9_O_196),
    .O_197(n9_O_197),
    .O_198(n9_O_198),
    .O_199(n9_O_199)
  );
  FIFO n10 ( // @[Top.scala 44:21]
    .clock(n10_clock),
    .reset(n10_reset),
    .valid_up(n10_valid_up),
    .valid_down(n10_valid_down),
    .I_0(n10_I_0),
    .I_1(n10_I_1),
    .I_2(n10_I_2),
    .I_3(n10_I_3),
    .I_4(n10_I_4),
    .I_5(n10_I_5),
    .I_6(n10_I_6),
    .I_7(n10_I_7),
    .I_8(n10_I_8),
    .I_9(n10_I_9),
    .I_10(n10_I_10),
    .I_11(n10_I_11),
    .I_12(n10_I_12),
    .I_13(n10_I_13),
    .I_14(n10_I_14),
    .I_15(n10_I_15),
    .I_16(n10_I_16),
    .I_17(n10_I_17),
    .I_18(n10_I_18),
    .I_19(n10_I_19),
    .I_20(n10_I_20),
    .I_21(n10_I_21),
    .I_22(n10_I_22),
    .I_23(n10_I_23),
    .I_24(n10_I_24),
    .I_25(n10_I_25),
    .I_26(n10_I_26),
    .I_27(n10_I_27),
    .I_28(n10_I_28),
    .I_29(n10_I_29),
    .I_30(n10_I_30),
    .I_31(n10_I_31),
    .I_32(n10_I_32),
    .I_33(n10_I_33),
    .I_34(n10_I_34),
    .I_35(n10_I_35),
    .I_36(n10_I_36),
    .I_37(n10_I_37),
    .I_38(n10_I_38),
    .I_39(n10_I_39),
    .I_40(n10_I_40),
    .I_41(n10_I_41),
    .I_42(n10_I_42),
    .I_43(n10_I_43),
    .I_44(n10_I_44),
    .I_45(n10_I_45),
    .I_46(n10_I_46),
    .I_47(n10_I_47),
    .I_48(n10_I_48),
    .I_49(n10_I_49),
    .I_50(n10_I_50),
    .I_51(n10_I_51),
    .I_52(n10_I_52),
    .I_53(n10_I_53),
    .I_54(n10_I_54),
    .I_55(n10_I_55),
    .I_56(n10_I_56),
    .I_57(n10_I_57),
    .I_58(n10_I_58),
    .I_59(n10_I_59),
    .I_60(n10_I_60),
    .I_61(n10_I_61),
    .I_62(n10_I_62),
    .I_63(n10_I_63),
    .I_64(n10_I_64),
    .I_65(n10_I_65),
    .I_66(n10_I_66),
    .I_67(n10_I_67),
    .I_68(n10_I_68),
    .I_69(n10_I_69),
    .I_70(n10_I_70),
    .I_71(n10_I_71),
    .I_72(n10_I_72),
    .I_73(n10_I_73),
    .I_74(n10_I_74),
    .I_75(n10_I_75),
    .I_76(n10_I_76),
    .I_77(n10_I_77),
    .I_78(n10_I_78),
    .I_79(n10_I_79),
    .I_80(n10_I_80),
    .I_81(n10_I_81),
    .I_82(n10_I_82),
    .I_83(n10_I_83),
    .I_84(n10_I_84),
    .I_85(n10_I_85),
    .I_86(n10_I_86),
    .I_87(n10_I_87),
    .I_88(n10_I_88),
    .I_89(n10_I_89),
    .I_90(n10_I_90),
    .I_91(n10_I_91),
    .I_92(n10_I_92),
    .I_93(n10_I_93),
    .I_94(n10_I_94),
    .I_95(n10_I_95),
    .I_96(n10_I_96),
    .I_97(n10_I_97),
    .I_98(n10_I_98),
    .I_99(n10_I_99),
    .I_100(n10_I_100),
    .I_101(n10_I_101),
    .I_102(n10_I_102),
    .I_103(n10_I_103),
    .I_104(n10_I_104),
    .I_105(n10_I_105),
    .I_106(n10_I_106),
    .I_107(n10_I_107),
    .I_108(n10_I_108),
    .I_109(n10_I_109),
    .I_110(n10_I_110),
    .I_111(n10_I_111),
    .I_112(n10_I_112),
    .I_113(n10_I_113),
    .I_114(n10_I_114),
    .I_115(n10_I_115),
    .I_116(n10_I_116),
    .I_117(n10_I_117),
    .I_118(n10_I_118),
    .I_119(n10_I_119),
    .I_120(n10_I_120),
    .I_121(n10_I_121),
    .I_122(n10_I_122),
    .I_123(n10_I_123),
    .I_124(n10_I_124),
    .I_125(n10_I_125),
    .I_126(n10_I_126),
    .I_127(n10_I_127),
    .I_128(n10_I_128),
    .I_129(n10_I_129),
    .I_130(n10_I_130),
    .I_131(n10_I_131),
    .I_132(n10_I_132),
    .I_133(n10_I_133),
    .I_134(n10_I_134),
    .I_135(n10_I_135),
    .I_136(n10_I_136),
    .I_137(n10_I_137),
    .I_138(n10_I_138),
    .I_139(n10_I_139),
    .I_140(n10_I_140),
    .I_141(n10_I_141),
    .I_142(n10_I_142),
    .I_143(n10_I_143),
    .I_144(n10_I_144),
    .I_145(n10_I_145),
    .I_146(n10_I_146),
    .I_147(n10_I_147),
    .I_148(n10_I_148),
    .I_149(n10_I_149),
    .I_150(n10_I_150),
    .I_151(n10_I_151),
    .I_152(n10_I_152),
    .I_153(n10_I_153),
    .I_154(n10_I_154),
    .I_155(n10_I_155),
    .I_156(n10_I_156),
    .I_157(n10_I_157),
    .I_158(n10_I_158),
    .I_159(n10_I_159),
    .I_160(n10_I_160),
    .I_161(n10_I_161),
    .I_162(n10_I_162),
    .I_163(n10_I_163),
    .I_164(n10_I_164),
    .I_165(n10_I_165),
    .I_166(n10_I_166),
    .I_167(n10_I_167),
    .I_168(n10_I_168),
    .I_169(n10_I_169),
    .I_170(n10_I_170),
    .I_171(n10_I_171),
    .I_172(n10_I_172),
    .I_173(n10_I_173),
    .I_174(n10_I_174),
    .I_175(n10_I_175),
    .I_176(n10_I_176),
    .I_177(n10_I_177),
    .I_178(n10_I_178),
    .I_179(n10_I_179),
    .I_180(n10_I_180),
    .I_181(n10_I_181),
    .I_182(n10_I_182),
    .I_183(n10_I_183),
    .I_184(n10_I_184),
    .I_185(n10_I_185),
    .I_186(n10_I_186),
    .I_187(n10_I_187),
    .I_188(n10_I_188),
    .I_189(n10_I_189),
    .I_190(n10_I_190),
    .I_191(n10_I_191),
    .I_192(n10_I_192),
    .I_193(n10_I_193),
    .I_194(n10_I_194),
    .I_195(n10_I_195),
    .I_196(n10_I_196),
    .I_197(n10_I_197),
    .I_198(n10_I_198),
    .I_199(n10_I_199),
    .O_0(n10_O_0),
    .O_1(n10_O_1),
    .O_2(n10_O_2),
    .O_3(n10_O_3),
    .O_4(n10_O_4),
    .O_5(n10_O_5),
    .O_6(n10_O_6),
    .O_7(n10_O_7),
    .O_8(n10_O_8),
    .O_9(n10_O_9),
    .O_10(n10_O_10),
    .O_11(n10_O_11),
    .O_12(n10_O_12),
    .O_13(n10_O_13),
    .O_14(n10_O_14),
    .O_15(n10_O_15),
    .O_16(n10_O_16),
    .O_17(n10_O_17),
    .O_18(n10_O_18),
    .O_19(n10_O_19),
    .O_20(n10_O_20),
    .O_21(n10_O_21),
    .O_22(n10_O_22),
    .O_23(n10_O_23),
    .O_24(n10_O_24),
    .O_25(n10_O_25),
    .O_26(n10_O_26),
    .O_27(n10_O_27),
    .O_28(n10_O_28),
    .O_29(n10_O_29),
    .O_30(n10_O_30),
    .O_31(n10_O_31),
    .O_32(n10_O_32),
    .O_33(n10_O_33),
    .O_34(n10_O_34),
    .O_35(n10_O_35),
    .O_36(n10_O_36),
    .O_37(n10_O_37),
    .O_38(n10_O_38),
    .O_39(n10_O_39),
    .O_40(n10_O_40),
    .O_41(n10_O_41),
    .O_42(n10_O_42),
    .O_43(n10_O_43),
    .O_44(n10_O_44),
    .O_45(n10_O_45),
    .O_46(n10_O_46),
    .O_47(n10_O_47),
    .O_48(n10_O_48),
    .O_49(n10_O_49),
    .O_50(n10_O_50),
    .O_51(n10_O_51),
    .O_52(n10_O_52),
    .O_53(n10_O_53),
    .O_54(n10_O_54),
    .O_55(n10_O_55),
    .O_56(n10_O_56),
    .O_57(n10_O_57),
    .O_58(n10_O_58),
    .O_59(n10_O_59),
    .O_60(n10_O_60),
    .O_61(n10_O_61),
    .O_62(n10_O_62),
    .O_63(n10_O_63),
    .O_64(n10_O_64),
    .O_65(n10_O_65),
    .O_66(n10_O_66),
    .O_67(n10_O_67),
    .O_68(n10_O_68),
    .O_69(n10_O_69),
    .O_70(n10_O_70),
    .O_71(n10_O_71),
    .O_72(n10_O_72),
    .O_73(n10_O_73),
    .O_74(n10_O_74),
    .O_75(n10_O_75),
    .O_76(n10_O_76),
    .O_77(n10_O_77),
    .O_78(n10_O_78),
    .O_79(n10_O_79),
    .O_80(n10_O_80),
    .O_81(n10_O_81),
    .O_82(n10_O_82),
    .O_83(n10_O_83),
    .O_84(n10_O_84),
    .O_85(n10_O_85),
    .O_86(n10_O_86),
    .O_87(n10_O_87),
    .O_88(n10_O_88),
    .O_89(n10_O_89),
    .O_90(n10_O_90),
    .O_91(n10_O_91),
    .O_92(n10_O_92),
    .O_93(n10_O_93),
    .O_94(n10_O_94),
    .O_95(n10_O_95),
    .O_96(n10_O_96),
    .O_97(n10_O_97),
    .O_98(n10_O_98),
    .O_99(n10_O_99),
    .O_100(n10_O_100),
    .O_101(n10_O_101),
    .O_102(n10_O_102),
    .O_103(n10_O_103),
    .O_104(n10_O_104),
    .O_105(n10_O_105),
    .O_106(n10_O_106),
    .O_107(n10_O_107),
    .O_108(n10_O_108),
    .O_109(n10_O_109),
    .O_110(n10_O_110),
    .O_111(n10_O_111),
    .O_112(n10_O_112),
    .O_113(n10_O_113),
    .O_114(n10_O_114),
    .O_115(n10_O_115),
    .O_116(n10_O_116),
    .O_117(n10_O_117),
    .O_118(n10_O_118),
    .O_119(n10_O_119),
    .O_120(n10_O_120),
    .O_121(n10_O_121),
    .O_122(n10_O_122),
    .O_123(n10_O_123),
    .O_124(n10_O_124),
    .O_125(n10_O_125),
    .O_126(n10_O_126),
    .O_127(n10_O_127),
    .O_128(n10_O_128),
    .O_129(n10_O_129),
    .O_130(n10_O_130),
    .O_131(n10_O_131),
    .O_132(n10_O_132),
    .O_133(n10_O_133),
    .O_134(n10_O_134),
    .O_135(n10_O_135),
    .O_136(n10_O_136),
    .O_137(n10_O_137),
    .O_138(n10_O_138),
    .O_139(n10_O_139),
    .O_140(n10_O_140),
    .O_141(n10_O_141),
    .O_142(n10_O_142),
    .O_143(n10_O_143),
    .O_144(n10_O_144),
    .O_145(n10_O_145),
    .O_146(n10_O_146),
    .O_147(n10_O_147),
    .O_148(n10_O_148),
    .O_149(n10_O_149),
    .O_150(n10_O_150),
    .O_151(n10_O_151),
    .O_152(n10_O_152),
    .O_153(n10_O_153),
    .O_154(n10_O_154),
    .O_155(n10_O_155),
    .O_156(n10_O_156),
    .O_157(n10_O_157),
    .O_158(n10_O_158),
    .O_159(n10_O_159),
    .O_160(n10_O_160),
    .O_161(n10_O_161),
    .O_162(n10_O_162),
    .O_163(n10_O_163),
    .O_164(n10_O_164),
    .O_165(n10_O_165),
    .O_166(n10_O_166),
    .O_167(n10_O_167),
    .O_168(n10_O_168),
    .O_169(n10_O_169),
    .O_170(n10_O_170),
    .O_171(n10_O_171),
    .O_172(n10_O_172),
    .O_173(n10_O_173),
    .O_174(n10_O_174),
    .O_175(n10_O_175),
    .O_176(n10_O_176),
    .O_177(n10_O_177),
    .O_178(n10_O_178),
    .O_179(n10_O_179),
    .O_180(n10_O_180),
    .O_181(n10_O_181),
    .O_182(n10_O_182),
    .O_183(n10_O_183),
    .O_184(n10_O_184),
    .O_185(n10_O_185),
    .O_186(n10_O_186),
    .O_187(n10_O_187),
    .O_188(n10_O_188),
    .O_189(n10_O_189),
    .O_190(n10_O_190),
    .O_191(n10_O_191),
    .O_192(n10_O_192),
    .O_193(n10_O_193),
    .O_194(n10_O_194),
    .O_195(n10_O_195),
    .O_196(n10_O_196),
    .O_197(n10_O_197),
    .O_198(n10_O_198),
    .O_199(n10_O_199)
  );
  assign valid_down = n10_valid_down; // @[Top.scala 48:16]
  assign O_0 = n10_O_0; // @[Top.scala 47:7]
  assign O_1 = n10_O_1; // @[Top.scala 47:7]
  assign O_2 = n10_O_2; // @[Top.scala 47:7]
  assign O_3 = n10_O_3; // @[Top.scala 47:7]
  assign O_4 = n10_O_4; // @[Top.scala 47:7]
  assign O_5 = n10_O_5; // @[Top.scala 47:7]
  assign O_6 = n10_O_6; // @[Top.scala 47:7]
  assign O_7 = n10_O_7; // @[Top.scala 47:7]
  assign O_8 = n10_O_8; // @[Top.scala 47:7]
  assign O_9 = n10_O_9; // @[Top.scala 47:7]
  assign O_10 = n10_O_10; // @[Top.scala 47:7]
  assign O_11 = n10_O_11; // @[Top.scala 47:7]
  assign O_12 = n10_O_12; // @[Top.scala 47:7]
  assign O_13 = n10_O_13; // @[Top.scala 47:7]
  assign O_14 = n10_O_14; // @[Top.scala 47:7]
  assign O_15 = n10_O_15; // @[Top.scala 47:7]
  assign O_16 = n10_O_16; // @[Top.scala 47:7]
  assign O_17 = n10_O_17; // @[Top.scala 47:7]
  assign O_18 = n10_O_18; // @[Top.scala 47:7]
  assign O_19 = n10_O_19; // @[Top.scala 47:7]
  assign O_20 = n10_O_20; // @[Top.scala 47:7]
  assign O_21 = n10_O_21; // @[Top.scala 47:7]
  assign O_22 = n10_O_22; // @[Top.scala 47:7]
  assign O_23 = n10_O_23; // @[Top.scala 47:7]
  assign O_24 = n10_O_24; // @[Top.scala 47:7]
  assign O_25 = n10_O_25; // @[Top.scala 47:7]
  assign O_26 = n10_O_26; // @[Top.scala 47:7]
  assign O_27 = n10_O_27; // @[Top.scala 47:7]
  assign O_28 = n10_O_28; // @[Top.scala 47:7]
  assign O_29 = n10_O_29; // @[Top.scala 47:7]
  assign O_30 = n10_O_30; // @[Top.scala 47:7]
  assign O_31 = n10_O_31; // @[Top.scala 47:7]
  assign O_32 = n10_O_32; // @[Top.scala 47:7]
  assign O_33 = n10_O_33; // @[Top.scala 47:7]
  assign O_34 = n10_O_34; // @[Top.scala 47:7]
  assign O_35 = n10_O_35; // @[Top.scala 47:7]
  assign O_36 = n10_O_36; // @[Top.scala 47:7]
  assign O_37 = n10_O_37; // @[Top.scala 47:7]
  assign O_38 = n10_O_38; // @[Top.scala 47:7]
  assign O_39 = n10_O_39; // @[Top.scala 47:7]
  assign O_40 = n10_O_40; // @[Top.scala 47:7]
  assign O_41 = n10_O_41; // @[Top.scala 47:7]
  assign O_42 = n10_O_42; // @[Top.scala 47:7]
  assign O_43 = n10_O_43; // @[Top.scala 47:7]
  assign O_44 = n10_O_44; // @[Top.scala 47:7]
  assign O_45 = n10_O_45; // @[Top.scala 47:7]
  assign O_46 = n10_O_46; // @[Top.scala 47:7]
  assign O_47 = n10_O_47; // @[Top.scala 47:7]
  assign O_48 = n10_O_48; // @[Top.scala 47:7]
  assign O_49 = n10_O_49; // @[Top.scala 47:7]
  assign O_50 = n10_O_50; // @[Top.scala 47:7]
  assign O_51 = n10_O_51; // @[Top.scala 47:7]
  assign O_52 = n10_O_52; // @[Top.scala 47:7]
  assign O_53 = n10_O_53; // @[Top.scala 47:7]
  assign O_54 = n10_O_54; // @[Top.scala 47:7]
  assign O_55 = n10_O_55; // @[Top.scala 47:7]
  assign O_56 = n10_O_56; // @[Top.scala 47:7]
  assign O_57 = n10_O_57; // @[Top.scala 47:7]
  assign O_58 = n10_O_58; // @[Top.scala 47:7]
  assign O_59 = n10_O_59; // @[Top.scala 47:7]
  assign O_60 = n10_O_60; // @[Top.scala 47:7]
  assign O_61 = n10_O_61; // @[Top.scala 47:7]
  assign O_62 = n10_O_62; // @[Top.scala 47:7]
  assign O_63 = n10_O_63; // @[Top.scala 47:7]
  assign O_64 = n10_O_64; // @[Top.scala 47:7]
  assign O_65 = n10_O_65; // @[Top.scala 47:7]
  assign O_66 = n10_O_66; // @[Top.scala 47:7]
  assign O_67 = n10_O_67; // @[Top.scala 47:7]
  assign O_68 = n10_O_68; // @[Top.scala 47:7]
  assign O_69 = n10_O_69; // @[Top.scala 47:7]
  assign O_70 = n10_O_70; // @[Top.scala 47:7]
  assign O_71 = n10_O_71; // @[Top.scala 47:7]
  assign O_72 = n10_O_72; // @[Top.scala 47:7]
  assign O_73 = n10_O_73; // @[Top.scala 47:7]
  assign O_74 = n10_O_74; // @[Top.scala 47:7]
  assign O_75 = n10_O_75; // @[Top.scala 47:7]
  assign O_76 = n10_O_76; // @[Top.scala 47:7]
  assign O_77 = n10_O_77; // @[Top.scala 47:7]
  assign O_78 = n10_O_78; // @[Top.scala 47:7]
  assign O_79 = n10_O_79; // @[Top.scala 47:7]
  assign O_80 = n10_O_80; // @[Top.scala 47:7]
  assign O_81 = n10_O_81; // @[Top.scala 47:7]
  assign O_82 = n10_O_82; // @[Top.scala 47:7]
  assign O_83 = n10_O_83; // @[Top.scala 47:7]
  assign O_84 = n10_O_84; // @[Top.scala 47:7]
  assign O_85 = n10_O_85; // @[Top.scala 47:7]
  assign O_86 = n10_O_86; // @[Top.scala 47:7]
  assign O_87 = n10_O_87; // @[Top.scala 47:7]
  assign O_88 = n10_O_88; // @[Top.scala 47:7]
  assign O_89 = n10_O_89; // @[Top.scala 47:7]
  assign O_90 = n10_O_90; // @[Top.scala 47:7]
  assign O_91 = n10_O_91; // @[Top.scala 47:7]
  assign O_92 = n10_O_92; // @[Top.scala 47:7]
  assign O_93 = n10_O_93; // @[Top.scala 47:7]
  assign O_94 = n10_O_94; // @[Top.scala 47:7]
  assign O_95 = n10_O_95; // @[Top.scala 47:7]
  assign O_96 = n10_O_96; // @[Top.scala 47:7]
  assign O_97 = n10_O_97; // @[Top.scala 47:7]
  assign O_98 = n10_O_98; // @[Top.scala 47:7]
  assign O_99 = n10_O_99; // @[Top.scala 47:7]
  assign O_100 = n10_O_100; // @[Top.scala 47:7]
  assign O_101 = n10_O_101; // @[Top.scala 47:7]
  assign O_102 = n10_O_102; // @[Top.scala 47:7]
  assign O_103 = n10_O_103; // @[Top.scala 47:7]
  assign O_104 = n10_O_104; // @[Top.scala 47:7]
  assign O_105 = n10_O_105; // @[Top.scala 47:7]
  assign O_106 = n10_O_106; // @[Top.scala 47:7]
  assign O_107 = n10_O_107; // @[Top.scala 47:7]
  assign O_108 = n10_O_108; // @[Top.scala 47:7]
  assign O_109 = n10_O_109; // @[Top.scala 47:7]
  assign O_110 = n10_O_110; // @[Top.scala 47:7]
  assign O_111 = n10_O_111; // @[Top.scala 47:7]
  assign O_112 = n10_O_112; // @[Top.scala 47:7]
  assign O_113 = n10_O_113; // @[Top.scala 47:7]
  assign O_114 = n10_O_114; // @[Top.scala 47:7]
  assign O_115 = n10_O_115; // @[Top.scala 47:7]
  assign O_116 = n10_O_116; // @[Top.scala 47:7]
  assign O_117 = n10_O_117; // @[Top.scala 47:7]
  assign O_118 = n10_O_118; // @[Top.scala 47:7]
  assign O_119 = n10_O_119; // @[Top.scala 47:7]
  assign O_120 = n10_O_120; // @[Top.scala 47:7]
  assign O_121 = n10_O_121; // @[Top.scala 47:7]
  assign O_122 = n10_O_122; // @[Top.scala 47:7]
  assign O_123 = n10_O_123; // @[Top.scala 47:7]
  assign O_124 = n10_O_124; // @[Top.scala 47:7]
  assign O_125 = n10_O_125; // @[Top.scala 47:7]
  assign O_126 = n10_O_126; // @[Top.scala 47:7]
  assign O_127 = n10_O_127; // @[Top.scala 47:7]
  assign O_128 = n10_O_128; // @[Top.scala 47:7]
  assign O_129 = n10_O_129; // @[Top.scala 47:7]
  assign O_130 = n10_O_130; // @[Top.scala 47:7]
  assign O_131 = n10_O_131; // @[Top.scala 47:7]
  assign O_132 = n10_O_132; // @[Top.scala 47:7]
  assign O_133 = n10_O_133; // @[Top.scala 47:7]
  assign O_134 = n10_O_134; // @[Top.scala 47:7]
  assign O_135 = n10_O_135; // @[Top.scala 47:7]
  assign O_136 = n10_O_136; // @[Top.scala 47:7]
  assign O_137 = n10_O_137; // @[Top.scala 47:7]
  assign O_138 = n10_O_138; // @[Top.scala 47:7]
  assign O_139 = n10_O_139; // @[Top.scala 47:7]
  assign O_140 = n10_O_140; // @[Top.scala 47:7]
  assign O_141 = n10_O_141; // @[Top.scala 47:7]
  assign O_142 = n10_O_142; // @[Top.scala 47:7]
  assign O_143 = n10_O_143; // @[Top.scala 47:7]
  assign O_144 = n10_O_144; // @[Top.scala 47:7]
  assign O_145 = n10_O_145; // @[Top.scala 47:7]
  assign O_146 = n10_O_146; // @[Top.scala 47:7]
  assign O_147 = n10_O_147; // @[Top.scala 47:7]
  assign O_148 = n10_O_148; // @[Top.scala 47:7]
  assign O_149 = n10_O_149; // @[Top.scala 47:7]
  assign O_150 = n10_O_150; // @[Top.scala 47:7]
  assign O_151 = n10_O_151; // @[Top.scala 47:7]
  assign O_152 = n10_O_152; // @[Top.scala 47:7]
  assign O_153 = n10_O_153; // @[Top.scala 47:7]
  assign O_154 = n10_O_154; // @[Top.scala 47:7]
  assign O_155 = n10_O_155; // @[Top.scala 47:7]
  assign O_156 = n10_O_156; // @[Top.scala 47:7]
  assign O_157 = n10_O_157; // @[Top.scala 47:7]
  assign O_158 = n10_O_158; // @[Top.scala 47:7]
  assign O_159 = n10_O_159; // @[Top.scala 47:7]
  assign O_160 = n10_O_160; // @[Top.scala 47:7]
  assign O_161 = n10_O_161; // @[Top.scala 47:7]
  assign O_162 = n10_O_162; // @[Top.scala 47:7]
  assign O_163 = n10_O_163; // @[Top.scala 47:7]
  assign O_164 = n10_O_164; // @[Top.scala 47:7]
  assign O_165 = n10_O_165; // @[Top.scala 47:7]
  assign O_166 = n10_O_166; // @[Top.scala 47:7]
  assign O_167 = n10_O_167; // @[Top.scala 47:7]
  assign O_168 = n10_O_168; // @[Top.scala 47:7]
  assign O_169 = n10_O_169; // @[Top.scala 47:7]
  assign O_170 = n10_O_170; // @[Top.scala 47:7]
  assign O_171 = n10_O_171; // @[Top.scala 47:7]
  assign O_172 = n10_O_172; // @[Top.scala 47:7]
  assign O_173 = n10_O_173; // @[Top.scala 47:7]
  assign O_174 = n10_O_174; // @[Top.scala 47:7]
  assign O_175 = n10_O_175; // @[Top.scala 47:7]
  assign O_176 = n10_O_176; // @[Top.scala 47:7]
  assign O_177 = n10_O_177; // @[Top.scala 47:7]
  assign O_178 = n10_O_178; // @[Top.scala 47:7]
  assign O_179 = n10_O_179; // @[Top.scala 47:7]
  assign O_180 = n10_O_180; // @[Top.scala 47:7]
  assign O_181 = n10_O_181; // @[Top.scala 47:7]
  assign O_182 = n10_O_182; // @[Top.scala 47:7]
  assign O_183 = n10_O_183; // @[Top.scala 47:7]
  assign O_184 = n10_O_184; // @[Top.scala 47:7]
  assign O_185 = n10_O_185; // @[Top.scala 47:7]
  assign O_186 = n10_O_186; // @[Top.scala 47:7]
  assign O_187 = n10_O_187; // @[Top.scala 47:7]
  assign O_188 = n10_O_188; // @[Top.scala 47:7]
  assign O_189 = n10_O_189; // @[Top.scala 47:7]
  assign O_190 = n10_O_190; // @[Top.scala 47:7]
  assign O_191 = n10_O_191; // @[Top.scala 47:7]
  assign O_192 = n10_O_192; // @[Top.scala 47:7]
  assign O_193 = n10_O_193; // @[Top.scala 47:7]
  assign O_194 = n10_O_194; // @[Top.scala 47:7]
  assign O_195 = n10_O_195; // @[Top.scala 47:7]
  assign O_196 = n10_O_196; // @[Top.scala 47:7]
  assign O_197 = n10_O_197; // @[Top.scala 47:7]
  assign O_198 = n10_O_198; // @[Top.scala 47:7]
  assign O_199 = n10_O_199; // @[Top.scala 47:7]
  assign n1_clock = clock;
  assign n1_reset = reset;
  assign n1_valid_up = valid_up; // @[Top.scala 34:17]
  assign n1_I_0 = I_0; // @[Top.scala 33:10]
  assign n1_I_1 = I_1; // @[Top.scala 33:10]
  assign n1_I_2 = I_2; // @[Top.scala 33:10]
  assign n1_I_3 = I_3; // @[Top.scala 33:10]
  assign n1_I_4 = I_4; // @[Top.scala 33:10]
  assign n1_I_5 = I_5; // @[Top.scala 33:10]
  assign n1_I_6 = I_6; // @[Top.scala 33:10]
  assign n1_I_7 = I_7; // @[Top.scala 33:10]
  assign n1_I_8 = I_8; // @[Top.scala 33:10]
  assign n1_I_9 = I_9; // @[Top.scala 33:10]
  assign n1_I_10 = I_10; // @[Top.scala 33:10]
  assign n1_I_11 = I_11; // @[Top.scala 33:10]
  assign n1_I_12 = I_12; // @[Top.scala 33:10]
  assign n1_I_13 = I_13; // @[Top.scala 33:10]
  assign n1_I_14 = I_14; // @[Top.scala 33:10]
  assign n1_I_15 = I_15; // @[Top.scala 33:10]
  assign n1_I_16 = I_16; // @[Top.scala 33:10]
  assign n1_I_17 = I_17; // @[Top.scala 33:10]
  assign n1_I_18 = I_18; // @[Top.scala 33:10]
  assign n1_I_19 = I_19; // @[Top.scala 33:10]
  assign n1_I_20 = I_20; // @[Top.scala 33:10]
  assign n1_I_21 = I_21; // @[Top.scala 33:10]
  assign n1_I_22 = I_22; // @[Top.scala 33:10]
  assign n1_I_23 = I_23; // @[Top.scala 33:10]
  assign n1_I_24 = I_24; // @[Top.scala 33:10]
  assign n1_I_25 = I_25; // @[Top.scala 33:10]
  assign n1_I_26 = I_26; // @[Top.scala 33:10]
  assign n1_I_27 = I_27; // @[Top.scala 33:10]
  assign n1_I_28 = I_28; // @[Top.scala 33:10]
  assign n1_I_29 = I_29; // @[Top.scala 33:10]
  assign n1_I_30 = I_30; // @[Top.scala 33:10]
  assign n1_I_31 = I_31; // @[Top.scala 33:10]
  assign n1_I_32 = I_32; // @[Top.scala 33:10]
  assign n1_I_33 = I_33; // @[Top.scala 33:10]
  assign n1_I_34 = I_34; // @[Top.scala 33:10]
  assign n1_I_35 = I_35; // @[Top.scala 33:10]
  assign n1_I_36 = I_36; // @[Top.scala 33:10]
  assign n1_I_37 = I_37; // @[Top.scala 33:10]
  assign n1_I_38 = I_38; // @[Top.scala 33:10]
  assign n1_I_39 = I_39; // @[Top.scala 33:10]
  assign n1_I_40 = I_40; // @[Top.scala 33:10]
  assign n1_I_41 = I_41; // @[Top.scala 33:10]
  assign n1_I_42 = I_42; // @[Top.scala 33:10]
  assign n1_I_43 = I_43; // @[Top.scala 33:10]
  assign n1_I_44 = I_44; // @[Top.scala 33:10]
  assign n1_I_45 = I_45; // @[Top.scala 33:10]
  assign n1_I_46 = I_46; // @[Top.scala 33:10]
  assign n1_I_47 = I_47; // @[Top.scala 33:10]
  assign n1_I_48 = I_48; // @[Top.scala 33:10]
  assign n1_I_49 = I_49; // @[Top.scala 33:10]
  assign n1_I_50 = I_50; // @[Top.scala 33:10]
  assign n1_I_51 = I_51; // @[Top.scala 33:10]
  assign n1_I_52 = I_52; // @[Top.scala 33:10]
  assign n1_I_53 = I_53; // @[Top.scala 33:10]
  assign n1_I_54 = I_54; // @[Top.scala 33:10]
  assign n1_I_55 = I_55; // @[Top.scala 33:10]
  assign n1_I_56 = I_56; // @[Top.scala 33:10]
  assign n1_I_57 = I_57; // @[Top.scala 33:10]
  assign n1_I_58 = I_58; // @[Top.scala 33:10]
  assign n1_I_59 = I_59; // @[Top.scala 33:10]
  assign n1_I_60 = I_60; // @[Top.scala 33:10]
  assign n1_I_61 = I_61; // @[Top.scala 33:10]
  assign n1_I_62 = I_62; // @[Top.scala 33:10]
  assign n1_I_63 = I_63; // @[Top.scala 33:10]
  assign n1_I_64 = I_64; // @[Top.scala 33:10]
  assign n1_I_65 = I_65; // @[Top.scala 33:10]
  assign n1_I_66 = I_66; // @[Top.scala 33:10]
  assign n1_I_67 = I_67; // @[Top.scala 33:10]
  assign n1_I_68 = I_68; // @[Top.scala 33:10]
  assign n1_I_69 = I_69; // @[Top.scala 33:10]
  assign n1_I_70 = I_70; // @[Top.scala 33:10]
  assign n1_I_71 = I_71; // @[Top.scala 33:10]
  assign n1_I_72 = I_72; // @[Top.scala 33:10]
  assign n1_I_73 = I_73; // @[Top.scala 33:10]
  assign n1_I_74 = I_74; // @[Top.scala 33:10]
  assign n1_I_75 = I_75; // @[Top.scala 33:10]
  assign n1_I_76 = I_76; // @[Top.scala 33:10]
  assign n1_I_77 = I_77; // @[Top.scala 33:10]
  assign n1_I_78 = I_78; // @[Top.scala 33:10]
  assign n1_I_79 = I_79; // @[Top.scala 33:10]
  assign n1_I_80 = I_80; // @[Top.scala 33:10]
  assign n1_I_81 = I_81; // @[Top.scala 33:10]
  assign n1_I_82 = I_82; // @[Top.scala 33:10]
  assign n1_I_83 = I_83; // @[Top.scala 33:10]
  assign n1_I_84 = I_84; // @[Top.scala 33:10]
  assign n1_I_85 = I_85; // @[Top.scala 33:10]
  assign n1_I_86 = I_86; // @[Top.scala 33:10]
  assign n1_I_87 = I_87; // @[Top.scala 33:10]
  assign n1_I_88 = I_88; // @[Top.scala 33:10]
  assign n1_I_89 = I_89; // @[Top.scala 33:10]
  assign n1_I_90 = I_90; // @[Top.scala 33:10]
  assign n1_I_91 = I_91; // @[Top.scala 33:10]
  assign n1_I_92 = I_92; // @[Top.scala 33:10]
  assign n1_I_93 = I_93; // @[Top.scala 33:10]
  assign n1_I_94 = I_94; // @[Top.scala 33:10]
  assign n1_I_95 = I_95; // @[Top.scala 33:10]
  assign n1_I_96 = I_96; // @[Top.scala 33:10]
  assign n1_I_97 = I_97; // @[Top.scala 33:10]
  assign n1_I_98 = I_98; // @[Top.scala 33:10]
  assign n1_I_99 = I_99; // @[Top.scala 33:10]
  assign n1_I_100 = I_100; // @[Top.scala 33:10]
  assign n1_I_101 = I_101; // @[Top.scala 33:10]
  assign n1_I_102 = I_102; // @[Top.scala 33:10]
  assign n1_I_103 = I_103; // @[Top.scala 33:10]
  assign n1_I_104 = I_104; // @[Top.scala 33:10]
  assign n1_I_105 = I_105; // @[Top.scala 33:10]
  assign n1_I_106 = I_106; // @[Top.scala 33:10]
  assign n1_I_107 = I_107; // @[Top.scala 33:10]
  assign n1_I_108 = I_108; // @[Top.scala 33:10]
  assign n1_I_109 = I_109; // @[Top.scala 33:10]
  assign n1_I_110 = I_110; // @[Top.scala 33:10]
  assign n1_I_111 = I_111; // @[Top.scala 33:10]
  assign n1_I_112 = I_112; // @[Top.scala 33:10]
  assign n1_I_113 = I_113; // @[Top.scala 33:10]
  assign n1_I_114 = I_114; // @[Top.scala 33:10]
  assign n1_I_115 = I_115; // @[Top.scala 33:10]
  assign n1_I_116 = I_116; // @[Top.scala 33:10]
  assign n1_I_117 = I_117; // @[Top.scala 33:10]
  assign n1_I_118 = I_118; // @[Top.scala 33:10]
  assign n1_I_119 = I_119; // @[Top.scala 33:10]
  assign n1_I_120 = I_120; // @[Top.scala 33:10]
  assign n1_I_121 = I_121; // @[Top.scala 33:10]
  assign n1_I_122 = I_122; // @[Top.scala 33:10]
  assign n1_I_123 = I_123; // @[Top.scala 33:10]
  assign n1_I_124 = I_124; // @[Top.scala 33:10]
  assign n1_I_125 = I_125; // @[Top.scala 33:10]
  assign n1_I_126 = I_126; // @[Top.scala 33:10]
  assign n1_I_127 = I_127; // @[Top.scala 33:10]
  assign n1_I_128 = I_128; // @[Top.scala 33:10]
  assign n1_I_129 = I_129; // @[Top.scala 33:10]
  assign n1_I_130 = I_130; // @[Top.scala 33:10]
  assign n1_I_131 = I_131; // @[Top.scala 33:10]
  assign n1_I_132 = I_132; // @[Top.scala 33:10]
  assign n1_I_133 = I_133; // @[Top.scala 33:10]
  assign n1_I_134 = I_134; // @[Top.scala 33:10]
  assign n1_I_135 = I_135; // @[Top.scala 33:10]
  assign n1_I_136 = I_136; // @[Top.scala 33:10]
  assign n1_I_137 = I_137; // @[Top.scala 33:10]
  assign n1_I_138 = I_138; // @[Top.scala 33:10]
  assign n1_I_139 = I_139; // @[Top.scala 33:10]
  assign n1_I_140 = I_140; // @[Top.scala 33:10]
  assign n1_I_141 = I_141; // @[Top.scala 33:10]
  assign n1_I_142 = I_142; // @[Top.scala 33:10]
  assign n1_I_143 = I_143; // @[Top.scala 33:10]
  assign n1_I_144 = I_144; // @[Top.scala 33:10]
  assign n1_I_145 = I_145; // @[Top.scala 33:10]
  assign n1_I_146 = I_146; // @[Top.scala 33:10]
  assign n1_I_147 = I_147; // @[Top.scala 33:10]
  assign n1_I_148 = I_148; // @[Top.scala 33:10]
  assign n1_I_149 = I_149; // @[Top.scala 33:10]
  assign n1_I_150 = I_150; // @[Top.scala 33:10]
  assign n1_I_151 = I_151; // @[Top.scala 33:10]
  assign n1_I_152 = I_152; // @[Top.scala 33:10]
  assign n1_I_153 = I_153; // @[Top.scala 33:10]
  assign n1_I_154 = I_154; // @[Top.scala 33:10]
  assign n1_I_155 = I_155; // @[Top.scala 33:10]
  assign n1_I_156 = I_156; // @[Top.scala 33:10]
  assign n1_I_157 = I_157; // @[Top.scala 33:10]
  assign n1_I_158 = I_158; // @[Top.scala 33:10]
  assign n1_I_159 = I_159; // @[Top.scala 33:10]
  assign n1_I_160 = I_160; // @[Top.scala 33:10]
  assign n1_I_161 = I_161; // @[Top.scala 33:10]
  assign n1_I_162 = I_162; // @[Top.scala 33:10]
  assign n1_I_163 = I_163; // @[Top.scala 33:10]
  assign n1_I_164 = I_164; // @[Top.scala 33:10]
  assign n1_I_165 = I_165; // @[Top.scala 33:10]
  assign n1_I_166 = I_166; // @[Top.scala 33:10]
  assign n1_I_167 = I_167; // @[Top.scala 33:10]
  assign n1_I_168 = I_168; // @[Top.scala 33:10]
  assign n1_I_169 = I_169; // @[Top.scala 33:10]
  assign n1_I_170 = I_170; // @[Top.scala 33:10]
  assign n1_I_171 = I_171; // @[Top.scala 33:10]
  assign n1_I_172 = I_172; // @[Top.scala 33:10]
  assign n1_I_173 = I_173; // @[Top.scala 33:10]
  assign n1_I_174 = I_174; // @[Top.scala 33:10]
  assign n1_I_175 = I_175; // @[Top.scala 33:10]
  assign n1_I_176 = I_176; // @[Top.scala 33:10]
  assign n1_I_177 = I_177; // @[Top.scala 33:10]
  assign n1_I_178 = I_178; // @[Top.scala 33:10]
  assign n1_I_179 = I_179; // @[Top.scala 33:10]
  assign n1_I_180 = I_180; // @[Top.scala 33:10]
  assign n1_I_181 = I_181; // @[Top.scala 33:10]
  assign n1_I_182 = I_182; // @[Top.scala 33:10]
  assign n1_I_183 = I_183; // @[Top.scala 33:10]
  assign n1_I_184 = I_184; // @[Top.scala 33:10]
  assign n1_I_185 = I_185; // @[Top.scala 33:10]
  assign n1_I_186 = I_186; // @[Top.scala 33:10]
  assign n1_I_187 = I_187; // @[Top.scala 33:10]
  assign n1_I_188 = I_188; // @[Top.scala 33:10]
  assign n1_I_189 = I_189; // @[Top.scala 33:10]
  assign n1_I_190 = I_190; // @[Top.scala 33:10]
  assign n1_I_191 = I_191; // @[Top.scala 33:10]
  assign n1_I_192 = I_192; // @[Top.scala 33:10]
  assign n1_I_193 = I_193; // @[Top.scala 33:10]
  assign n1_I_194 = I_194; // @[Top.scala 33:10]
  assign n1_I_195 = I_195; // @[Top.scala 33:10]
  assign n1_I_196 = I_196; // @[Top.scala 33:10]
  assign n1_I_197 = I_197; // @[Top.scala 33:10]
  assign n1_I_198 = I_198; // @[Top.scala 33:10]
  assign n1_I_199 = I_199; // @[Top.scala 33:10]
  assign n7_clock = clock;
  assign n7_reset = reset;
  assign n7_valid_up = n1_valid_down; // @[Top.scala 37:17]
  assign n7_I_0 = n1_O_0; // @[Top.scala 36:10]
  assign n7_I_1 = n1_O_1; // @[Top.scala 36:10]
  assign n7_I_2 = n1_O_2; // @[Top.scala 36:10]
  assign n7_I_3 = n1_O_3; // @[Top.scala 36:10]
  assign n7_I_4 = n1_O_4; // @[Top.scala 36:10]
  assign n7_I_5 = n1_O_5; // @[Top.scala 36:10]
  assign n7_I_6 = n1_O_6; // @[Top.scala 36:10]
  assign n7_I_7 = n1_O_7; // @[Top.scala 36:10]
  assign n7_I_8 = n1_O_8; // @[Top.scala 36:10]
  assign n7_I_9 = n1_O_9; // @[Top.scala 36:10]
  assign n7_I_10 = n1_O_10; // @[Top.scala 36:10]
  assign n7_I_11 = n1_O_11; // @[Top.scala 36:10]
  assign n7_I_12 = n1_O_12; // @[Top.scala 36:10]
  assign n7_I_13 = n1_O_13; // @[Top.scala 36:10]
  assign n7_I_14 = n1_O_14; // @[Top.scala 36:10]
  assign n7_I_15 = n1_O_15; // @[Top.scala 36:10]
  assign n7_I_16 = n1_O_16; // @[Top.scala 36:10]
  assign n7_I_17 = n1_O_17; // @[Top.scala 36:10]
  assign n7_I_18 = n1_O_18; // @[Top.scala 36:10]
  assign n7_I_19 = n1_O_19; // @[Top.scala 36:10]
  assign n7_I_20 = n1_O_20; // @[Top.scala 36:10]
  assign n7_I_21 = n1_O_21; // @[Top.scala 36:10]
  assign n7_I_22 = n1_O_22; // @[Top.scala 36:10]
  assign n7_I_23 = n1_O_23; // @[Top.scala 36:10]
  assign n7_I_24 = n1_O_24; // @[Top.scala 36:10]
  assign n7_I_25 = n1_O_25; // @[Top.scala 36:10]
  assign n7_I_26 = n1_O_26; // @[Top.scala 36:10]
  assign n7_I_27 = n1_O_27; // @[Top.scala 36:10]
  assign n7_I_28 = n1_O_28; // @[Top.scala 36:10]
  assign n7_I_29 = n1_O_29; // @[Top.scala 36:10]
  assign n7_I_30 = n1_O_30; // @[Top.scala 36:10]
  assign n7_I_31 = n1_O_31; // @[Top.scala 36:10]
  assign n7_I_32 = n1_O_32; // @[Top.scala 36:10]
  assign n7_I_33 = n1_O_33; // @[Top.scala 36:10]
  assign n7_I_34 = n1_O_34; // @[Top.scala 36:10]
  assign n7_I_35 = n1_O_35; // @[Top.scala 36:10]
  assign n7_I_36 = n1_O_36; // @[Top.scala 36:10]
  assign n7_I_37 = n1_O_37; // @[Top.scala 36:10]
  assign n7_I_38 = n1_O_38; // @[Top.scala 36:10]
  assign n7_I_39 = n1_O_39; // @[Top.scala 36:10]
  assign n7_I_40 = n1_O_40; // @[Top.scala 36:10]
  assign n7_I_41 = n1_O_41; // @[Top.scala 36:10]
  assign n7_I_42 = n1_O_42; // @[Top.scala 36:10]
  assign n7_I_43 = n1_O_43; // @[Top.scala 36:10]
  assign n7_I_44 = n1_O_44; // @[Top.scala 36:10]
  assign n7_I_45 = n1_O_45; // @[Top.scala 36:10]
  assign n7_I_46 = n1_O_46; // @[Top.scala 36:10]
  assign n7_I_47 = n1_O_47; // @[Top.scala 36:10]
  assign n7_I_48 = n1_O_48; // @[Top.scala 36:10]
  assign n7_I_49 = n1_O_49; // @[Top.scala 36:10]
  assign n7_I_50 = n1_O_50; // @[Top.scala 36:10]
  assign n7_I_51 = n1_O_51; // @[Top.scala 36:10]
  assign n7_I_52 = n1_O_52; // @[Top.scala 36:10]
  assign n7_I_53 = n1_O_53; // @[Top.scala 36:10]
  assign n7_I_54 = n1_O_54; // @[Top.scala 36:10]
  assign n7_I_55 = n1_O_55; // @[Top.scala 36:10]
  assign n7_I_56 = n1_O_56; // @[Top.scala 36:10]
  assign n7_I_57 = n1_O_57; // @[Top.scala 36:10]
  assign n7_I_58 = n1_O_58; // @[Top.scala 36:10]
  assign n7_I_59 = n1_O_59; // @[Top.scala 36:10]
  assign n7_I_60 = n1_O_60; // @[Top.scala 36:10]
  assign n7_I_61 = n1_O_61; // @[Top.scala 36:10]
  assign n7_I_62 = n1_O_62; // @[Top.scala 36:10]
  assign n7_I_63 = n1_O_63; // @[Top.scala 36:10]
  assign n7_I_64 = n1_O_64; // @[Top.scala 36:10]
  assign n7_I_65 = n1_O_65; // @[Top.scala 36:10]
  assign n7_I_66 = n1_O_66; // @[Top.scala 36:10]
  assign n7_I_67 = n1_O_67; // @[Top.scala 36:10]
  assign n7_I_68 = n1_O_68; // @[Top.scala 36:10]
  assign n7_I_69 = n1_O_69; // @[Top.scala 36:10]
  assign n7_I_70 = n1_O_70; // @[Top.scala 36:10]
  assign n7_I_71 = n1_O_71; // @[Top.scala 36:10]
  assign n7_I_72 = n1_O_72; // @[Top.scala 36:10]
  assign n7_I_73 = n1_O_73; // @[Top.scala 36:10]
  assign n7_I_74 = n1_O_74; // @[Top.scala 36:10]
  assign n7_I_75 = n1_O_75; // @[Top.scala 36:10]
  assign n7_I_76 = n1_O_76; // @[Top.scala 36:10]
  assign n7_I_77 = n1_O_77; // @[Top.scala 36:10]
  assign n7_I_78 = n1_O_78; // @[Top.scala 36:10]
  assign n7_I_79 = n1_O_79; // @[Top.scala 36:10]
  assign n7_I_80 = n1_O_80; // @[Top.scala 36:10]
  assign n7_I_81 = n1_O_81; // @[Top.scala 36:10]
  assign n7_I_82 = n1_O_82; // @[Top.scala 36:10]
  assign n7_I_83 = n1_O_83; // @[Top.scala 36:10]
  assign n7_I_84 = n1_O_84; // @[Top.scala 36:10]
  assign n7_I_85 = n1_O_85; // @[Top.scala 36:10]
  assign n7_I_86 = n1_O_86; // @[Top.scala 36:10]
  assign n7_I_87 = n1_O_87; // @[Top.scala 36:10]
  assign n7_I_88 = n1_O_88; // @[Top.scala 36:10]
  assign n7_I_89 = n1_O_89; // @[Top.scala 36:10]
  assign n7_I_90 = n1_O_90; // @[Top.scala 36:10]
  assign n7_I_91 = n1_O_91; // @[Top.scala 36:10]
  assign n7_I_92 = n1_O_92; // @[Top.scala 36:10]
  assign n7_I_93 = n1_O_93; // @[Top.scala 36:10]
  assign n7_I_94 = n1_O_94; // @[Top.scala 36:10]
  assign n7_I_95 = n1_O_95; // @[Top.scala 36:10]
  assign n7_I_96 = n1_O_96; // @[Top.scala 36:10]
  assign n7_I_97 = n1_O_97; // @[Top.scala 36:10]
  assign n7_I_98 = n1_O_98; // @[Top.scala 36:10]
  assign n7_I_99 = n1_O_99; // @[Top.scala 36:10]
  assign n7_I_100 = n1_O_100; // @[Top.scala 36:10]
  assign n7_I_101 = n1_O_101; // @[Top.scala 36:10]
  assign n7_I_102 = n1_O_102; // @[Top.scala 36:10]
  assign n7_I_103 = n1_O_103; // @[Top.scala 36:10]
  assign n7_I_104 = n1_O_104; // @[Top.scala 36:10]
  assign n7_I_105 = n1_O_105; // @[Top.scala 36:10]
  assign n7_I_106 = n1_O_106; // @[Top.scala 36:10]
  assign n7_I_107 = n1_O_107; // @[Top.scala 36:10]
  assign n7_I_108 = n1_O_108; // @[Top.scala 36:10]
  assign n7_I_109 = n1_O_109; // @[Top.scala 36:10]
  assign n7_I_110 = n1_O_110; // @[Top.scala 36:10]
  assign n7_I_111 = n1_O_111; // @[Top.scala 36:10]
  assign n7_I_112 = n1_O_112; // @[Top.scala 36:10]
  assign n7_I_113 = n1_O_113; // @[Top.scala 36:10]
  assign n7_I_114 = n1_O_114; // @[Top.scala 36:10]
  assign n7_I_115 = n1_O_115; // @[Top.scala 36:10]
  assign n7_I_116 = n1_O_116; // @[Top.scala 36:10]
  assign n7_I_117 = n1_O_117; // @[Top.scala 36:10]
  assign n7_I_118 = n1_O_118; // @[Top.scala 36:10]
  assign n7_I_119 = n1_O_119; // @[Top.scala 36:10]
  assign n7_I_120 = n1_O_120; // @[Top.scala 36:10]
  assign n7_I_121 = n1_O_121; // @[Top.scala 36:10]
  assign n7_I_122 = n1_O_122; // @[Top.scala 36:10]
  assign n7_I_123 = n1_O_123; // @[Top.scala 36:10]
  assign n7_I_124 = n1_O_124; // @[Top.scala 36:10]
  assign n7_I_125 = n1_O_125; // @[Top.scala 36:10]
  assign n7_I_126 = n1_O_126; // @[Top.scala 36:10]
  assign n7_I_127 = n1_O_127; // @[Top.scala 36:10]
  assign n7_I_128 = n1_O_128; // @[Top.scala 36:10]
  assign n7_I_129 = n1_O_129; // @[Top.scala 36:10]
  assign n7_I_130 = n1_O_130; // @[Top.scala 36:10]
  assign n7_I_131 = n1_O_131; // @[Top.scala 36:10]
  assign n7_I_132 = n1_O_132; // @[Top.scala 36:10]
  assign n7_I_133 = n1_O_133; // @[Top.scala 36:10]
  assign n7_I_134 = n1_O_134; // @[Top.scala 36:10]
  assign n7_I_135 = n1_O_135; // @[Top.scala 36:10]
  assign n7_I_136 = n1_O_136; // @[Top.scala 36:10]
  assign n7_I_137 = n1_O_137; // @[Top.scala 36:10]
  assign n7_I_138 = n1_O_138; // @[Top.scala 36:10]
  assign n7_I_139 = n1_O_139; // @[Top.scala 36:10]
  assign n7_I_140 = n1_O_140; // @[Top.scala 36:10]
  assign n7_I_141 = n1_O_141; // @[Top.scala 36:10]
  assign n7_I_142 = n1_O_142; // @[Top.scala 36:10]
  assign n7_I_143 = n1_O_143; // @[Top.scala 36:10]
  assign n7_I_144 = n1_O_144; // @[Top.scala 36:10]
  assign n7_I_145 = n1_O_145; // @[Top.scala 36:10]
  assign n7_I_146 = n1_O_146; // @[Top.scala 36:10]
  assign n7_I_147 = n1_O_147; // @[Top.scala 36:10]
  assign n7_I_148 = n1_O_148; // @[Top.scala 36:10]
  assign n7_I_149 = n1_O_149; // @[Top.scala 36:10]
  assign n7_I_150 = n1_O_150; // @[Top.scala 36:10]
  assign n7_I_151 = n1_O_151; // @[Top.scala 36:10]
  assign n7_I_152 = n1_O_152; // @[Top.scala 36:10]
  assign n7_I_153 = n1_O_153; // @[Top.scala 36:10]
  assign n7_I_154 = n1_O_154; // @[Top.scala 36:10]
  assign n7_I_155 = n1_O_155; // @[Top.scala 36:10]
  assign n7_I_156 = n1_O_156; // @[Top.scala 36:10]
  assign n7_I_157 = n1_O_157; // @[Top.scala 36:10]
  assign n7_I_158 = n1_O_158; // @[Top.scala 36:10]
  assign n7_I_159 = n1_O_159; // @[Top.scala 36:10]
  assign n7_I_160 = n1_O_160; // @[Top.scala 36:10]
  assign n7_I_161 = n1_O_161; // @[Top.scala 36:10]
  assign n7_I_162 = n1_O_162; // @[Top.scala 36:10]
  assign n7_I_163 = n1_O_163; // @[Top.scala 36:10]
  assign n7_I_164 = n1_O_164; // @[Top.scala 36:10]
  assign n7_I_165 = n1_O_165; // @[Top.scala 36:10]
  assign n7_I_166 = n1_O_166; // @[Top.scala 36:10]
  assign n7_I_167 = n1_O_167; // @[Top.scala 36:10]
  assign n7_I_168 = n1_O_168; // @[Top.scala 36:10]
  assign n7_I_169 = n1_O_169; // @[Top.scala 36:10]
  assign n7_I_170 = n1_O_170; // @[Top.scala 36:10]
  assign n7_I_171 = n1_O_171; // @[Top.scala 36:10]
  assign n7_I_172 = n1_O_172; // @[Top.scala 36:10]
  assign n7_I_173 = n1_O_173; // @[Top.scala 36:10]
  assign n7_I_174 = n1_O_174; // @[Top.scala 36:10]
  assign n7_I_175 = n1_O_175; // @[Top.scala 36:10]
  assign n7_I_176 = n1_O_176; // @[Top.scala 36:10]
  assign n7_I_177 = n1_O_177; // @[Top.scala 36:10]
  assign n7_I_178 = n1_O_178; // @[Top.scala 36:10]
  assign n7_I_179 = n1_O_179; // @[Top.scala 36:10]
  assign n7_I_180 = n1_O_180; // @[Top.scala 36:10]
  assign n7_I_181 = n1_O_181; // @[Top.scala 36:10]
  assign n7_I_182 = n1_O_182; // @[Top.scala 36:10]
  assign n7_I_183 = n1_O_183; // @[Top.scala 36:10]
  assign n7_I_184 = n1_O_184; // @[Top.scala 36:10]
  assign n7_I_185 = n1_O_185; // @[Top.scala 36:10]
  assign n7_I_186 = n1_O_186; // @[Top.scala 36:10]
  assign n7_I_187 = n1_O_187; // @[Top.scala 36:10]
  assign n7_I_188 = n1_O_188; // @[Top.scala 36:10]
  assign n7_I_189 = n1_O_189; // @[Top.scala 36:10]
  assign n7_I_190 = n1_O_190; // @[Top.scala 36:10]
  assign n7_I_191 = n1_O_191; // @[Top.scala 36:10]
  assign n7_I_192 = n1_O_192; // @[Top.scala 36:10]
  assign n7_I_193 = n1_O_193; // @[Top.scala 36:10]
  assign n7_I_194 = n1_O_194; // @[Top.scala 36:10]
  assign n7_I_195 = n1_O_195; // @[Top.scala 36:10]
  assign n7_I_196 = n1_O_196; // @[Top.scala 36:10]
  assign n7_I_197 = n1_O_197; // @[Top.scala 36:10]
  assign n7_I_198 = n1_O_198; // @[Top.scala 36:10]
  assign n7_I_199 = n1_O_199; // @[Top.scala 36:10]
  assign n8_clock = clock;
  assign n8_reset = reset;
  assign n8_valid_up = n7_valid_down; // @[Top.scala 40:17]
  assign n8_I_0 = n7_O_0; // @[Top.scala 39:10]
  assign n8_I_1 = n7_O_1; // @[Top.scala 39:10]
  assign n8_I_2 = n7_O_2; // @[Top.scala 39:10]
  assign n8_I_3 = n7_O_3; // @[Top.scala 39:10]
  assign n8_I_4 = n7_O_4; // @[Top.scala 39:10]
  assign n8_I_5 = n7_O_5; // @[Top.scala 39:10]
  assign n8_I_6 = n7_O_6; // @[Top.scala 39:10]
  assign n8_I_7 = n7_O_7; // @[Top.scala 39:10]
  assign n8_I_8 = n7_O_8; // @[Top.scala 39:10]
  assign n8_I_9 = n7_O_9; // @[Top.scala 39:10]
  assign n8_I_10 = n7_O_10; // @[Top.scala 39:10]
  assign n8_I_11 = n7_O_11; // @[Top.scala 39:10]
  assign n8_I_12 = n7_O_12; // @[Top.scala 39:10]
  assign n8_I_13 = n7_O_13; // @[Top.scala 39:10]
  assign n8_I_14 = n7_O_14; // @[Top.scala 39:10]
  assign n8_I_15 = n7_O_15; // @[Top.scala 39:10]
  assign n8_I_16 = n7_O_16; // @[Top.scala 39:10]
  assign n8_I_17 = n7_O_17; // @[Top.scala 39:10]
  assign n8_I_18 = n7_O_18; // @[Top.scala 39:10]
  assign n8_I_19 = n7_O_19; // @[Top.scala 39:10]
  assign n8_I_20 = n7_O_20; // @[Top.scala 39:10]
  assign n8_I_21 = n7_O_21; // @[Top.scala 39:10]
  assign n8_I_22 = n7_O_22; // @[Top.scala 39:10]
  assign n8_I_23 = n7_O_23; // @[Top.scala 39:10]
  assign n8_I_24 = n7_O_24; // @[Top.scala 39:10]
  assign n8_I_25 = n7_O_25; // @[Top.scala 39:10]
  assign n8_I_26 = n7_O_26; // @[Top.scala 39:10]
  assign n8_I_27 = n7_O_27; // @[Top.scala 39:10]
  assign n8_I_28 = n7_O_28; // @[Top.scala 39:10]
  assign n8_I_29 = n7_O_29; // @[Top.scala 39:10]
  assign n8_I_30 = n7_O_30; // @[Top.scala 39:10]
  assign n8_I_31 = n7_O_31; // @[Top.scala 39:10]
  assign n8_I_32 = n7_O_32; // @[Top.scala 39:10]
  assign n8_I_33 = n7_O_33; // @[Top.scala 39:10]
  assign n8_I_34 = n7_O_34; // @[Top.scala 39:10]
  assign n8_I_35 = n7_O_35; // @[Top.scala 39:10]
  assign n8_I_36 = n7_O_36; // @[Top.scala 39:10]
  assign n8_I_37 = n7_O_37; // @[Top.scala 39:10]
  assign n8_I_38 = n7_O_38; // @[Top.scala 39:10]
  assign n8_I_39 = n7_O_39; // @[Top.scala 39:10]
  assign n8_I_40 = n7_O_40; // @[Top.scala 39:10]
  assign n8_I_41 = n7_O_41; // @[Top.scala 39:10]
  assign n8_I_42 = n7_O_42; // @[Top.scala 39:10]
  assign n8_I_43 = n7_O_43; // @[Top.scala 39:10]
  assign n8_I_44 = n7_O_44; // @[Top.scala 39:10]
  assign n8_I_45 = n7_O_45; // @[Top.scala 39:10]
  assign n8_I_46 = n7_O_46; // @[Top.scala 39:10]
  assign n8_I_47 = n7_O_47; // @[Top.scala 39:10]
  assign n8_I_48 = n7_O_48; // @[Top.scala 39:10]
  assign n8_I_49 = n7_O_49; // @[Top.scala 39:10]
  assign n8_I_50 = n7_O_50; // @[Top.scala 39:10]
  assign n8_I_51 = n7_O_51; // @[Top.scala 39:10]
  assign n8_I_52 = n7_O_52; // @[Top.scala 39:10]
  assign n8_I_53 = n7_O_53; // @[Top.scala 39:10]
  assign n8_I_54 = n7_O_54; // @[Top.scala 39:10]
  assign n8_I_55 = n7_O_55; // @[Top.scala 39:10]
  assign n8_I_56 = n7_O_56; // @[Top.scala 39:10]
  assign n8_I_57 = n7_O_57; // @[Top.scala 39:10]
  assign n8_I_58 = n7_O_58; // @[Top.scala 39:10]
  assign n8_I_59 = n7_O_59; // @[Top.scala 39:10]
  assign n8_I_60 = n7_O_60; // @[Top.scala 39:10]
  assign n8_I_61 = n7_O_61; // @[Top.scala 39:10]
  assign n8_I_62 = n7_O_62; // @[Top.scala 39:10]
  assign n8_I_63 = n7_O_63; // @[Top.scala 39:10]
  assign n8_I_64 = n7_O_64; // @[Top.scala 39:10]
  assign n8_I_65 = n7_O_65; // @[Top.scala 39:10]
  assign n8_I_66 = n7_O_66; // @[Top.scala 39:10]
  assign n8_I_67 = n7_O_67; // @[Top.scala 39:10]
  assign n8_I_68 = n7_O_68; // @[Top.scala 39:10]
  assign n8_I_69 = n7_O_69; // @[Top.scala 39:10]
  assign n8_I_70 = n7_O_70; // @[Top.scala 39:10]
  assign n8_I_71 = n7_O_71; // @[Top.scala 39:10]
  assign n8_I_72 = n7_O_72; // @[Top.scala 39:10]
  assign n8_I_73 = n7_O_73; // @[Top.scala 39:10]
  assign n8_I_74 = n7_O_74; // @[Top.scala 39:10]
  assign n8_I_75 = n7_O_75; // @[Top.scala 39:10]
  assign n8_I_76 = n7_O_76; // @[Top.scala 39:10]
  assign n8_I_77 = n7_O_77; // @[Top.scala 39:10]
  assign n8_I_78 = n7_O_78; // @[Top.scala 39:10]
  assign n8_I_79 = n7_O_79; // @[Top.scala 39:10]
  assign n8_I_80 = n7_O_80; // @[Top.scala 39:10]
  assign n8_I_81 = n7_O_81; // @[Top.scala 39:10]
  assign n8_I_82 = n7_O_82; // @[Top.scala 39:10]
  assign n8_I_83 = n7_O_83; // @[Top.scala 39:10]
  assign n8_I_84 = n7_O_84; // @[Top.scala 39:10]
  assign n8_I_85 = n7_O_85; // @[Top.scala 39:10]
  assign n8_I_86 = n7_O_86; // @[Top.scala 39:10]
  assign n8_I_87 = n7_O_87; // @[Top.scala 39:10]
  assign n8_I_88 = n7_O_88; // @[Top.scala 39:10]
  assign n8_I_89 = n7_O_89; // @[Top.scala 39:10]
  assign n8_I_90 = n7_O_90; // @[Top.scala 39:10]
  assign n8_I_91 = n7_O_91; // @[Top.scala 39:10]
  assign n8_I_92 = n7_O_92; // @[Top.scala 39:10]
  assign n8_I_93 = n7_O_93; // @[Top.scala 39:10]
  assign n8_I_94 = n7_O_94; // @[Top.scala 39:10]
  assign n8_I_95 = n7_O_95; // @[Top.scala 39:10]
  assign n8_I_96 = n7_O_96; // @[Top.scala 39:10]
  assign n8_I_97 = n7_O_97; // @[Top.scala 39:10]
  assign n8_I_98 = n7_O_98; // @[Top.scala 39:10]
  assign n8_I_99 = n7_O_99; // @[Top.scala 39:10]
  assign n8_I_100 = n7_O_100; // @[Top.scala 39:10]
  assign n8_I_101 = n7_O_101; // @[Top.scala 39:10]
  assign n8_I_102 = n7_O_102; // @[Top.scala 39:10]
  assign n8_I_103 = n7_O_103; // @[Top.scala 39:10]
  assign n8_I_104 = n7_O_104; // @[Top.scala 39:10]
  assign n8_I_105 = n7_O_105; // @[Top.scala 39:10]
  assign n8_I_106 = n7_O_106; // @[Top.scala 39:10]
  assign n8_I_107 = n7_O_107; // @[Top.scala 39:10]
  assign n8_I_108 = n7_O_108; // @[Top.scala 39:10]
  assign n8_I_109 = n7_O_109; // @[Top.scala 39:10]
  assign n8_I_110 = n7_O_110; // @[Top.scala 39:10]
  assign n8_I_111 = n7_O_111; // @[Top.scala 39:10]
  assign n8_I_112 = n7_O_112; // @[Top.scala 39:10]
  assign n8_I_113 = n7_O_113; // @[Top.scala 39:10]
  assign n8_I_114 = n7_O_114; // @[Top.scala 39:10]
  assign n8_I_115 = n7_O_115; // @[Top.scala 39:10]
  assign n8_I_116 = n7_O_116; // @[Top.scala 39:10]
  assign n8_I_117 = n7_O_117; // @[Top.scala 39:10]
  assign n8_I_118 = n7_O_118; // @[Top.scala 39:10]
  assign n8_I_119 = n7_O_119; // @[Top.scala 39:10]
  assign n8_I_120 = n7_O_120; // @[Top.scala 39:10]
  assign n8_I_121 = n7_O_121; // @[Top.scala 39:10]
  assign n8_I_122 = n7_O_122; // @[Top.scala 39:10]
  assign n8_I_123 = n7_O_123; // @[Top.scala 39:10]
  assign n8_I_124 = n7_O_124; // @[Top.scala 39:10]
  assign n8_I_125 = n7_O_125; // @[Top.scala 39:10]
  assign n8_I_126 = n7_O_126; // @[Top.scala 39:10]
  assign n8_I_127 = n7_O_127; // @[Top.scala 39:10]
  assign n8_I_128 = n7_O_128; // @[Top.scala 39:10]
  assign n8_I_129 = n7_O_129; // @[Top.scala 39:10]
  assign n8_I_130 = n7_O_130; // @[Top.scala 39:10]
  assign n8_I_131 = n7_O_131; // @[Top.scala 39:10]
  assign n8_I_132 = n7_O_132; // @[Top.scala 39:10]
  assign n8_I_133 = n7_O_133; // @[Top.scala 39:10]
  assign n8_I_134 = n7_O_134; // @[Top.scala 39:10]
  assign n8_I_135 = n7_O_135; // @[Top.scala 39:10]
  assign n8_I_136 = n7_O_136; // @[Top.scala 39:10]
  assign n8_I_137 = n7_O_137; // @[Top.scala 39:10]
  assign n8_I_138 = n7_O_138; // @[Top.scala 39:10]
  assign n8_I_139 = n7_O_139; // @[Top.scala 39:10]
  assign n8_I_140 = n7_O_140; // @[Top.scala 39:10]
  assign n8_I_141 = n7_O_141; // @[Top.scala 39:10]
  assign n8_I_142 = n7_O_142; // @[Top.scala 39:10]
  assign n8_I_143 = n7_O_143; // @[Top.scala 39:10]
  assign n8_I_144 = n7_O_144; // @[Top.scala 39:10]
  assign n8_I_145 = n7_O_145; // @[Top.scala 39:10]
  assign n8_I_146 = n7_O_146; // @[Top.scala 39:10]
  assign n8_I_147 = n7_O_147; // @[Top.scala 39:10]
  assign n8_I_148 = n7_O_148; // @[Top.scala 39:10]
  assign n8_I_149 = n7_O_149; // @[Top.scala 39:10]
  assign n8_I_150 = n7_O_150; // @[Top.scala 39:10]
  assign n8_I_151 = n7_O_151; // @[Top.scala 39:10]
  assign n8_I_152 = n7_O_152; // @[Top.scala 39:10]
  assign n8_I_153 = n7_O_153; // @[Top.scala 39:10]
  assign n8_I_154 = n7_O_154; // @[Top.scala 39:10]
  assign n8_I_155 = n7_O_155; // @[Top.scala 39:10]
  assign n8_I_156 = n7_O_156; // @[Top.scala 39:10]
  assign n8_I_157 = n7_O_157; // @[Top.scala 39:10]
  assign n8_I_158 = n7_O_158; // @[Top.scala 39:10]
  assign n8_I_159 = n7_O_159; // @[Top.scala 39:10]
  assign n8_I_160 = n7_O_160; // @[Top.scala 39:10]
  assign n8_I_161 = n7_O_161; // @[Top.scala 39:10]
  assign n8_I_162 = n7_O_162; // @[Top.scala 39:10]
  assign n8_I_163 = n7_O_163; // @[Top.scala 39:10]
  assign n8_I_164 = n7_O_164; // @[Top.scala 39:10]
  assign n8_I_165 = n7_O_165; // @[Top.scala 39:10]
  assign n8_I_166 = n7_O_166; // @[Top.scala 39:10]
  assign n8_I_167 = n7_O_167; // @[Top.scala 39:10]
  assign n8_I_168 = n7_O_168; // @[Top.scala 39:10]
  assign n8_I_169 = n7_O_169; // @[Top.scala 39:10]
  assign n8_I_170 = n7_O_170; // @[Top.scala 39:10]
  assign n8_I_171 = n7_O_171; // @[Top.scala 39:10]
  assign n8_I_172 = n7_O_172; // @[Top.scala 39:10]
  assign n8_I_173 = n7_O_173; // @[Top.scala 39:10]
  assign n8_I_174 = n7_O_174; // @[Top.scala 39:10]
  assign n8_I_175 = n7_O_175; // @[Top.scala 39:10]
  assign n8_I_176 = n7_O_176; // @[Top.scala 39:10]
  assign n8_I_177 = n7_O_177; // @[Top.scala 39:10]
  assign n8_I_178 = n7_O_178; // @[Top.scala 39:10]
  assign n8_I_179 = n7_O_179; // @[Top.scala 39:10]
  assign n8_I_180 = n7_O_180; // @[Top.scala 39:10]
  assign n8_I_181 = n7_O_181; // @[Top.scala 39:10]
  assign n8_I_182 = n7_O_182; // @[Top.scala 39:10]
  assign n8_I_183 = n7_O_183; // @[Top.scala 39:10]
  assign n8_I_184 = n7_O_184; // @[Top.scala 39:10]
  assign n8_I_185 = n7_O_185; // @[Top.scala 39:10]
  assign n8_I_186 = n7_O_186; // @[Top.scala 39:10]
  assign n8_I_187 = n7_O_187; // @[Top.scala 39:10]
  assign n8_I_188 = n7_O_188; // @[Top.scala 39:10]
  assign n8_I_189 = n7_O_189; // @[Top.scala 39:10]
  assign n8_I_190 = n7_O_190; // @[Top.scala 39:10]
  assign n8_I_191 = n7_O_191; // @[Top.scala 39:10]
  assign n8_I_192 = n7_O_192; // @[Top.scala 39:10]
  assign n8_I_193 = n7_O_193; // @[Top.scala 39:10]
  assign n8_I_194 = n7_O_194; // @[Top.scala 39:10]
  assign n8_I_195 = n7_O_195; // @[Top.scala 39:10]
  assign n8_I_196 = n7_O_196; // @[Top.scala 39:10]
  assign n8_I_197 = n7_O_197; // @[Top.scala 39:10]
  assign n8_I_198 = n7_O_198; // @[Top.scala 39:10]
  assign n8_I_199 = n7_O_199; // @[Top.scala 39:10]
  assign n9_clock = clock;
  assign n9_reset = reset;
  assign n9_valid_up = n8_valid_down; // @[Top.scala 43:17]
  assign n9_I_0 = n8_O_0; // @[Top.scala 42:10]
  assign n9_I_1 = n8_O_1; // @[Top.scala 42:10]
  assign n9_I_2 = n8_O_2; // @[Top.scala 42:10]
  assign n9_I_3 = n8_O_3; // @[Top.scala 42:10]
  assign n9_I_4 = n8_O_4; // @[Top.scala 42:10]
  assign n9_I_5 = n8_O_5; // @[Top.scala 42:10]
  assign n9_I_6 = n8_O_6; // @[Top.scala 42:10]
  assign n9_I_7 = n8_O_7; // @[Top.scala 42:10]
  assign n9_I_8 = n8_O_8; // @[Top.scala 42:10]
  assign n9_I_9 = n8_O_9; // @[Top.scala 42:10]
  assign n9_I_10 = n8_O_10; // @[Top.scala 42:10]
  assign n9_I_11 = n8_O_11; // @[Top.scala 42:10]
  assign n9_I_12 = n8_O_12; // @[Top.scala 42:10]
  assign n9_I_13 = n8_O_13; // @[Top.scala 42:10]
  assign n9_I_14 = n8_O_14; // @[Top.scala 42:10]
  assign n9_I_15 = n8_O_15; // @[Top.scala 42:10]
  assign n9_I_16 = n8_O_16; // @[Top.scala 42:10]
  assign n9_I_17 = n8_O_17; // @[Top.scala 42:10]
  assign n9_I_18 = n8_O_18; // @[Top.scala 42:10]
  assign n9_I_19 = n8_O_19; // @[Top.scala 42:10]
  assign n9_I_20 = n8_O_20; // @[Top.scala 42:10]
  assign n9_I_21 = n8_O_21; // @[Top.scala 42:10]
  assign n9_I_22 = n8_O_22; // @[Top.scala 42:10]
  assign n9_I_23 = n8_O_23; // @[Top.scala 42:10]
  assign n9_I_24 = n8_O_24; // @[Top.scala 42:10]
  assign n9_I_25 = n8_O_25; // @[Top.scala 42:10]
  assign n9_I_26 = n8_O_26; // @[Top.scala 42:10]
  assign n9_I_27 = n8_O_27; // @[Top.scala 42:10]
  assign n9_I_28 = n8_O_28; // @[Top.scala 42:10]
  assign n9_I_29 = n8_O_29; // @[Top.scala 42:10]
  assign n9_I_30 = n8_O_30; // @[Top.scala 42:10]
  assign n9_I_31 = n8_O_31; // @[Top.scala 42:10]
  assign n9_I_32 = n8_O_32; // @[Top.scala 42:10]
  assign n9_I_33 = n8_O_33; // @[Top.scala 42:10]
  assign n9_I_34 = n8_O_34; // @[Top.scala 42:10]
  assign n9_I_35 = n8_O_35; // @[Top.scala 42:10]
  assign n9_I_36 = n8_O_36; // @[Top.scala 42:10]
  assign n9_I_37 = n8_O_37; // @[Top.scala 42:10]
  assign n9_I_38 = n8_O_38; // @[Top.scala 42:10]
  assign n9_I_39 = n8_O_39; // @[Top.scala 42:10]
  assign n9_I_40 = n8_O_40; // @[Top.scala 42:10]
  assign n9_I_41 = n8_O_41; // @[Top.scala 42:10]
  assign n9_I_42 = n8_O_42; // @[Top.scala 42:10]
  assign n9_I_43 = n8_O_43; // @[Top.scala 42:10]
  assign n9_I_44 = n8_O_44; // @[Top.scala 42:10]
  assign n9_I_45 = n8_O_45; // @[Top.scala 42:10]
  assign n9_I_46 = n8_O_46; // @[Top.scala 42:10]
  assign n9_I_47 = n8_O_47; // @[Top.scala 42:10]
  assign n9_I_48 = n8_O_48; // @[Top.scala 42:10]
  assign n9_I_49 = n8_O_49; // @[Top.scala 42:10]
  assign n9_I_50 = n8_O_50; // @[Top.scala 42:10]
  assign n9_I_51 = n8_O_51; // @[Top.scala 42:10]
  assign n9_I_52 = n8_O_52; // @[Top.scala 42:10]
  assign n9_I_53 = n8_O_53; // @[Top.scala 42:10]
  assign n9_I_54 = n8_O_54; // @[Top.scala 42:10]
  assign n9_I_55 = n8_O_55; // @[Top.scala 42:10]
  assign n9_I_56 = n8_O_56; // @[Top.scala 42:10]
  assign n9_I_57 = n8_O_57; // @[Top.scala 42:10]
  assign n9_I_58 = n8_O_58; // @[Top.scala 42:10]
  assign n9_I_59 = n8_O_59; // @[Top.scala 42:10]
  assign n9_I_60 = n8_O_60; // @[Top.scala 42:10]
  assign n9_I_61 = n8_O_61; // @[Top.scala 42:10]
  assign n9_I_62 = n8_O_62; // @[Top.scala 42:10]
  assign n9_I_63 = n8_O_63; // @[Top.scala 42:10]
  assign n9_I_64 = n8_O_64; // @[Top.scala 42:10]
  assign n9_I_65 = n8_O_65; // @[Top.scala 42:10]
  assign n9_I_66 = n8_O_66; // @[Top.scala 42:10]
  assign n9_I_67 = n8_O_67; // @[Top.scala 42:10]
  assign n9_I_68 = n8_O_68; // @[Top.scala 42:10]
  assign n9_I_69 = n8_O_69; // @[Top.scala 42:10]
  assign n9_I_70 = n8_O_70; // @[Top.scala 42:10]
  assign n9_I_71 = n8_O_71; // @[Top.scala 42:10]
  assign n9_I_72 = n8_O_72; // @[Top.scala 42:10]
  assign n9_I_73 = n8_O_73; // @[Top.scala 42:10]
  assign n9_I_74 = n8_O_74; // @[Top.scala 42:10]
  assign n9_I_75 = n8_O_75; // @[Top.scala 42:10]
  assign n9_I_76 = n8_O_76; // @[Top.scala 42:10]
  assign n9_I_77 = n8_O_77; // @[Top.scala 42:10]
  assign n9_I_78 = n8_O_78; // @[Top.scala 42:10]
  assign n9_I_79 = n8_O_79; // @[Top.scala 42:10]
  assign n9_I_80 = n8_O_80; // @[Top.scala 42:10]
  assign n9_I_81 = n8_O_81; // @[Top.scala 42:10]
  assign n9_I_82 = n8_O_82; // @[Top.scala 42:10]
  assign n9_I_83 = n8_O_83; // @[Top.scala 42:10]
  assign n9_I_84 = n8_O_84; // @[Top.scala 42:10]
  assign n9_I_85 = n8_O_85; // @[Top.scala 42:10]
  assign n9_I_86 = n8_O_86; // @[Top.scala 42:10]
  assign n9_I_87 = n8_O_87; // @[Top.scala 42:10]
  assign n9_I_88 = n8_O_88; // @[Top.scala 42:10]
  assign n9_I_89 = n8_O_89; // @[Top.scala 42:10]
  assign n9_I_90 = n8_O_90; // @[Top.scala 42:10]
  assign n9_I_91 = n8_O_91; // @[Top.scala 42:10]
  assign n9_I_92 = n8_O_92; // @[Top.scala 42:10]
  assign n9_I_93 = n8_O_93; // @[Top.scala 42:10]
  assign n9_I_94 = n8_O_94; // @[Top.scala 42:10]
  assign n9_I_95 = n8_O_95; // @[Top.scala 42:10]
  assign n9_I_96 = n8_O_96; // @[Top.scala 42:10]
  assign n9_I_97 = n8_O_97; // @[Top.scala 42:10]
  assign n9_I_98 = n8_O_98; // @[Top.scala 42:10]
  assign n9_I_99 = n8_O_99; // @[Top.scala 42:10]
  assign n9_I_100 = n8_O_100; // @[Top.scala 42:10]
  assign n9_I_101 = n8_O_101; // @[Top.scala 42:10]
  assign n9_I_102 = n8_O_102; // @[Top.scala 42:10]
  assign n9_I_103 = n8_O_103; // @[Top.scala 42:10]
  assign n9_I_104 = n8_O_104; // @[Top.scala 42:10]
  assign n9_I_105 = n8_O_105; // @[Top.scala 42:10]
  assign n9_I_106 = n8_O_106; // @[Top.scala 42:10]
  assign n9_I_107 = n8_O_107; // @[Top.scala 42:10]
  assign n9_I_108 = n8_O_108; // @[Top.scala 42:10]
  assign n9_I_109 = n8_O_109; // @[Top.scala 42:10]
  assign n9_I_110 = n8_O_110; // @[Top.scala 42:10]
  assign n9_I_111 = n8_O_111; // @[Top.scala 42:10]
  assign n9_I_112 = n8_O_112; // @[Top.scala 42:10]
  assign n9_I_113 = n8_O_113; // @[Top.scala 42:10]
  assign n9_I_114 = n8_O_114; // @[Top.scala 42:10]
  assign n9_I_115 = n8_O_115; // @[Top.scala 42:10]
  assign n9_I_116 = n8_O_116; // @[Top.scala 42:10]
  assign n9_I_117 = n8_O_117; // @[Top.scala 42:10]
  assign n9_I_118 = n8_O_118; // @[Top.scala 42:10]
  assign n9_I_119 = n8_O_119; // @[Top.scala 42:10]
  assign n9_I_120 = n8_O_120; // @[Top.scala 42:10]
  assign n9_I_121 = n8_O_121; // @[Top.scala 42:10]
  assign n9_I_122 = n8_O_122; // @[Top.scala 42:10]
  assign n9_I_123 = n8_O_123; // @[Top.scala 42:10]
  assign n9_I_124 = n8_O_124; // @[Top.scala 42:10]
  assign n9_I_125 = n8_O_125; // @[Top.scala 42:10]
  assign n9_I_126 = n8_O_126; // @[Top.scala 42:10]
  assign n9_I_127 = n8_O_127; // @[Top.scala 42:10]
  assign n9_I_128 = n8_O_128; // @[Top.scala 42:10]
  assign n9_I_129 = n8_O_129; // @[Top.scala 42:10]
  assign n9_I_130 = n8_O_130; // @[Top.scala 42:10]
  assign n9_I_131 = n8_O_131; // @[Top.scala 42:10]
  assign n9_I_132 = n8_O_132; // @[Top.scala 42:10]
  assign n9_I_133 = n8_O_133; // @[Top.scala 42:10]
  assign n9_I_134 = n8_O_134; // @[Top.scala 42:10]
  assign n9_I_135 = n8_O_135; // @[Top.scala 42:10]
  assign n9_I_136 = n8_O_136; // @[Top.scala 42:10]
  assign n9_I_137 = n8_O_137; // @[Top.scala 42:10]
  assign n9_I_138 = n8_O_138; // @[Top.scala 42:10]
  assign n9_I_139 = n8_O_139; // @[Top.scala 42:10]
  assign n9_I_140 = n8_O_140; // @[Top.scala 42:10]
  assign n9_I_141 = n8_O_141; // @[Top.scala 42:10]
  assign n9_I_142 = n8_O_142; // @[Top.scala 42:10]
  assign n9_I_143 = n8_O_143; // @[Top.scala 42:10]
  assign n9_I_144 = n8_O_144; // @[Top.scala 42:10]
  assign n9_I_145 = n8_O_145; // @[Top.scala 42:10]
  assign n9_I_146 = n8_O_146; // @[Top.scala 42:10]
  assign n9_I_147 = n8_O_147; // @[Top.scala 42:10]
  assign n9_I_148 = n8_O_148; // @[Top.scala 42:10]
  assign n9_I_149 = n8_O_149; // @[Top.scala 42:10]
  assign n9_I_150 = n8_O_150; // @[Top.scala 42:10]
  assign n9_I_151 = n8_O_151; // @[Top.scala 42:10]
  assign n9_I_152 = n8_O_152; // @[Top.scala 42:10]
  assign n9_I_153 = n8_O_153; // @[Top.scala 42:10]
  assign n9_I_154 = n8_O_154; // @[Top.scala 42:10]
  assign n9_I_155 = n8_O_155; // @[Top.scala 42:10]
  assign n9_I_156 = n8_O_156; // @[Top.scala 42:10]
  assign n9_I_157 = n8_O_157; // @[Top.scala 42:10]
  assign n9_I_158 = n8_O_158; // @[Top.scala 42:10]
  assign n9_I_159 = n8_O_159; // @[Top.scala 42:10]
  assign n9_I_160 = n8_O_160; // @[Top.scala 42:10]
  assign n9_I_161 = n8_O_161; // @[Top.scala 42:10]
  assign n9_I_162 = n8_O_162; // @[Top.scala 42:10]
  assign n9_I_163 = n8_O_163; // @[Top.scala 42:10]
  assign n9_I_164 = n8_O_164; // @[Top.scala 42:10]
  assign n9_I_165 = n8_O_165; // @[Top.scala 42:10]
  assign n9_I_166 = n8_O_166; // @[Top.scala 42:10]
  assign n9_I_167 = n8_O_167; // @[Top.scala 42:10]
  assign n9_I_168 = n8_O_168; // @[Top.scala 42:10]
  assign n9_I_169 = n8_O_169; // @[Top.scala 42:10]
  assign n9_I_170 = n8_O_170; // @[Top.scala 42:10]
  assign n9_I_171 = n8_O_171; // @[Top.scala 42:10]
  assign n9_I_172 = n8_O_172; // @[Top.scala 42:10]
  assign n9_I_173 = n8_O_173; // @[Top.scala 42:10]
  assign n9_I_174 = n8_O_174; // @[Top.scala 42:10]
  assign n9_I_175 = n8_O_175; // @[Top.scala 42:10]
  assign n9_I_176 = n8_O_176; // @[Top.scala 42:10]
  assign n9_I_177 = n8_O_177; // @[Top.scala 42:10]
  assign n9_I_178 = n8_O_178; // @[Top.scala 42:10]
  assign n9_I_179 = n8_O_179; // @[Top.scala 42:10]
  assign n9_I_180 = n8_O_180; // @[Top.scala 42:10]
  assign n9_I_181 = n8_O_181; // @[Top.scala 42:10]
  assign n9_I_182 = n8_O_182; // @[Top.scala 42:10]
  assign n9_I_183 = n8_O_183; // @[Top.scala 42:10]
  assign n9_I_184 = n8_O_184; // @[Top.scala 42:10]
  assign n9_I_185 = n8_O_185; // @[Top.scala 42:10]
  assign n9_I_186 = n8_O_186; // @[Top.scala 42:10]
  assign n9_I_187 = n8_O_187; // @[Top.scala 42:10]
  assign n9_I_188 = n8_O_188; // @[Top.scala 42:10]
  assign n9_I_189 = n8_O_189; // @[Top.scala 42:10]
  assign n9_I_190 = n8_O_190; // @[Top.scala 42:10]
  assign n9_I_191 = n8_O_191; // @[Top.scala 42:10]
  assign n9_I_192 = n8_O_192; // @[Top.scala 42:10]
  assign n9_I_193 = n8_O_193; // @[Top.scala 42:10]
  assign n9_I_194 = n8_O_194; // @[Top.scala 42:10]
  assign n9_I_195 = n8_O_195; // @[Top.scala 42:10]
  assign n9_I_196 = n8_O_196; // @[Top.scala 42:10]
  assign n9_I_197 = n8_O_197; // @[Top.scala 42:10]
  assign n9_I_198 = n8_O_198; // @[Top.scala 42:10]
  assign n9_I_199 = n8_O_199; // @[Top.scala 42:10]
  assign n10_clock = clock;
  assign n10_reset = reset;
  assign n10_valid_up = n9_valid_down; // @[Top.scala 46:18]
  assign n10_I_0 = n9_O_0; // @[Top.scala 45:11]
  assign n10_I_1 = n9_O_1; // @[Top.scala 45:11]
  assign n10_I_2 = n9_O_2; // @[Top.scala 45:11]
  assign n10_I_3 = n9_O_3; // @[Top.scala 45:11]
  assign n10_I_4 = n9_O_4; // @[Top.scala 45:11]
  assign n10_I_5 = n9_O_5; // @[Top.scala 45:11]
  assign n10_I_6 = n9_O_6; // @[Top.scala 45:11]
  assign n10_I_7 = n9_O_7; // @[Top.scala 45:11]
  assign n10_I_8 = n9_O_8; // @[Top.scala 45:11]
  assign n10_I_9 = n9_O_9; // @[Top.scala 45:11]
  assign n10_I_10 = n9_O_10; // @[Top.scala 45:11]
  assign n10_I_11 = n9_O_11; // @[Top.scala 45:11]
  assign n10_I_12 = n9_O_12; // @[Top.scala 45:11]
  assign n10_I_13 = n9_O_13; // @[Top.scala 45:11]
  assign n10_I_14 = n9_O_14; // @[Top.scala 45:11]
  assign n10_I_15 = n9_O_15; // @[Top.scala 45:11]
  assign n10_I_16 = n9_O_16; // @[Top.scala 45:11]
  assign n10_I_17 = n9_O_17; // @[Top.scala 45:11]
  assign n10_I_18 = n9_O_18; // @[Top.scala 45:11]
  assign n10_I_19 = n9_O_19; // @[Top.scala 45:11]
  assign n10_I_20 = n9_O_20; // @[Top.scala 45:11]
  assign n10_I_21 = n9_O_21; // @[Top.scala 45:11]
  assign n10_I_22 = n9_O_22; // @[Top.scala 45:11]
  assign n10_I_23 = n9_O_23; // @[Top.scala 45:11]
  assign n10_I_24 = n9_O_24; // @[Top.scala 45:11]
  assign n10_I_25 = n9_O_25; // @[Top.scala 45:11]
  assign n10_I_26 = n9_O_26; // @[Top.scala 45:11]
  assign n10_I_27 = n9_O_27; // @[Top.scala 45:11]
  assign n10_I_28 = n9_O_28; // @[Top.scala 45:11]
  assign n10_I_29 = n9_O_29; // @[Top.scala 45:11]
  assign n10_I_30 = n9_O_30; // @[Top.scala 45:11]
  assign n10_I_31 = n9_O_31; // @[Top.scala 45:11]
  assign n10_I_32 = n9_O_32; // @[Top.scala 45:11]
  assign n10_I_33 = n9_O_33; // @[Top.scala 45:11]
  assign n10_I_34 = n9_O_34; // @[Top.scala 45:11]
  assign n10_I_35 = n9_O_35; // @[Top.scala 45:11]
  assign n10_I_36 = n9_O_36; // @[Top.scala 45:11]
  assign n10_I_37 = n9_O_37; // @[Top.scala 45:11]
  assign n10_I_38 = n9_O_38; // @[Top.scala 45:11]
  assign n10_I_39 = n9_O_39; // @[Top.scala 45:11]
  assign n10_I_40 = n9_O_40; // @[Top.scala 45:11]
  assign n10_I_41 = n9_O_41; // @[Top.scala 45:11]
  assign n10_I_42 = n9_O_42; // @[Top.scala 45:11]
  assign n10_I_43 = n9_O_43; // @[Top.scala 45:11]
  assign n10_I_44 = n9_O_44; // @[Top.scala 45:11]
  assign n10_I_45 = n9_O_45; // @[Top.scala 45:11]
  assign n10_I_46 = n9_O_46; // @[Top.scala 45:11]
  assign n10_I_47 = n9_O_47; // @[Top.scala 45:11]
  assign n10_I_48 = n9_O_48; // @[Top.scala 45:11]
  assign n10_I_49 = n9_O_49; // @[Top.scala 45:11]
  assign n10_I_50 = n9_O_50; // @[Top.scala 45:11]
  assign n10_I_51 = n9_O_51; // @[Top.scala 45:11]
  assign n10_I_52 = n9_O_52; // @[Top.scala 45:11]
  assign n10_I_53 = n9_O_53; // @[Top.scala 45:11]
  assign n10_I_54 = n9_O_54; // @[Top.scala 45:11]
  assign n10_I_55 = n9_O_55; // @[Top.scala 45:11]
  assign n10_I_56 = n9_O_56; // @[Top.scala 45:11]
  assign n10_I_57 = n9_O_57; // @[Top.scala 45:11]
  assign n10_I_58 = n9_O_58; // @[Top.scala 45:11]
  assign n10_I_59 = n9_O_59; // @[Top.scala 45:11]
  assign n10_I_60 = n9_O_60; // @[Top.scala 45:11]
  assign n10_I_61 = n9_O_61; // @[Top.scala 45:11]
  assign n10_I_62 = n9_O_62; // @[Top.scala 45:11]
  assign n10_I_63 = n9_O_63; // @[Top.scala 45:11]
  assign n10_I_64 = n9_O_64; // @[Top.scala 45:11]
  assign n10_I_65 = n9_O_65; // @[Top.scala 45:11]
  assign n10_I_66 = n9_O_66; // @[Top.scala 45:11]
  assign n10_I_67 = n9_O_67; // @[Top.scala 45:11]
  assign n10_I_68 = n9_O_68; // @[Top.scala 45:11]
  assign n10_I_69 = n9_O_69; // @[Top.scala 45:11]
  assign n10_I_70 = n9_O_70; // @[Top.scala 45:11]
  assign n10_I_71 = n9_O_71; // @[Top.scala 45:11]
  assign n10_I_72 = n9_O_72; // @[Top.scala 45:11]
  assign n10_I_73 = n9_O_73; // @[Top.scala 45:11]
  assign n10_I_74 = n9_O_74; // @[Top.scala 45:11]
  assign n10_I_75 = n9_O_75; // @[Top.scala 45:11]
  assign n10_I_76 = n9_O_76; // @[Top.scala 45:11]
  assign n10_I_77 = n9_O_77; // @[Top.scala 45:11]
  assign n10_I_78 = n9_O_78; // @[Top.scala 45:11]
  assign n10_I_79 = n9_O_79; // @[Top.scala 45:11]
  assign n10_I_80 = n9_O_80; // @[Top.scala 45:11]
  assign n10_I_81 = n9_O_81; // @[Top.scala 45:11]
  assign n10_I_82 = n9_O_82; // @[Top.scala 45:11]
  assign n10_I_83 = n9_O_83; // @[Top.scala 45:11]
  assign n10_I_84 = n9_O_84; // @[Top.scala 45:11]
  assign n10_I_85 = n9_O_85; // @[Top.scala 45:11]
  assign n10_I_86 = n9_O_86; // @[Top.scala 45:11]
  assign n10_I_87 = n9_O_87; // @[Top.scala 45:11]
  assign n10_I_88 = n9_O_88; // @[Top.scala 45:11]
  assign n10_I_89 = n9_O_89; // @[Top.scala 45:11]
  assign n10_I_90 = n9_O_90; // @[Top.scala 45:11]
  assign n10_I_91 = n9_O_91; // @[Top.scala 45:11]
  assign n10_I_92 = n9_O_92; // @[Top.scala 45:11]
  assign n10_I_93 = n9_O_93; // @[Top.scala 45:11]
  assign n10_I_94 = n9_O_94; // @[Top.scala 45:11]
  assign n10_I_95 = n9_O_95; // @[Top.scala 45:11]
  assign n10_I_96 = n9_O_96; // @[Top.scala 45:11]
  assign n10_I_97 = n9_O_97; // @[Top.scala 45:11]
  assign n10_I_98 = n9_O_98; // @[Top.scala 45:11]
  assign n10_I_99 = n9_O_99; // @[Top.scala 45:11]
  assign n10_I_100 = n9_O_100; // @[Top.scala 45:11]
  assign n10_I_101 = n9_O_101; // @[Top.scala 45:11]
  assign n10_I_102 = n9_O_102; // @[Top.scala 45:11]
  assign n10_I_103 = n9_O_103; // @[Top.scala 45:11]
  assign n10_I_104 = n9_O_104; // @[Top.scala 45:11]
  assign n10_I_105 = n9_O_105; // @[Top.scala 45:11]
  assign n10_I_106 = n9_O_106; // @[Top.scala 45:11]
  assign n10_I_107 = n9_O_107; // @[Top.scala 45:11]
  assign n10_I_108 = n9_O_108; // @[Top.scala 45:11]
  assign n10_I_109 = n9_O_109; // @[Top.scala 45:11]
  assign n10_I_110 = n9_O_110; // @[Top.scala 45:11]
  assign n10_I_111 = n9_O_111; // @[Top.scala 45:11]
  assign n10_I_112 = n9_O_112; // @[Top.scala 45:11]
  assign n10_I_113 = n9_O_113; // @[Top.scala 45:11]
  assign n10_I_114 = n9_O_114; // @[Top.scala 45:11]
  assign n10_I_115 = n9_O_115; // @[Top.scala 45:11]
  assign n10_I_116 = n9_O_116; // @[Top.scala 45:11]
  assign n10_I_117 = n9_O_117; // @[Top.scala 45:11]
  assign n10_I_118 = n9_O_118; // @[Top.scala 45:11]
  assign n10_I_119 = n9_O_119; // @[Top.scala 45:11]
  assign n10_I_120 = n9_O_120; // @[Top.scala 45:11]
  assign n10_I_121 = n9_O_121; // @[Top.scala 45:11]
  assign n10_I_122 = n9_O_122; // @[Top.scala 45:11]
  assign n10_I_123 = n9_O_123; // @[Top.scala 45:11]
  assign n10_I_124 = n9_O_124; // @[Top.scala 45:11]
  assign n10_I_125 = n9_O_125; // @[Top.scala 45:11]
  assign n10_I_126 = n9_O_126; // @[Top.scala 45:11]
  assign n10_I_127 = n9_O_127; // @[Top.scala 45:11]
  assign n10_I_128 = n9_O_128; // @[Top.scala 45:11]
  assign n10_I_129 = n9_O_129; // @[Top.scala 45:11]
  assign n10_I_130 = n9_O_130; // @[Top.scala 45:11]
  assign n10_I_131 = n9_O_131; // @[Top.scala 45:11]
  assign n10_I_132 = n9_O_132; // @[Top.scala 45:11]
  assign n10_I_133 = n9_O_133; // @[Top.scala 45:11]
  assign n10_I_134 = n9_O_134; // @[Top.scala 45:11]
  assign n10_I_135 = n9_O_135; // @[Top.scala 45:11]
  assign n10_I_136 = n9_O_136; // @[Top.scala 45:11]
  assign n10_I_137 = n9_O_137; // @[Top.scala 45:11]
  assign n10_I_138 = n9_O_138; // @[Top.scala 45:11]
  assign n10_I_139 = n9_O_139; // @[Top.scala 45:11]
  assign n10_I_140 = n9_O_140; // @[Top.scala 45:11]
  assign n10_I_141 = n9_O_141; // @[Top.scala 45:11]
  assign n10_I_142 = n9_O_142; // @[Top.scala 45:11]
  assign n10_I_143 = n9_O_143; // @[Top.scala 45:11]
  assign n10_I_144 = n9_O_144; // @[Top.scala 45:11]
  assign n10_I_145 = n9_O_145; // @[Top.scala 45:11]
  assign n10_I_146 = n9_O_146; // @[Top.scala 45:11]
  assign n10_I_147 = n9_O_147; // @[Top.scala 45:11]
  assign n10_I_148 = n9_O_148; // @[Top.scala 45:11]
  assign n10_I_149 = n9_O_149; // @[Top.scala 45:11]
  assign n10_I_150 = n9_O_150; // @[Top.scala 45:11]
  assign n10_I_151 = n9_O_151; // @[Top.scala 45:11]
  assign n10_I_152 = n9_O_152; // @[Top.scala 45:11]
  assign n10_I_153 = n9_O_153; // @[Top.scala 45:11]
  assign n10_I_154 = n9_O_154; // @[Top.scala 45:11]
  assign n10_I_155 = n9_O_155; // @[Top.scala 45:11]
  assign n10_I_156 = n9_O_156; // @[Top.scala 45:11]
  assign n10_I_157 = n9_O_157; // @[Top.scala 45:11]
  assign n10_I_158 = n9_O_158; // @[Top.scala 45:11]
  assign n10_I_159 = n9_O_159; // @[Top.scala 45:11]
  assign n10_I_160 = n9_O_160; // @[Top.scala 45:11]
  assign n10_I_161 = n9_O_161; // @[Top.scala 45:11]
  assign n10_I_162 = n9_O_162; // @[Top.scala 45:11]
  assign n10_I_163 = n9_O_163; // @[Top.scala 45:11]
  assign n10_I_164 = n9_O_164; // @[Top.scala 45:11]
  assign n10_I_165 = n9_O_165; // @[Top.scala 45:11]
  assign n10_I_166 = n9_O_166; // @[Top.scala 45:11]
  assign n10_I_167 = n9_O_167; // @[Top.scala 45:11]
  assign n10_I_168 = n9_O_168; // @[Top.scala 45:11]
  assign n10_I_169 = n9_O_169; // @[Top.scala 45:11]
  assign n10_I_170 = n9_O_170; // @[Top.scala 45:11]
  assign n10_I_171 = n9_O_171; // @[Top.scala 45:11]
  assign n10_I_172 = n9_O_172; // @[Top.scala 45:11]
  assign n10_I_173 = n9_O_173; // @[Top.scala 45:11]
  assign n10_I_174 = n9_O_174; // @[Top.scala 45:11]
  assign n10_I_175 = n9_O_175; // @[Top.scala 45:11]
  assign n10_I_176 = n9_O_176; // @[Top.scala 45:11]
  assign n10_I_177 = n9_O_177; // @[Top.scala 45:11]
  assign n10_I_178 = n9_O_178; // @[Top.scala 45:11]
  assign n10_I_179 = n9_O_179; // @[Top.scala 45:11]
  assign n10_I_180 = n9_O_180; // @[Top.scala 45:11]
  assign n10_I_181 = n9_O_181; // @[Top.scala 45:11]
  assign n10_I_182 = n9_O_182; // @[Top.scala 45:11]
  assign n10_I_183 = n9_O_183; // @[Top.scala 45:11]
  assign n10_I_184 = n9_O_184; // @[Top.scala 45:11]
  assign n10_I_185 = n9_O_185; // @[Top.scala 45:11]
  assign n10_I_186 = n9_O_186; // @[Top.scala 45:11]
  assign n10_I_187 = n9_O_187; // @[Top.scala 45:11]
  assign n10_I_188 = n9_O_188; // @[Top.scala 45:11]
  assign n10_I_189 = n9_O_189; // @[Top.scala 45:11]
  assign n10_I_190 = n9_O_190; // @[Top.scala 45:11]
  assign n10_I_191 = n9_O_191; // @[Top.scala 45:11]
  assign n10_I_192 = n9_O_192; // @[Top.scala 45:11]
  assign n10_I_193 = n9_O_193; // @[Top.scala 45:11]
  assign n10_I_194 = n9_O_194; // @[Top.scala 45:11]
  assign n10_I_195 = n9_O_195; // @[Top.scala 45:11]
  assign n10_I_196 = n9_O_196; // @[Top.scala 45:11]
  assign n10_I_197 = n9_O_197; // @[Top.scala 45:11]
  assign n10_I_198 = n9_O_198; // @[Top.scala 45:11]
  assign n10_I_199 = n9_O_199; // @[Top.scala 45:11]
endmodule
