module FIFO(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  input  [7:0] I_4,
  input  [7:0] I_5,
  input  [7:0] I_6,
  input  [7:0] I_7,
  input  [7:0] I_8,
  input  [7:0] I_9,
  input  [7:0] I_10,
  input  [7:0] I_11,
  input  [7:0] I_12,
  input  [7:0] I_13,
  input  [7:0] I_14,
  input  [7:0] I_15,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15
);
  reg [7:0] _T__0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg [7:0] _T__1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_1;
  reg [7:0] _T__2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_2;
  reg [7:0] _T__3; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_3;
  reg [7:0] _T__4; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_4;
  reg [7:0] _T__5; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_5;
  reg [7:0] _T__6; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_6;
  reg [7:0] _T__7; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_7;
  reg [7:0] _T__8; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_8;
  reg [7:0] _T__9; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_9;
  reg [7:0] _T__10; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_10;
  reg [7:0] _T__11; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_11;
  reg [7:0] _T__12; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_12;
  reg [7:0] _T__13; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_13;
  reg [7:0] _T__14; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_14;
  reg [7:0] _T__15; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_15;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_16;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O_0 = _T__0; // @[FIFO.scala 14:7]
  assign O_1 = _T__1; // @[FIFO.scala 14:7]
  assign O_2 = _T__2; // @[FIFO.scala 14:7]
  assign O_3 = _T__3; // @[FIFO.scala 14:7]
  assign O_4 = _T__4; // @[FIFO.scala 14:7]
  assign O_5 = _T__5; // @[FIFO.scala 14:7]
  assign O_6 = _T__6; // @[FIFO.scala 14:7]
  assign O_7 = _T__7; // @[FIFO.scala 14:7]
  assign O_8 = _T__8; // @[FIFO.scala 14:7]
  assign O_9 = _T__9; // @[FIFO.scala 14:7]
  assign O_10 = _T__10; // @[FIFO.scala 14:7]
  assign O_11 = _T__11; // @[FIFO.scala 14:7]
  assign O_12 = _T__12; // @[FIFO.scala 14:7]
  assign O_13 = _T__13; // @[FIFO.scala 14:7]
  assign O_14 = _T__14; // @[FIFO.scala 14:7]
  assign O_15 = _T__15; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T__0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T__1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__3 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T__4 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T__5 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__6 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__7 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T__8 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T__9 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T__10 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T__11 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T__12 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T__13 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T__14 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T__15 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_1 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T__0 <= I_0;
    _T__1 <= I_1;
    _T__2 <= I_2;
    _T__3 <= I_3;
    _T__4 <= I_4;
    _T__5 <= I_5;
    _T__6 <= I_6;
    _T__7 <= I_7;
    _T__8 <= I_8;
    _T__9 <= I_9;
    _T__10 <= I_10;
    _T__11 <= I_11;
    _T__12 <= I_12;
    _T__13 <= I_13;
    _T__14 <= I_14;
    _T__15 <= I_15;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module ShiftS(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  input  [7:0] I_4,
  input  [7:0] I_5,
  input  [7:0] I_6,
  input  [7:0] I_7,
  input  [7:0] I_8,
  input  [7:0] I_9,
  input  [7:0] I_10,
  input  [7:0] I_11,
  input  [7:0] I_12,
  input  [7:0] I_13,
  input  [7:0] I_14,
  input  [7:0] I_15,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15
);
  assign valid_down = valid_up; // @[ShiftS.scala 24:14]
  assign O_0 = I_12; // @[ShiftS.scala 21:31]
  assign O_1 = I_13; // @[ShiftS.scala 21:31]
  assign O_2 = I_14; // @[ShiftS.scala 21:31]
  assign O_3 = I_15; // @[ShiftS.scala 21:31]
  assign O_4 = I_0; // @[ShiftS.scala 21:31]
  assign O_5 = I_1; // @[ShiftS.scala 21:31]
  assign O_6 = I_2; // @[ShiftS.scala 21:31]
  assign O_7 = I_3; // @[ShiftS.scala 21:31]
  assign O_8 = I_4; // @[ShiftS.scala 21:31]
  assign O_9 = I_5; // @[ShiftS.scala 21:31]
  assign O_10 = I_6; // @[ShiftS.scala 21:31]
  assign O_11 = I_7; // @[ShiftS.scala 21:31]
  assign O_12 = I_8; // @[ShiftS.scala 21:31]
  assign O_13 = I_9; // @[ShiftS.scala 21:31]
  assign O_14 = I_10; // @[ShiftS.scala 21:31]
  assign O_15 = I_11; // @[ShiftS.scala 21:31]
endmodule
module ShiftS_2(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  input  [7:0] I_4,
  input  [7:0] I_5,
  input  [7:0] I_6,
  input  [7:0] I_7,
  input  [7:0] I_8,
  input  [7:0] I_9,
  input  [7:0] I_10,
  input  [7:0] I_11,
  input  [7:0] I_12,
  input  [7:0] I_13,
  input  [7:0] I_14,
  input  [7:0] I_15,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15
);
  assign valid_down = valid_up; // @[ShiftS.scala 24:14]
  assign O_0 = I_15; // @[ShiftS.scala 21:31]
  assign O_1 = I_0; // @[ShiftS.scala 21:31]
  assign O_2 = I_1; // @[ShiftS.scala 21:31]
  assign O_3 = I_2; // @[ShiftS.scala 21:31]
  assign O_4 = I_3; // @[ShiftS.scala 21:31]
  assign O_5 = I_4; // @[ShiftS.scala 21:31]
  assign O_6 = I_5; // @[ShiftS.scala 21:31]
  assign O_7 = I_6; // @[ShiftS.scala 21:31]
  assign O_8 = I_7; // @[ShiftS.scala 21:31]
  assign O_9 = I_8; // @[ShiftS.scala 21:31]
  assign O_10 = I_9; // @[ShiftS.scala 21:31]
  assign O_11 = I_10; // @[ShiftS.scala 21:31]
  assign O_12 = I_11; // @[ShiftS.scala 21:31]
  assign O_13 = I_12; // @[ShiftS.scala 21:31]
  assign O_14 = I_13; // @[ShiftS.scala 21:31]
  assign O_15 = I_14; // @[ShiftS.scala 21:31]
endmodule
module SSeqTupleCreator(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  input  [7:0] I1,
  output [7:0] O_0,
  output [7:0] O_1
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0 = I0; // @[Tuple.scala 12:32]
  assign O_1 = I1; // @[Tuple.scala 13:32]
endmodule
module Map2S(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I0_2,
  input  [7:0] I0_3,
  input  [7:0] I0_4,
  input  [7:0] I0_5,
  input  [7:0] I0_6,
  input  [7:0] I0_7,
  input  [7:0] I0_8,
  input  [7:0] I0_9,
  input  [7:0] I0_10,
  input  [7:0] I0_11,
  input  [7:0] I0_12,
  input  [7:0] I0_13,
  input  [7:0] I0_14,
  input  [7:0] I0_15,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  input  [7:0] I1_3,
  input  [7:0] I1_4,
  input  [7:0] I1_5,
  input  [7:0] I1_6,
  input  [7:0] I1_7,
  input  [7:0] I1_8,
  input  [7:0] I1_9,
  input  [7:0] I1_10,
  input  [7:0] I1_11,
  input  [7:0] I1_12,
  input  [7:0] I1_13,
  input  [7:0] I1_14,
  input  [7:0] I1_15,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_3_0,
  output [7:0] O_3_1,
  output [7:0] O_4_0,
  output [7:0] O_4_1,
  output [7:0] O_5_0,
  output [7:0] O_5_1,
  output [7:0] O_6_0,
  output [7:0] O_6_1,
  output [7:0] O_7_0,
  output [7:0] O_7_1,
  output [7:0] O_8_0,
  output [7:0] O_8_1,
  output [7:0] O_9_0,
  output [7:0] O_9_1,
  output [7:0] O_10_0,
  output [7:0] O_10_1,
  output [7:0] O_11_0,
  output [7:0] O_11_1,
  output [7:0] O_12_0,
  output [7:0] O_12_1,
  output [7:0] O_13_0,
  output [7:0] O_13_1,
  output [7:0] O_14_0,
  output [7:0] O_14_1,
  output [7:0] O_15_0,
  output [7:0] O_15_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_1; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  SSeqTupleCreator fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1)
  );
  SSeqTupleCreator other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1)
  );
  SSeqTupleCreator other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1)
  );
  SSeqTupleCreator other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0(other_ops_2_I0),
    .I1(other_ops_2_I1),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1)
  );
  SSeqTupleCreator other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0(other_ops_3_I0),
    .I1(other_ops_3_I1),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1)
  );
  SSeqTupleCreator other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0(other_ops_4_I0),
    .I1(other_ops_4_I1),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1)
  );
  SSeqTupleCreator other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0(other_ops_5_I0),
    .I1(other_ops_5_I1),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1)
  );
  SSeqTupleCreator other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0(other_ops_6_I0),
    .I1(other_ops_6_I1),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1)
  );
  SSeqTupleCreator other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0(other_ops_7_I0),
    .I1(other_ops_7_I1),
    .O_0(other_ops_7_O_0),
    .O_1(other_ops_7_O_1)
  );
  SSeqTupleCreator other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0(other_ops_8_I0),
    .I1(other_ops_8_I1),
    .O_0(other_ops_8_O_0),
    .O_1(other_ops_8_O_1)
  );
  SSeqTupleCreator other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0(other_ops_9_I0),
    .I1(other_ops_9_I1),
    .O_0(other_ops_9_O_0),
    .O_1(other_ops_9_O_1)
  );
  SSeqTupleCreator other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0(other_ops_10_I0),
    .I1(other_ops_10_I1),
    .O_0(other_ops_10_O_0),
    .O_1(other_ops_10_O_1)
  );
  SSeqTupleCreator other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0(other_ops_11_I0),
    .I1(other_ops_11_I1),
    .O_0(other_ops_11_O_0),
    .O_1(other_ops_11_O_1)
  );
  SSeqTupleCreator other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0(other_ops_12_I0),
    .I1(other_ops_12_I1),
    .O_0(other_ops_12_O_0),
    .O_1(other_ops_12_O_1)
  );
  SSeqTupleCreator other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0(other_ops_13_I0),
    .I1(other_ops_13_I1),
    .O_0(other_ops_13_O_0),
    .O_1(other_ops_13_O_1)
  );
  SSeqTupleCreator other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0(other_ops_14_I0),
    .I1(other_ops_14_I1),
    .O_0(other_ops_14_O_0),
    .O_1(other_ops_14_O_1)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_1_0 = other_ops_0_O_0; // @[Map2S.scala 24:12]
  assign O_1_1 = other_ops_0_O_1; // @[Map2S.scala 24:12]
  assign O_2_0 = other_ops_1_O_0; // @[Map2S.scala 24:12]
  assign O_2_1 = other_ops_1_O_1; // @[Map2S.scala 24:12]
  assign O_3_0 = other_ops_2_O_0; // @[Map2S.scala 24:12]
  assign O_3_1 = other_ops_2_O_1; // @[Map2S.scala 24:12]
  assign O_4_0 = other_ops_3_O_0; // @[Map2S.scala 24:12]
  assign O_4_1 = other_ops_3_O_1; // @[Map2S.scala 24:12]
  assign O_5_0 = other_ops_4_O_0; // @[Map2S.scala 24:12]
  assign O_5_1 = other_ops_4_O_1; // @[Map2S.scala 24:12]
  assign O_6_0 = other_ops_5_O_0; // @[Map2S.scala 24:12]
  assign O_6_1 = other_ops_5_O_1; // @[Map2S.scala 24:12]
  assign O_7_0 = other_ops_6_O_0; // @[Map2S.scala 24:12]
  assign O_7_1 = other_ops_6_O_1; // @[Map2S.scala 24:12]
  assign O_8_0 = other_ops_7_O_0; // @[Map2S.scala 24:12]
  assign O_8_1 = other_ops_7_O_1; // @[Map2S.scala 24:12]
  assign O_9_0 = other_ops_8_O_0; // @[Map2S.scala 24:12]
  assign O_9_1 = other_ops_8_O_1; // @[Map2S.scala 24:12]
  assign O_10_0 = other_ops_9_O_0; // @[Map2S.scala 24:12]
  assign O_10_1 = other_ops_9_O_1; // @[Map2S.scala 24:12]
  assign O_11_0 = other_ops_10_O_0; // @[Map2S.scala 24:12]
  assign O_11_1 = other_ops_10_O_1; // @[Map2S.scala 24:12]
  assign O_12_0 = other_ops_11_O_0; // @[Map2S.scala 24:12]
  assign O_12_1 = other_ops_11_O_1; // @[Map2S.scala 24:12]
  assign O_13_0 = other_ops_12_O_0; // @[Map2S.scala 24:12]
  assign O_13_1 = other_ops_12_O_1; // @[Map2S.scala 24:12]
  assign O_14_0 = other_ops_13_O_0; // @[Map2S.scala 24:12]
  assign O_14_1 = other_ops_13_O_1; // @[Map2S.scala 24:12]
  assign O_15_0 = other_ops_14_O_0; // @[Map2S.scala 24:12]
  assign O_15_1 = other_ops_14_O_1; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0 = I0_3; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0 = I0_4; // @[Map2S.scala 22:43]
  assign other_ops_3_I1 = I1_4; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0 = I0_5; // @[Map2S.scala 22:43]
  assign other_ops_4_I1 = I1_5; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0 = I0_6; // @[Map2S.scala 22:43]
  assign other_ops_5_I1 = I1_6; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0 = I0_7; // @[Map2S.scala 22:43]
  assign other_ops_6_I1 = I1_7; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0 = I0_8; // @[Map2S.scala 22:43]
  assign other_ops_7_I1 = I1_8; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0 = I0_9; // @[Map2S.scala 22:43]
  assign other_ops_8_I1 = I1_9; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0 = I0_10; // @[Map2S.scala 22:43]
  assign other_ops_9_I1 = I1_10; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0 = I0_11; // @[Map2S.scala 22:43]
  assign other_ops_10_I1 = I1_11; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0 = I0_12; // @[Map2S.scala 22:43]
  assign other_ops_11_I1 = I1_12; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0 = I0_13; // @[Map2S.scala 22:43]
  assign other_ops_12_I1 = I1_13; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0 = I0_14; // @[Map2S.scala 22:43]
  assign other_ops_13_I1 = I1_14; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0 = I0_15; // @[Map2S.scala 22:43]
  assign other_ops_14_I1 = I1_15; // @[Map2S.scala 23:43]
endmodule
module SSeqTupleAppender(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I1,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0 = I0_0; // @[Tuple.scala 24:34]
  assign O_1 = I0_1; // @[Tuple.scala 24:34]
  assign O_2 = I1; // @[Tuple.scala 26:32]
endmodule
module Map2S_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_2_0,
  input  [7:0] I0_2_1,
  input  [7:0] I0_3_0,
  input  [7:0] I0_3_1,
  input  [7:0] I0_4_0,
  input  [7:0] I0_4_1,
  input  [7:0] I0_5_0,
  input  [7:0] I0_5_1,
  input  [7:0] I0_6_0,
  input  [7:0] I0_6_1,
  input  [7:0] I0_7_0,
  input  [7:0] I0_7_1,
  input  [7:0] I0_8_0,
  input  [7:0] I0_8_1,
  input  [7:0] I0_9_0,
  input  [7:0] I0_9_1,
  input  [7:0] I0_10_0,
  input  [7:0] I0_10_1,
  input  [7:0] I0_11_0,
  input  [7:0] I0_11_1,
  input  [7:0] I0_12_0,
  input  [7:0] I0_12_1,
  input  [7:0] I0_13_0,
  input  [7:0] I0_13_1,
  input  [7:0] I0_14_0,
  input  [7:0] I0_14_1,
  input  [7:0] I0_15_0,
  input  [7:0] I0_15_1,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  input  [7:0] I1_3,
  input  [7:0] I1_4,
  input  [7:0] I1_5,
  input  [7:0] I1_6,
  input  [7:0] I1_7,
  input  [7:0] I1_8,
  input  [7:0] I1_9,
  input  [7:0] I1_10,
  input  [7:0] I1_11,
  input  [7:0] I1_12,
  input  [7:0] I1_13,
  input  [7:0] I1_14,
  input  [7:0] I1_15,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2,
  output [7:0] O_3_0,
  output [7:0] O_3_1,
  output [7:0] O_3_2,
  output [7:0] O_4_0,
  output [7:0] O_4_1,
  output [7:0] O_4_2,
  output [7:0] O_5_0,
  output [7:0] O_5_1,
  output [7:0] O_5_2,
  output [7:0] O_6_0,
  output [7:0] O_6_1,
  output [7:0] O_6_2,
  output [7:0] O_7_0,
  output [7:0] O_7_1,
  output [7:0] O_7_2,
  output [7:0] O_8_0,
  output [7:0] O_8_1,
  output [7:0] O_8_2,
  output [7:0] O_9_0,
  output [7:0] O_9_1,
  output [7:0] O_9_2,
  output [7:0] O_10_0,
  output [7:0] O_10_1,
  output [7:0] O_10_2,
  output [7:0] O_11_0,
  output [7:0] O_11_1,
  output [7:0] O_11_2,
  output [7:0] O_12_0,
  output [7:0] O_12_1,
  output [7:0] O_12_2,
  output [7:0] O_13_0,
  output [7:0] O_13_1,
  output [7:0] O_13_2,
  output [7:0] O_14_0,
  output [7:0] O_14_1,
  output [7:0] O_14_2,
  output [7:0] O_15_0,
  output [7:0] O_15_1,
  output [7:0] O_15_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  SSeqTupleAppender fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  SSeqTupleAppender other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I1(other_ops_0_I1),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  SSeqTupleAppender other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I1(other_ops_1_I1),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  SSeqTupleAppender other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0(other_ops_2_I0_0),
    .I0_1(other_ops_2_I0_1),
    .I1(other_ops_2_I1),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1),
    .O_2(other_ops_2_O_2)
  );
  SSeqTupleAppender other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0(other_ops_3_I0_0),
    .I0_1(other_ops_3_I0_1),
    .I1(other_ops_3_I1),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1),
    .O_2(other_ops_3_O_2)
  );
  SSeqTupleAppender other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0(other_ops_4_I0_0),
    .I0_1(other_ops_4_I0_1),
    .I1(other_ops_4_I1),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1),
    .O_2(other_ops_4_O_2)
  );
  SSeqTupleAppender other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0(other_ops_5_I0_0),
    .I0_1(other_ops_5_I0_1),
    .I1(other_ops_5_I1),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1),
    .O_2(other_ops_5_O_2)
  );
  SSeqTupleAppender other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0(other_ops_6_I0_0),
    .I0_1(other_ops_6_I0_1),
    .I1(other_ops_6_I1),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1),
    .O_2(other_ops_6_O_2)
  );
  SSeqTupleAppender other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0(other_ops_7_I0_0),
    .I0_1(other_ops_7_I0_1),
    .I1(other_ops_7_I1),
    .O_0(other_ops_7_O_0),
    .O_1(other_ops_7_O_1),
    .O_2(other_ops_7_O_2)
  );
  SSeqTupleAppender other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0(other_ops_8_I0_0),
    .I0_1(other_ops_8_I0_1),
    .I1(other_ops_8_I1),
    .O_0(other_ops_8_O_0),
    .O_1(other_ops_8_O_1),
    .O_2(other_ops_8_O_2)
  );
  SSeqTupleAppender other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0(other_ops_9_I0_0),
    .I0_1(other_ops_9_I0_1),
    .I1(other_ops_9_I1),
    .O_0(other_ops_9_O_0),
    .O_1(other_ops_9_O_1),
    .O_2(other_ops_9_O_2)
  );
  SSeqTupleAppender other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0(other_ops_10_I0_0),
    .I0_1(other_ops_10_I0_1),
    .I1(other_ops_10_I1),
    .O_0(other_ops_10_O_0),
    .O_1(other_ops_10_O_1),
    .O_2(other_ops_10_O_2)
  );
  SSeqTupleAppender other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0(other_ops_11_I0_0),
    .I0_1(other_ops_11_I0_1),
    .I1(other_ops_11_I1),
    .O_0(other_ops_11_O_0),
    .O_1(other_ops_11_O_1),
    .O_2(other_ops_11_O_2)
  );
  SSeqTupleAppender other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0(other_ops_12_I0_0),
    .I0_1(other_ops_12_I0_1),
    .I1(other_ops_12_I1),
    .O_0(other_ops_12_O_0),
    .O_1(other_ops_12_O_1),
    .O_2(other_ops_12_O_2)
  );
  SSeqTupleAppender other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0(other_ops_13_I0_0),
    .I0_1(other_ops_13_I0_1),
    .I1(other_ops_13_I1),
    .O_0(other_ops_13_O_0),
    .O_1(other_ops_13_O_1),
    .O_2(other_ops_13_O_2)
  );
  SSeqTupleAppender other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0(other_ops_14_I0_0),
    .I0_1(other_ops_14_I0_1),
    .I1(other_ops_14_I1),
    .O_0(other_ops_14_O_0),
    .O_1(other_ops_14_O_1),
    .O_2(other_ops_14_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_0_2 = fst_op_O_2; // @[Map2S.scala 19:8]
  assign O_1_0 = other_ops_0_O_0; // @[Map2S.scala 24:12]
  assign O_1_1 = other_ops_0_O_1; // @[Map2S.scala 24:12]
  assign O_1_2 = other_ops_0_O_2; // @[Map2S.scala 24:12]
  assign O_2_0 = other_ops_1_O_0; // @[Map2S.scala 24:12]
  assign O_2_1 = other_ops_1_O_1; // @[Map2S.scala 24:12]
  assign O_2_2 = other_ops_1_O_2; // @[Map2S.scala 24:12]
  assign O_3_0 = other_ops_2_O_0; // @[Map2S.scala 24:12]
  assign O_3_1 = other_ops_2_O_1; // @[Map2S.scala 24:12]
  assign O_3_2 = other_ops_2_O_2; // @[Map2S.scala 24:12]
  assign O_4_0 = other_ops_3_O_0; // @[Map2S.scala 24:12]
  assign O_4_1 = other_ops_3_O_1; // @[Map2S.scala 24:12]
  assign O_4_2 = other_ops_3_O_2; // @[Map2S.scala 24:12]
  assign O_5_0 = other_ops_4_O_0; // @[Map2S.scala 24:12]
  assign O_5_1 = other_ops_4_O_1; // @[Map2S.scala 24:12]
  assign O_5_2 = other_ops_4_O_2; // @[Map2S.scala 24:12]
  assign O_6_0 = other_ops_5_O_0; // @[Map2S.scala 24:12]
  assign O_6_1 = other_ops_5_O_1; // @[Map2S.scala 24:12]
  assign O_6_2 = other_ops_5_O_2; // @[Map2S.scala 24:12]
  assign O_7_0 = other_ops_6_O_0; // @[Map2S.scala 24:12]
  assign O_7_1 = other_ops_6_O_1; // @[Map2S.scala 24:12]
  assign O_7_2 = other_ops_6_O_2; // @[Map2S.scala 24:12]
  assign O_8_0 = other_ops_7_O_0; // @[Map2S.scala 24:12]
  assign O_8_1 = other_ops_7_O_1; // @[Map2S.scala 24:12]
  assign O_8_2 = other_ops_7_O_2; // @[Map2S.scala 24:12]
  assign O_9_0 = other_ops_8_O_0; // @[Map2S.scala 24:12]
  assign O_9_1 = other_ops_8_O_1; // @[Map2S.scala 24:12]
  assign O_9_2 = other_ops_8_O_2; // @[Map2S.scala 24:12]
  assign O_10_0 = other_ops_9_O_0; // @[Map2S.scala 24:12]
  assign O_10_1 = other_ops_9_O_1; // @[Map2S.scala 24:12]
  assign O_10_2 = other_ops_9_O_2; // @[Map2S.scala 24:12]
  assign O_11_0 = other_ops_10_O_0; // @[Map2S.scala 24:12]
  assign O_11_1 = other_ops_10_O_1; // @[Map2S.scala 24:12]
  assign O_11_2 = other_ops_10_O_2; // @[Map2S.scala 24:12]
  assign O_12_0 = other_ops_11_O_0; // @[Map2S.scala 24:12]
  assign O_12_1 = other_ops_11_O_1; // @[Map2S.scala 24:12]
  assign O_12_2 = other_ops_11_O_2; // @[Map2S.scala 24:12]
  assign O_13_0 = other_ops_12_O_0; // @[Map2S.scala 24:12]
  assign O_13_1 = other_ops_12_O_1; // @[Map2S.scala 24:12]
  assign O_13_2 = other_ops_12_O_2; // @[Map2S.scala 24:12]
  assign O_14_0 = other_ops_13_O_0; // @[Map2S.scala 24:12]
  assign O_14_1 = other_ops_13_O_1; // @[Map2S.scala 24:12]
  assign O_14_2 = other_ops_13_O_2; // @[Map2S.scala 24:12]
  assign O_15_0 = other_ops_14_O_0; // @[Map2S.scala 24:12]
  assign O_15_1 = other_ops_14_O_1; // @[Map2S.scala 24:12]
  assign O_15_2 = other_ops_14_O_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0 = I0_3_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1 = I0_3_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0 = I0_4_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1 = I0_4_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I1 = I1_4; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0 = I0_5_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1 = I0_5_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I1 = I1_5; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0 = I0_6_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1 = I0_6_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I1 = I1_6; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0 = I0_7_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1 = I0_7_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I1 = I1_7; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0 = I0_8_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1 = I0_8_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I1 = I1_8; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0 = I0_9_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1 = I0_9_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I1 = I1_9; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0 = I0_10_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1 = I0_10_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I1 = I1_10; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0 = I0_11_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1 = I0_11_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I1 = I1_11; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0 = I0_12_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1 = I0_12_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I1 = I1_12; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0 = I0_13_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1 = I0_13_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I1 = I1_13; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0 = I0_14_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1 = I0_14_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I1 = I1_14; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0 = I0_15_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1 = I0_15_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I1 = I1_15; // @[Map2S.scala 23:43]
endmodule
module PartitionS(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_2_2,
  input  [7:0] I_3_0,
  input  [7:0] I_3_1,
  input  [7:0] I_3_2,
  input  [7:0] I_4_0,
  input  [7:0] I_4_1,
  input  [7:0] I_4_2,
  input  [7:0] I_5_0,
  input  [7:0] I_5_1,
  input  [7:0] I_5_2,
  input  [7:0] I_6_0,
  input  [7:0] I_6_1,
  input  [7:0] I_6_2,
  input  [7:0] I_7_0,
  input  [7:0] I_7_1,
  input  [7:0] I_7_2,
  input  [7:0] I_8_0,
  input  [7:0] I_8_1,
  input  [7:0] I_8_2,
  input  [7:0] I_9_0,
  input  [7:0] I_9_1,
  input  [7:0] I_9_2,
  input  [7:0] I_10_0,
  input  [7:0] I_10_1,
  input  [7:0] I_10_2,
  input  [7:0] I_11_0,
  input  [7:0] I_11_1,
  input  [7:0] I_11_2,
  input  [7:0] I_12_0,
  input  [7:0] I_12_1,
  input  [7:0] I_12_2,
  input  [7:0] I_13_0,
  input  [7:0] I_13_1,
  input  [7:0] I_13_2,
  input  [7:0] I_14_0,
  input  [7:0] I_14_1,
  input  [7:0] I_14_2,
  input  [7:0] I_15_0,
  input  [7:0] I_15_1,
  input  [7:0] I_15_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_0_2,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_0_2,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_0_2,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_0_2,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_0_2,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_0_2,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_0_2,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_0_2
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0 = I_0_0; // @[Partition.scala 15:39]
  assign O_0_0_1 = I_0_1; // @[Partition.scala 15:39]
  assign O_0_0_2 = I_0_2; // @[Partition.scala 15:39]
  assign O_1_0_0 = I_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1 = I_1_1; // @[Partition.scala 15:39]
  assign O_1_0_2 = I_1_2; // @[Partition.scala 15:39]
  assign O_2_0_0 = I_2_0; // @[Partition.scala 15:39]
  assign O_2_0_1 = I_2_1; // @[Partition.scala 15:39]
  assign O_2_0_2 = I_2_2; // @[Partition.scala 15:39]
  assign O_3_0_0 = I_3_0; // @[Partition.scala 15:39]
  assign O_3_0_1 = I_3_1; // @[Partition.scala 15:39]
  assign O_3_0_2 = I_3_2; // @[Partition.scala 15:39]
  assign O_4_0_0 = I_4_0; // @[Partition.scala 15:39]
  assign O_4_0_1 = I_4_1; // @[Partition.scala 15:39]
  assign O_4_0_2 = I_4_2; // @[Partition.scala 15:39]
  assign O_5_0_0 = I_5_0; // @[Partition.scala 15:39]
  assign O_5_0_1 = I_5_1; // @[Partition.scala 15:39]
  assign O_5_0_2 = I_5_2; // @[Partition.scala 15:39]
  assign O_6_0_0 = I_6_0; // @[Partition.scala 15:39]
  assign O_6_0_1 = I_6_1; // @[Partition.scala 15:39]
  assign O_6_0_2 = I_6_2; // @[Partition.scala 15:39]
  assign O_7_0_0 = I_7_0; // @[Partition.scala 15:39]
  assign O_7_0_1 = I_7_1; // @[Partition.scala 15:39]
  assign O_7_0_2 = I_7_2; // @[Partition.scala 15:39]
  assign O_8_0_0 = I_8_0; // @[Partition.scala 15:39]
  assign O_8_0_1 = I_8_1; // @[Partition.scala 15:39]
  assign O_8_0_2 = I_8_2; // @[Partition.scala 15:39]
  assign O_9_0_0 = I_9_0; // @[Partition.scala 15:39]
  assign O_9_0_1 = I_9_1; // @[Partition.scala 15:39]
  assign O_9_0_2 = I_9_2; // @[Partition.scala 15:39]
  assign O_10_0_0 = I_10_0; // @[Partition.scala 15:39]
  assign O_10_0_1 = I_10_1; // @[Partition.scala 15:39]
  assign O_10_0_2 = I_10_2; // @[Partition.scala 15:39]
  assign O_11_0_0 = I_11_0; // @[Partition.scala 15:39]
  assign O_11_0_1 = I_11_1; // @[Partition.scala 15:39]
  assign O_11_0_2 = I_11_2; // @[Partition.scala 15:39]
  assign O_12_0_0 = I_12_0; // @[Partition.scala 15:39]
  assign O_12_0_1 = I_12_1; // @[Partition.scala 15:39]
  assign O_12_0_2 = I_12_2; // @[Partition.scala 15:39]
  assign O_13_0_0 = I_13_0; // @[Partition.scala 15:39]
  assign O_13_0_1 = I_13_1; // @[Partition.scala 15:39]
  assign O_13_0_2 = I_13_2; // @[Partition.scala 15:39]
  assign O_14_0_0 = I_14_0; // @[Partition.scala 15:39]
  assign O_14_0_1 = I_14_1; // @[Partition.scala 15:39]
  assign O_14_0_2 = I_14_2; // @[Partition.scala 15:39]
  assign O_15_0_0 = I_15_0; // @[Partition.scala 15:39]
  assign O_15_0_1 = I_15_1; // @[Partition.scala 15:39]
  assign O_15_0_2 = I_15_2; // @[Partition.scala 15:39]
endmodule
module SSeqTupleToSSeq(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0 = I_0; // @[Tuple.scala 41:5]
  assign O_1 = I_1; // @[Tuple.scala 41:5]
  assign O_2 = I_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0(op_inst_I_0),
    .I_1(op_inst_I_1),
    .I_2(op_inst_I_2),
    .O_0(op_inst_O_0),
    .O_1(op_inst_O_1),
    .O_2(op_inst_O_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0 = op_inst_O_0; // @[Remove1S.scala 14:5]
  assign O_1 = op_inst_O_1; // @[Remove1S.scala 14:5]
  assign O_2 = op_inst_O_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0 = I_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1 = I_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2 = I_0_2; // @[Remove1S.scala 13:13]
endmodule
module MapS(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_2_0_2,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_3_0_2,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_4_0_2,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_5_0_2,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_6_0_2,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_7_0_2,
  input  [7:0] I_8_0_0,
  input  [7:0] I_8_0_1,
  input  [7:0] I_8_0_2,
  input  [7:0] I_9_0_0,
  input  [7:0] I_9_0_1,
  input  [7:0] I_9_0_2,
  input  [7:0] I_10_0_0,
  input  [7:0] I_10_0_1,
  input  [7:0] I_10_0_2,
  input  [7:0] I_11_0_0,
  input  [7:0] I_11_0_1,
  input  [7:0] I_11_0_2,
  input  [7:0] I_12_0_0,
  input  [7:0] I_12_0_1,
  input  [7:0] I_12_0_2,
  input  [7:0] I_13_0_0,
  input  [7:0] I_13_0_1,
  input  [7:0] I_13_0_2,
  input  [7:0] I_14_0_0,
  input  [7:0] I_14_0_1,
  input  [7:0] I_14_0_2,
  input  [7:0] I_15_0_0,
  input  [7:0] I_15_0_1,
  input  [7:0] I_15_0_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2,
  output [7:0] O_3_0,
  output [7:0] O_3_1,
  output [7:0] O_3_2,
  output [7:0] O_4_0,
  output [7:0] O_4_1,
  output [7:0] O_4_2,
  output [7:0] O_5_0,
  output [7:0] O_5_1,
  output [7:0] O_5_2,
  output [7:0] O_6_0,
  output [7:0] O_6_1,
  output [7:0] O_6_2,
  output [7:0] O_7_0,
  output [7:0] O_7_1,
  output [7:0] O_7_2,
  output [7:0] O_8_0,
  output [7:0] O_8_1,
  output [7:0] O_8_2,
  output [7:0] O_9_0,
  output [7:0] O_9_1,
  output [7:0] O_9_2,
  output [7:0] O_10_0,
  output [7:0] O_10_1,
  output [7:0] O_10_2,
  output [7:0] O_11_0,
  output [7:0] O_11_1,
  output [7:0] O_11_2,
  output [7:0] O_12_0,
  output [7:0] O_12_1,
  output [7:0] O_12_2,
  output [7:0] O_13_0,
  output [7:0] O_13_1,
  output [7:0] O_13_2,
  output [7:0] O_14_0,
  output [7:0] O_14_1,
  output [7:0] O_14_2,
  output [7:0] O_15_0,
  output [7:0] O_15_1,
  output [7:0] O_15_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_2; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_2; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_2; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_2; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_2; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_2; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_2; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_2; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_2; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_2; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_2; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_2; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  Remove1S fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  Remove1S other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  Remove1S other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_0_2(other_ops_1_I_0_2),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  Remove1S other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_0_2(other_ops_2_I_0_2),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1),
    .O_2(other_ops_2_O_2)
  );
  Remove1S other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0(other_ops_3_I_0_0),
    .I_0_1(other_ops_3_I_0_1),
    .I_0_2(other_ops_3_I_0_2),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1),
    .O_2(other_ops_3_O_2)
  );
  Remove1S other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0(other_ops_4_I_0_0),
    .I_0_1(other_ops_4_I_0_1),
    .I_0_2(other_ops_4_I_0_2),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1),
    .O_2(other_ops_4_O_2)
  );
  Remove1S other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0(other_ops_5_I_0_0),
    .I_0_1(other_ops_5_I_0_1),
    .I_0_2(other_ops_5_I_0_2),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1),
    .O_2(other_ops_5_O_2)
  );
  Remove1S other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0(other_ops_6_I_0_0),
    .I_0_1(other_ops_6_I_0_1),
    .I_0_2(other_ops_6_I_0_2),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1),
    .O_2(other_ops_6_O_2)
  );
  Remove1S other_ops_7 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I_0_0(other_ops_7_I_0_0),
    .I_0_1(other_ops_7_I_0_1),
    .I_0_2(other_ops_7_I_0_2),
    .O_0(other_ops_7_O_0),
    .O_1(other_ops_7_O_1),
    .O_2(other_ops_7_O_2)
  );
  Remove1S other_ops_8 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I_0_0(other_ops_8_I_0_0),
    .I_0_1(other_ops_8_I_0_1),
    .I_0_2(other_ops_8_I_0_2),
    .O_0(other_ops_8_O_0),
    .O_1(other_ops_8_O_1),
    .O_2(other_ops_8_O_2)
  );
  Remove1S other_ops_9 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I_0_0(other_ops_9_I_0_0),
    .I_0_1(other_ops_9_I_0_1),
    .I_0_2(other_ops_9_I_0_2),
    .O_0(other_ops_9_O_0),
    .O_1(other_ops_9_O_1),
    .O_2(other_ops_9_O_2)
  );
  Remove1S other_ops_10 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I_0_0(other_ops_10_I_0_0),
    .I_0_1(other_ops_10_I_0_1),
    .I_0_2(other_ops_10_I_0_2),
    .O_0(other_ops_10_O_0),
    .O_1(other_ops_10_O_1),
    .O_2(other_ops_10_O_2)
  );
  Remove1S other_ops_11 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I_0_0(other_ops_11_I_0_0),
    .I_0_1(other_ops_11_I_0_1),
    .I_0_2(other_ops_11_I_0_2),
    .O_0(other_ops_11_O_0),
    .O_1(other_ops_11_O_1),
    .O_2(other_ops_11_O_2)
  );
  Remove1S other_ops_12 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I_0_0(other_ops_12_I_0_0),
    .I_0_1(other_ops_12_I_0_1),
    .I_0_2(other_ops_12_I_0_2),
    .O_0(other_ops_12_O_0),
    .O_1(other_ops_12_O_1),
    .O_2(other_ops_12_O_2)
  );
  Remove1S other_ops_13 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I_0_0(other_ops_13_I_0_0),
    .I_0_1(other_ops_13_I_0_1),
    .I_0_2(other_ops_13_I_0_2),
    .O_0(other_ops_13_O_0),
    .O_1(other_ops_13_O_1),
    .O_2(other_ops_13_O_2)
  );
  Remove1S other_ops_14 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I_0_0(other_ops_14_I_0_0),
    .I_0_1(other_ops_14_I_0_1),
    .I_0_2(other_ops_14_I_0_2),
    .O_0(other_ops_14_O_0),
    .O_1(other_ops_14_O_1),
    .O_2(other_ops_14_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_1_2 = other_ops_0_O_2; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign O_2_1 = other_ops_1_O_1; // @[MapS.scala 21:12]
  assign O_2_2 = other_ops_1_O_2; // @[MapS.scala 21:12]
  assign O_3_0 = other_ops_2_O_0; // @[MapS.scala 21:12]
  assign O_3_1 = other_ops_2_O_1; // @[MapS.scala 21:12]
  assign O_3_2 = other_ops_2_O_2; // @[MapS.scala 21:12]
  assign O_4_0 = other_ops_3_O_0; // @[MapS.scala 21:12]
  assign O_4_1 = other_ops_3_O_1; // @[MapS.scala 21:12]
  assign O_4_2 = other_ops_3_O_2; // @[MapS.scala 21:12]
  assign O_5_0 = other_ops_4_O_0; // @[MapS.scala 21:12]
  assign O_5_1 = other_ops_4_O_1; // @[MapS.scala 21:12]
  assign O_5_2 = other_ops_4_O_2; // @[MapS.scala 21:12]
  assign O_6_0 = other_ops_5_O_0; // @[MapS.scala 21:12]
  assign O_6_1 = other_ops_5_O_1; // @[MapS.scala 21:12]
  assign O_6_2 = other_ops_5_O_2; // @[MapS.scala 21:12]
  assign O_7_0 = other_ops_6_O_0; // @[MapS.scala 21:12]
  assign O_7_1 = other_ops_6_O_1; // @[MapS.scala 21:12]
  assign O_7_2 = other_ops_6_O_2; // @[MapS.scala 21:12]
  assign O_8_0 = other_ops_7_O_0; // @[MapS.scala 21:12]
  assign O_8_1 = other_ops_7_O_1; // @[MapS.scala 21:12]
  assign O_8_2 = other_ops_7_O_2; // @[MapS.scala 21:12]
  assign O_9_0 = other_ops_8_O_0; // @[MapS.scala 21:12]
  assign O_9_1 = other_ops_8_O_1; // @[MapS.scala 21:12]
  assign O_9_2 = other_ops_8_O_2; // @[MapS.scala 21:12]
  assign O_10_0 = other_ops_9_O_0; // @[MapS.scala 21:12]
  assign O_10_1 = other_ops_9_O_1; // @[MapS.scala 21:12]
  assign O_10_2 = other_ops_9_O_2; // @[MapS.scala 21:12]
  assign O_11_0 = other_ops_10_O_0; // @[MapS.scala 21:12]
  assign O_11_1 = other_ops_10_O_1; // @[MapS.scala 21:12]
  assign O_11_2 = other_ops_10_O_2; // @[MapS.scala 21:12]
  assign O_12_0 = other_ops_11_O_0; // @[MapS.scala 21:12]
  assign O_12_1 = other_ops_11_O_1; // @[MapS.scala 21:12]
  assign O_12_2 = other_ops_11_O_2; // @[MapS.scala 21:12]
  assign O_13_0 = other_ops_12_O_0; // @[MapS.scala 21:12]
  assign O_13_1 = other_ops_12_O_1; // @[MapS.scala 21:12]
  assign O_13_2 = other_ops_12_O_2; // @[MapS.scala 21:12]
  assign O_14_0 = other_ops_13_O_0; // @[MapS.scala 21:12]
  assign O_14_1 = other_ops_13_O_1; // @[MapS.scala 21:12]
  assign O_14_2 = other_ops_13_O_2; // @[MapS.scala 21:12]
  assign O_15_0 = other_ops_14_O_0; // @[MapS.scala 21:12]
  assign O_15_1 = other_ops_14_O_1; // @[MapS.scala 21:12]
  assign O_15_2 = other_ops_14_O_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2 = I_2_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2 = I_3_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0 = I_4_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1 = I_4_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2 = I_4_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0 = I_5_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1 = I_5_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2 = I_5_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0 = I_6_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1 = I_6_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2 = I_6_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0 = I_7_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1 = I_7_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2 = I_7_0_2; // @[MapS.scala 20:41]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I_0_0 = I_8_0_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1 = I_8_0_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2 = I_8_0_2; // @[MapS.scala 20:41]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I_0_0 = I_9_0_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1 = I_9_0_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2 = I_9_0_2; // @[MapS.scala 20:41]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I_0_0 = I_10_0_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1 = I_10_0_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2 = I_10_0_2; // @[MapS.scala 20:41]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I_0_0 = I_11_0_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1 = I_11_0_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2 = I_11_0_2; // @[MapS.scala 20:41]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I_0_0 = I_12_0_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1 = I_12_0_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2 = I_12_0_2; // @[MapS.scala 20:41]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I_0_0 = I_13_0_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1 = I_13_0_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2 = I_13_0_2; // @[MapS.scala 20:41]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I_0_0 = I_14_0_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1 = I_14_0_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2 = I_14_0_2; // @[MapS.scala 20:41]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I_0_0 = I_15_0_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1 = I_15_0_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2 = I_15_0_2; // @[MapS.scala 20:41]
endmodule
module SSeqTupleCreator_2(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I0_2,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0_0 = I0_0; // @[Tuple.scala 12:32]
  assign O_0_1 = I0_1; // @[Tuple.scala 12:32]
  assign O_0_2 = I0_2; // @[Tuple.scala 12:32]
  assign O_1_0 = I1_0; // @[Tuple.scala 13:32]
  assign O_1_1 = I1_1; // @[Tuple.scala 13:32]
  assign O_1_2 = I1_2; // @[Tuple.scala 13:32]
endmodule
module Map2S_4(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_0_2,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_1_2,
  input  [7:0] I0_2_0,
  input  [7:0] I0_2_1,
  input  [7:0] I0_2_2,
  input  [7:0] I0_3_0,
  input  [7:0] I0_3_1,
  input  [7:0] I0_3_2,
  input  [7:0] I0_4_0,
  input  [7:0] I0_4_1,
  input  [7:0] I0_4_2,
  input  [7:0] I0_5_0,
  input  [7:0] I0_5_1,
  input  [7:0] I0_5_2,
  input  [7:0] I0_6_0,
  input  [7:0] I0_6_1,
  input  [7:0] I0_6_2,
  input  [7:0] I0_7_0,
  input  [7:0] I0_7_1,
  input  [7:0] I0_7_2,
  input  [7:0] I0_8_0,
  input  [7:0] I0_8_1,
  input  [7:0] I0_8_2,
  input  [7:0] I0_9_0,
  input  [7:0] I0_9_1,
  input  [7:0] I0_9_2,
  input  [7:0] I0_10_0,
  input  [7:0] I0_10_1,
  input  [7:0] I0_10_2,
  input  [7:0] I0_11_0,
  input  [7:0] I0_11_1,
  input  [7:0] I0_11_2,
  input  [7:0] I0_12_0,
  input  [7:0] I0_12_1,
  input  [7:0] I0_12_2,
  input  [7:0] I0_13_0,
  input  [7:0] I0_13_1,
  input  [7:0] I0_13_2,
  input  [7:0] I0_14_0,
  input  [7:0] I0_14_1,
  input  [7:0] I0_14_2,
  input  [7:0] I0_15_0,
  input  [7:0] I0_15_1,
  input  [7:0] I0_15_2,
  input  [7:0] I1_0_0,
  input  [7:0] I1_0_1,
  input  [7:0] I1_0_2,
  input  [7:0] I1_1_0,
  input  [7:0] I1_1_1,
  input  [7:0] I1_1_2,
  input  [7:0] I1_2_0,
  input  [7:0] I1_2_1,
  input  [7:0] I1_2_2,
  input  [7:0] I1_3_0,
  input  [7:0] I1_3_1,
  input  [7:0] I1_3_2,
  input  [7:0] I1_4_0,
  input  [7:0] I1_4_1,
  input  [7:0] I1_4_2,
  input  [7:0] I1_5_0,
  input  [7:0] I1_5_1,
  input  [7:0] I1_5_2,
  input  [7:0] I1_6_0,
  input  [7:0] I1_6_1,
  input  [7:0] I1_6_2,
  input  [7:0] I1_7_0,
  input  [7:0] I1_7_1,
  input  [7:0] I1_7_2,
  input  [7:0] I1_8_0,
  input  [7:0] I1_8_1,
  input  [7:0] I1_8_2,
  input  [7:0] I1_9_0,
  input  [7:0] I1_9_1,
  input  [7:0] I1_9_2,
  input  [7:0] I1_10_0,
  input  [7:0] I1_10_1,
  input  [7:0] I1_10_2,
  input  [7:0] I1_11_0,
  input  [7:0] I1_11_1,
  input  [7:0] I1_11_2,
  input  [7:0] I1_12_0,
  input  [7:0] I1_12_1,
  input  [7:0] I1_12_2,
  input  [7:0] I1_13_0,
  input  [7:0] I1_13_1,
  input  [7:0] I1_13_2,
  input  [7:0] I1_14_0,
  input  [7:0] I1_14_1,
  input  [7:0] I1_14_2,
  input  [7:0] I1_15_0,
  input  [7:0] I1_15_1,
  input  [7:0] I1_15_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_2_1_0,
  output [7:0] O_2_1_1,
  output [7:0] O_2_1_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_3_1_0,
  output [7:0] O_3_1_1,
  output [7:0] O_3_1_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_4_1_0,
  output [7:0] O_4_1_1,
  output [7:0] O_4_1_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_5_1_0,
  output [7:0] O_5_1_1,
  output [7:0] O_5_1_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_6_1_0,
  output [7:0] O_6_1_1,
  output [7:0] O_6_1_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2,
  output [7:0] O_7_1_0,
  output [7:0] O_7_1_1,
  output [7:0] O_7_1_2,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_0_2,
  output [7:0] O_8_1_0,
  output [7:0] O_8_1_1,
  output [7:0] O_8_1_2,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_0_2,
  output [7:0] O_9_1_0,
  output [7:0] O_9_1_1,
  output [7:0] O_9_1_2,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_0_2,
  output [7:0] O_10_1_0,
  output [7:0] O_10_1_1,
  output [7:0] O_10_1_2,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_0_2,
  output [7:0] O_11_1_0,
  output [7:0] O_11_1_1,
  output [7:0] O_11_1_2,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_0_2,
  output [7:0] O_12_1_0,
  output [7:0] O_12_1_1,
  output [7:0] O_12_1_2,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_0_2,
  output [7:0] O_13_1_0,
  output [7:0] O_13_1_1,
  output [7:0] O_13_1_2,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_0_2,
  output [7:0] O_14_1_0,
  output [7:0] O_14_1_1,
  output [7:0] O_14_1_2,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_0_2,
  output [7:0] O_15_1_0,
  output [7:0] O_15_1_1,
  output [7:0] O_15_1_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_1_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  SSeqTupleCreator_2 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I0_2(other_ops_0_I0_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I0_2(other_ops_1_I0_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0(other_ops_2_I0_0),
    .I0_1(other_ops_2_I0_1),
    .I0_2(other_ops_2_I0_2),
    .I1_0(other_ops_2_I1_0),
    .I1_1(other_ops_2_I1_1),
    .I1_2(other_ops_2_I1_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0(other_ops_3_I0_0),
    .I0_1(other_ops_3_I0_1),
    .I0_2(other_ops_3_I0_2),
    .I1_0(other_ops_3_I1_0),
    .I1_1(other_ops_3_I1_1),
    .I1_2(other_ops_3_I1_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0(other_ops_4_I0_0),
    .I0_1(other_ops_4_I0_1),
    .I0_2(other_ops_4_I0_2),
    .I1_0(other_ops_4_I1_0),
    .I1_1(other_ops_4_I1_1),
    .I1_2(other_ops_4_I1_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0(other_ops_5_I0_0),
    .I0_1(other_ops_5_I0_1),
    .I0_2(other_ops_5_I0_2),
    .I1_0(other_ops_5_I1_0),
    .I1_1(other_ops_5_I1_1),
    .I1_2(other_ops_5_I1_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0(other_ops_6_I0_0),
    .I0_1(other_ops_6_I0_1),
    .I0_2(other_ops_6_I0_2),
    .I1_0(other_ops_6_I1_0),
    .I1_1(other_ops_6_I1_1),
    .I1_2(other_ops_6_I1_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0(other_ops_7_I0_0),
    .I0_1(other_ops_7_I0_1),
    .I0_2(other_ops_7_I0_2),
    .I1_0(other_ops_7_I1_0),
    .I1_1(other_ops_7_I1_1),
    .I1_2(other_ops_7_I1_2),
    .O_0_0(other_ops_7_O_0_0),
    .O_0_1(other_ops_7_O_0_1),
    .O_0_2(other_ops_7_O_0_2),
    .O_1_0(other_ops_7_O_1_0),
    .O_1_1(other_ops_7_O_1_1),
    .O_1_2(other_ops_7_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0(other_ops_8_I0_0),
    .I0_1(other_ops_8_I0_1),
    .I0_2(other_ops_8_I0_2),
    .I1_0(other_ops_8_I1_0),
    .I1_1(other_ops_8_I1_1),
    .I1_2(other_ops_8_I1_2),
    .O_0_0(other_ops_8_O_0_0),
    .O_0_1(other_ops_8_O_0_1),
    .O_0_2(other_ops_8_O_0_2),
    .O_1_0(other_ops_8_O_1_0),
    .O_1_1(other_ops_8_O_1_1),
    .O_1_2(other_ops_8_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0(other_ops_9_I0_0),
    .I0_1(other_ops_9_I0_1),
    .I0_2(other_ops_9_I0_2),
    .I1_0(other_ops_9_I1_0),
    .I1_1(other_ops_9_I1_1),
    .I1_2(other_ops_9_I1_2),
    .O_0_0(other_ops_9_O_0_0),
    .O_0_1(other_ops_9_O_0_1),
    .O_0_2(other_ops_9_O_0_2),
    .O_1_0(other_ops_9_O_1_0),
    .O_1_1(other_ops_9_O_1_1),
    .O_1_2(other_ops_9_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0(other_ops_10_I0_0),
    .I0_1(other_ops_10_I0_1),
    .I0_2(other_ops_10_I0_2),
    .I1_0(other_ops_10_I1_0),
    .I1_1(other_ops_10_I1_1),
    .I1_2(other_ops_10_I1_2),
    .O_0_0(other_ops_10_O_0_0),
    .O_0_1(other_ops_10_O_0_1),
    .O_0_2(other_ops_10_O_0_2),
    .O_1_0(other_ops_10_O_1_0),
    .O_1_1(other_ops_10_O_1_1),
    .O_1_2(other_ops_10_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0(other_ops_11_I0_0),
    .I0_1(other_ops_11_I0_1),
    .I0_2(other_ops_11_I0_2),
    .I1_0(other_ops_11_I1_0),
    .I1_1(other_ops_11_I1_1),
    .I1_2(other_ops_11_I1_2),
    .O_0_0(other_ops_11_O_0_0),
    .O_0_1(other_ops_11_O_0_1),
    .O_0_2(other_ops_11_O_0_2),
    .O_1_0(other_ops_11_O_1_0),
    .O_1_1(other_ops_11_O_1_1),
    .O_1_2(other_ops_11_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0(other_ops_12_I0_0),
    .I0_1(other_ops_12_I0_1),
    .I0_2(other_ops_12_I0_2),
    .I1_0(other_ops_12_I1_0),
    .I1_1(other_ops_12_I1_1),
    .I1_2(other_ops_12_I1_2),
    .O_0_0(other_ops_12_O_0_0),
    .O_0_1(other_ops_12_O_0_1),
    .O_0_2(other_ops_12_O_0_2),
    .O_1_0(other_ops_12_O_1_0),
    .O_1_1(other_ops_12_O_1_1),
    .O_1_2(other_ops_12_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0(other_ops_13_I0_0),
    .I0_1(other_ops_13_I0_1),
    .I0_2(other_ops_13_I0_2),
    .I1_0(other_ops_13_I1_0),
    .I1_1(other_ops_13_I1_1),
    .I1_2(other_ops_13_I1_2),
    .O_0_0(other_ops_13_O_0_0),
    .O_0_1(other_ops_13_O_0_1),
    .O_0_2(other_ops_13_O_0_2),
    .O_1_0(other_ops_13_O_1_0),
    .O_1_1(other_ops_13_O_1_1),
    .O_1_2(other_ops_13_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0(other_ops_14_I0_0),
    .I0_1(other_ops_14_I0_1),
    .I0_2(other_ops_14_I0_2),
    .I1_0(other_ops_14_I1_0),
    .I1_1(other_ops_14_I1_1),
    .I1_2(other_ops_14_I1_2),
    .O_0_0(other_ops_14_O_0_0),
    .O_0_1(other_ops_14_O_0_1),
    .O_0_2(other_ops_14_O_0_2),
    .O_1_0(other_ops_14_O_1_0),
    .O_1_1(other_ops_14_O_1_1),
    .O_1_2(other_ops_14_O_1_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[Map2S.scala 24:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[Map2S.scala 24:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[Map2S.scala 24:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[Map2S.scala 24:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[Map2S.scala 24:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[Map2S.scala 24:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[Map2S.scala 24:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[Map2S.scala 24:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[Map2S.scala 24:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[Map2S.scala 24:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[Map2S.scala 24:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[Map2S.scala 24:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[Map2S.scala 24:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[Map2S.scala 24:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[Map2S.scala 24:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[Map2S.scala 24:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[Map2S.scala 24:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[Map2S.scala 24:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[Map2S.scala 24:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[Map2S.scala 24:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[Map2S.scala 24:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[Map2S.scala 24:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[Map2S.scala 24:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[Map2S.scala 24:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[Map2S.scala 24:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[Map2S.scala 24:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[Map2S.scala 24:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[Map2S.scala 24:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[Map2S.scala 24:12]
  assign O_8_0_1 = other_ops_7_O_0_1; // @[Map2S.scala 24:12]
  assign O_8_0_2 = other_ops_7_O_0_2; // @[Map2S.scala 24:12]
  assign O_8_1_0 = other_ops_7_O_1_0; // @[Map2S.scala 24:12]
  assign O_8_1_1 = other_ops_7_O_1_1; // @[Map2S.scala 24:12]
  assign O_8_1_2 = other_ops_7_O_1_2; // @[Map2S.scala 24:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[Map2S.scala 24:12]
  assign O_9_0_1 = other_ops_8_O_0_1; // @[Map2S.scala 24:12]
  assign O_9_0_2 = other_ops_8_O_0_2; // @[Map2S.scala 24:12]
  assign O_9_1_0 = other_ops_8_O_1_0; // @[Map2S.scala 24:12]
  assign O_9_1_1 = other_ops_8_O_1_1; // @[Map2S.scala 24:12]
  assign O_9_1_2 = other_ops_8_O_1_2; // @[Map2S.scala 24:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[Map2S.scala 24:12]
  assign O_10_0_1 = other_ops_9_O_0_1; // @[Map2S.scala 24:12]
  assign O_10_0_2 = other_ops_9_O_0_2; // @[Map2S.scala 24:12]
  assign O_10_1_0 = other_ops_9_O_1_0; // @[Map2S.scala 24:12]
  assign O_10_1_1 = other_ops_9_O_1_1; // @[Map2S.scala 24:12]
  assign O_10_1_2 = other_ops_9_O_1_2; // @[Map2S.scala 24:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[Map2S.scala 24:12]
  assign O_11_0_1 = other_ops_10_O_0_1; // @[Map2S.scala 24:12]
  assign O_11_0_2 = other_ops_10_O_0_2; // @[Map2S.scala 24:12]
  assign O_11_1_0 = other_ops_10_O_1_0; // @[Map2S.scala 24:12]
  assign O_11_1_1 = other_ops_10_O_1_1; // @[Map2S.scala 24:12]
  assign O_11_1_2 = other_ops_10_O_1_2; // @[Map2S.scala 24:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[Map2S.scala 24:12]
  assign O_12_0_1 = other_ops_11_O_0_1; // @[Map2S.scala 24:12]
  assign O_12_0_2 = other_ops_11_O_0_2; // @[Map2S.scala 24:12]
  assign O_12_1_0 = other_ops_11_O_1_0; // @[Map2S.scala 24:12]
  assign O_12_1_1 = other_ops_11_O_1_1; // @[Map2S.scala 24:12]
  assign O_12_1_2 = other_ops_11_O_1_2; // @[Map2S.scala 24:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[Map2S.scala 24:12]
  assign O_13_0_1 = other_ops_12_O_0_1; // @[Map2S.scala 24:12]
  assign O_13_0_2 = other_ops_12_O_0_2; // @[Map2S.scala 24:12]
  assign O_13_1_0 = other_ops_12_O_1_0; // @[Map2S.scala 24:12]
  assign O_13_1_1 = other_ops_12_O_1_1; // @[Map2S.scala 24:12]
  assign O_13_1_2 = other_ops_12_O_1_2; // @[Map2S.scala 24:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[Map2S.scala 24:12]
  assign O_14_0_1 = other_ops_13_O_0_1; // @[Map2S.scala 24:12]
  assign O_14_0_2 = other_ops_13_O_0_2; // @[Map2S.scala 24:12]
  assign O_14_1_0 = other_ops_13_O_1_0; // @[Map2S.scala 24:12]
  assign O_14_1_1 = other_ops_13_O_1_1; // @[Map2S.scala 24:12]
  assign O_14_1_2 = other_ops_13_O_1_2; // @[Map2S.scala 24:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[Map2S.scala 24:12]
  assign O_15_0_1 = other_ops_14_O_0_1; // @[Map2S.scala 24:12]
  assign O_15_0_2 = other_ops_14_O_0_2; // @[Map2S.scala 24:12]
  assign O_15_1_0 = other_ops_14_O_1_0; // @[Map2S.scala 24:12]
  assign O_15_1_1 = other_ops_14_O_1_1; // @[Map2S.scala 24:12]
  assign O_15_1_2 = other_ops_14_O_1_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2 = I0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = I1_1_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = I1_1_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = I1_1_2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2 = I0_2_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = I1_2_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = I1_2_1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = I1_2_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0 = I0_3_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1 = I0_3_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_2 = I0_3_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0 = I1_3_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_1 = I1_3_1; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_2 = I1_3_2; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0 = I0_4_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1 = I0_4_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_2 = I0_4_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0 = I1_4_0; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_1 = I1_4_1; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_2 = I1_4_2; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0 = I0_5_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1 = I0_5_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_2 = I0_5_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0 = I1_5_0; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_1 = I1_5_1; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_2 = I1_5_2; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0 = I0_6_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1 = I0_6_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_2 = I0_6_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0 = I1_6_0; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_1 = I1_6_1; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_2 = I1_6_2; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0 = I0_7_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1 = I0_7_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_2 = I0_7_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0 = I1_7_0; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_1 = I1_7_1; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_2 = I1_7_2; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0 = I0_8_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1 = I0_8_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_2 = I0_8_2; // @[Map2S.scala 22:43]
  assign other_ops_7_I1_0 = I1_8_0; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_1 = I1_8_1; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_2 = I1_8_2; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0 = I0_9_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1 = I0_9_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_2 = I0_9_2; // @[Map2S.scala 22:43]
  assign other_ops_8_I1_0 = I1_9_0; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_1 = I1_9_1; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_2 = I1_9_2; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0 = I0_10_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1 = I0_10_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_2 = I0_10_2; // @[Map2S.scala 22:43]
  assign other_ops_9_I1_0 = I1_10_0; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_1 = I1_10_1; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_2 = I1_10_2; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0 = I0_11_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1 = I0_11_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_2 = I0_11_2; // @[Map2S.scala 22:43]
  assign other_ops_10_I1_0 = I1_11_0; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_1 = I1_11_1; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_2 = I1_11_2; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0 = I0_12_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1 = I0_12_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_2 = I0_12_2; // @[Map2S.scala 22:43]
  assign other_ops_11_I1_0 = I1_12_0; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_1 = I1_12_1; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_2 = I1_12_2; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0 = I0_13_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1 = I0_13_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_2 = I0_13_2; // @[Map2S.scala 22:43]
  assign other_ops_12_I1_0 = I1_13_0; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_1 = I1_13_1; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_2 = I1_13_2; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0 = I0_14_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1 = I0_14_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_2 = I0_14_2; // @[Map2S.scala 22:43]
  assign other_ops_13_I1_0 = I1_14_0; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_1 = I1_14_1; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_2 = I1_14_2; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0 = I0_15_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1 = I0_15_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_2 = I0_15_2; // @[Map2S.scala 22:43]
  assign other_ops_14_I1_0 = I1_15_0; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_1 = I1_15_1; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_2 = I1_15_2; // @[Map2S.scala 23:43]
endmodule
module SSeqTupleAppender_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_0_2,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_1_2,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0_0 = I0_0_0; // @[Tuple.scala 24:34]
  assign O_0_1 = I0_0_1; // @[Tuple.scala 24:34]
  assign O_0_2 = I0_0_2; // @[Tuple.scala 24:34]
  assign O_1_0 = I0_1_0; // @[Tuple.scala 24:34]
  assign O_1_1 = I0_1_1; // @[Tuple.scala 24:34]
  assign O_1_2 = I0_1_2; // @[Tuple.scala 24:34]
  assign O_2_0 = I1_0; // @[Tuple.scala 26:32]
  assign O_2_1 = I1_1; // @[Tuple.scala 26:32]
  assign O_2_2 = I1_2; // @[Tuple.scala 26:32]
endmodule
module Map2S_7(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_0_0_1,
  input  [7:0] I0_0_0_2,
  input  [7:0] I0_0_1_0,
  input  [7:0] I0_0_1_1,
  input  [7:0] I0_0_1_2,
  input  [7:0] I0_1_0_0,
  input  [7:0] I0_1_0_1,
  input  [7:0] I0_1_0_2,
  input  [7:0] I0_1_1_0,
  input  [7:0] I0_1_1_1,
  input  [7:0] I0_1_1_2,
  input  [7:0] I0_2_0_0,
  input  [7:0] I0_2_0_1,
  input  [7:0] I0_2_0_2,
  input  [7:0] I0_2_1_0,
  input  [7:0] I0_2_1_1,
  input  [7:0] I0_2_1_2,
  input  [7:0] I0_3_0_0,
  input  [7:0] I0_3_0_1,
  input  [7:0] I0_3_0_2,
  input  [7:0] I0_3_1_0,
  input  [7:0] I0_3_1_1,
  input  [7:0] I0_3_1_2,
  input  [7:0] I0_4_0_0,
  input  [7:0] I0_4_0_1,
  input  [7:0] I0_4_0_2,
  input  [7:0] I0_4_1_0,
  input  [7:0] I0_4_1_1,
  input  [7:0] I0_4_1_2,
  input  [7:0] I0_5_0_0,
  input  [7:0] I0_5_0_1,
  input  [7:0] I0_5_0_2,
  input  [7:0] I0_5_1_0,
  input  [7:0] I0_5_1_1,
  input  [7:0] I0_5_1_2,
  input  [7:0] I0_6_0_0,
  input  [7:0] I0_6_0_1,
  input  [7:0] I0_6_0_2,
  input  [7:0] I0_6_1_0,
  input  [7:0] I0_6_1_1,
  input  [7:0] I0_6_1_2,
  input  [7:0] I0_7_0_0,
  input  [7:0] I0_7_0_1,
  input  [7:0] I0_7_0_2,
  input  [7:0] I0_7_1_0,
  input  [7:0] I0_7_1_1,
  input  [7:0] I0_7_1_2,
  input  [7:0] I0_8_0_0,
  input  [7:0] I0_8_0_1,
  input  [7:0] I0_8_0_2,
  input  [7:0] I0_8_1_0,
  input  [7:0] I0_8_1_1,
  input  [7:0] I0_8_1_2,
  input  [7:0] I0_9_0_0,
  input  [7:0] I0_9_0_1,
  input  [7:0] I0_9_0_2,
  input  [7:0] I0_9_1_0,
  input  [7:0] I0_9_1_1,
  input  [7:0] I0_9_1_2,
  input  [7:0] I0_10_0_0,
  input  [7:0] I0_10_0_1,
  input  [7:0] I0_10_0_2,
  input  [7:0] I0_10_1_0,
  input  [7:0] I0_10_1_1,
  input  [7:0] I0_10_1_2,
  input  [7:0] I0_11_0_0,
  input  [7:0] I0_11_0_1,
  input  [7:0] I0_11_0_2,
  input  [7:0] I0_11_1_0,
  input  [7:0] I0_11_1_1,
  input  [7:0] I0_11_1_2,
  input  [7:0] I0_12_0_0,
  input  [7:0] I0_12_0_1,
  input  [7:0] I0_12_0_2,
  input  [7:0] I0_12_1_0,
  input  [7:0] I0_12_1_1,
  input  [7:0] I0_12_1_2,
  input  [7:0] I0_13_0_0,
  input  [7:0] I0_13_0_1,
  input  [7:0] I0_13_0_2,
  input  [7:0] I0_13_1_0,
  input  [7:0] I0_13_1_1,
  input  [7:0] I0_13_1_2,
  input  [7:0] I0_14_0_0,
  input  [7:0] I0_14_0_1,
  input  [7:0] I0_14_0_2,
  input  [7:0] I0_14_1_0,
  input  [7:0] I0_14_1_1,
  input  [7:0] I0_14_1_2,
  input  [7:0] I0_15_0_0,
  input  [7:0] I0_15_0_1,
  input  [7:0] I0_15_0_2,
  input  [7:0] I0_15_1_0,
  input  [7:0] I0_15_1_1,
  input  [7:0] I0_15_1_2,
  input  [7:0] I1_0_0,
  input  [7:0] I1_0_1,
  input  [7:0] I1_0_2,
  input  [7:0] I1_1_0,
  input  [7:0] I1_1_1,
  input  [7:0] I1_1_2,
  input  [7:0] I1_2_0,
  input  [7:0] I1_2_1,
  input  [7:0] I1_2_2,
  input  [7:0] I1_3_0,
  input  [7:0] I1_3_1,
  input  [7:0] I1_3_2,
  input  [7:0] I1_4_0,
  input  [7:0] I1_4_1,
  input  [7:0] I1_4_2,
  input  [7:0] I1_5_0,
  input  [7:0] I1_5_1,
  input  [7:0] I1_5_2,
  input  [7:0] I1_6_0,
  input  [7:0] I1_6_1,
  input  [7:0] I1_6_2,
  input  [7:0] I1_7_0,
  input  [7:0] I1_7_1,
  input  [7:0] I1_7_2,
  input  [7:0] I1_8_0,
  input  [7:0] I1_8_1,
  input  [7:0] I1_8_2,
  input  [7:0] I1_9_0,
  input  [7:0] I1_9_1,
  input  [7:0] I1_9_2,
  input  [7:0] I1_10_0,
  input  [7:0] I1_10_1,
  input  [7:0] I1_10_2,
  input  [7:0] I1_11_0,
  input  [7:0] I1_11_1,
  input  [7:0] I1_11_2,
  input  [7:0] I1_12_0,
  input  [7:0] I1_12_1,
  input  [7:0] I1_12_2,
  input  [7:0] I1_13_0,
  input  [7:0] I1_13_1,
  input  [7:0] I1_13_2,
  input  [7:0] I1_14_0,
  input  [7:0] I1_14_1,
  input  [7:0] I1_14_2,
  input  [7:0] I1_15_0,
  input  [7:0] I1_15_1,
  input  [7:0] I1_15_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_0_2_0,
  output [7:0] O_0_2_1,
  output [7:0] O_0_2_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2,
  output [7:0] O_1_2_0,
  output [7:0] O_1_2_1,
  output [7:0] O_1_2_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_2_1_0,
  output [7:0] O_2_1_1,
  output [7:0] O_2_1_2,
  output [7:0] O_2_2_0,
  output [7:0] O_2_2_1,
  output [7:0] O_2_2_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_3_1_0,
  output [7:0] O_3_1_1,
  output [7:0] O_3_1_2,
  output [7:0] O_3_2_0,
  output [7:0] O_3_2_1,
  output [7:0] O_3_2_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_4_1_0,
  output [7:0] O_4_1_1,
  output [7:0] O_4_1_2,
  output [7:0] O_4_2_0,
  output [7:0] O_4_2_1,
  output [7:0] O_4_2_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_5_1_0,
  output [7:0] O_5_1_1,
  output [7:0] O_5_1_2,
  output [7:0] O_5_2_0,
  output [7:0] O_5_2_1,
  output [7:0] O_5_2_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_6_1_0,
  output [7:0] O_6_1_1,
  output [7:0] O_6_1_2,
  output [7:0] O_6_2_0,
  output [7:0] O_6_2_1,
  output [7:0] O_6_2_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2,
  output [7:0] O_7_1_0,
  output [7:0] O_7_1_1,
  output [7:0] O_7_1_2,
  output [7:0] O_7_2_0,
  output [7:0] O_7_2_1,
  output [7:0] O_7_2_2,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_0_2,
  output [7:0] O_8_1_0,
  output [7:0] O_8_1_1,
  output [7:0] O_8_1_2,
  output [7:0] O_8_2_0,
  output [7:0] O_8_2_1,
  output [7:0] O_8_2_2,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_0_2,
  output [7:0] O_9_1_0,
  output [7:0] O_9_1_1,
  output [7:0] O_9_1_2,
  output [7:0] O_9_2_0,
  output [7:0] O_9_2_1,
  output [7:0] O_9_2_2,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_0_2,
  output [7:0] O_10_1_0,
  output [7:0] O_10_1_1,
  output [7:0] O_10_1_2,
  output [7:0] O_10_2_0,
  output [7:0] O_10_2_1,
  output [7:0] O_10_2_2,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_0_2,
  output [7:0] O_11_1_0,
  output [7:0] O_11_1_1,
  output [7:0] O_11_1_2,
  output [7:0] O_11_2_0,
  output [7:0] O_11_2_1,
  output [7:0] O_11_2_2,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_0_2,
  output [7:0] O_12_1_0,
  output [7:0] O_12_1_1,
  output [7:0] O_12_1_2,
  output [7:0] O_12_2_0,
  output [7:0] O_12_2_1,
  output [7:0] O_12_2_2,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_0_2,
  output [7:0] O_13_1_0,
  output [7:0] O_13_1_1,
  output [7:0] O_13_1_2,
  output [7:0] O_13_2_0,
  output [7:0] O_13_2_1,
  output [7:0] O_13_2_2,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_0_2,
  output [7:0] O_14_1_0,
  output [7:0] O_14_1_1,
  output [7:0] O_14_1_2,
  output [7:0] O_14_2_0,
  output [7:0] O_14_2_1,
  output [7:0] O_14_2_2,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_0_2,
  output [7:0] O_15_1_0,
  output [7:0] O_15_1_1,
  output [7:0] O_15_1_2,
  output [7:0] O_15_2_0,
  output [7:0] O_15_2_1,
  output [7:0] O_15_2_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_2_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  SSeqTupleAppender_3 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I0_0_2(fst_op_I0_0_2),
    .I0_1_0(fst_op_I0_1_0),
    .I0_1_1(fst_op_I0_1_1),
    .I0_1_2(fst_op_I0_1_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0(other_ops_0_I0_0_0),
    .I0_0_1(other_ops_0_I0_0_1),
    .I0_0_2(other_ops_0_I0_0_2),
    .I0_1_0(other_ops_0_I0_1_0),
    .I0_1_1(other_ops_0_I0_1_1),
    .I0_1_2(other_ops_0_I0_1_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2),
    .O_2_0(other_ops_0_O_2_0),
    .O_2_1(other_ops_0_O_2_1),
    .O_2_2(other_ops_0_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0_0(other_ops_1_I0_0_0),
    .I0_0_1(other_ops_1_I0_0_1),
    .I0_0_2(other_ops_1_I0_0_2),
    .I0_1_0(other_ops_1_I0_1_0),
    .I0_1_1(other_ops_1_I0_1_1),
    .I0_1_2(other_ops_1_I0_1_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2),
    .O_2_0(other_ops_1_O_2_0),
    .O_2_1(other_ops_1_O_2_1),
    .O_2_2(other_ops_1_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0_0(other_ops_2_I0_0_0),
    .I0_0_1(other_ops_2_I0_0_1),
    .I0_0_2(other_ops_2_I0_0_2),
    .I0_1_0(other_ops_2_I0_1_0),
    .I0_1_1(other_ops_2_I0_1_1),
    .I0_1_2(other_ops_2_I0_1_2),
    .I1_0(other_ops_2_I1_0),
    .I1_1(other_ops_2_I1_1),
    .I1_2(other_ops_2_I1_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2),
    .O_2_0(other_ops_2_O_2_0),
    .O_2_1(other_ops_2_O_2_1),
    .O_2_2(other_ops_2_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0_0(other_ops_3_I0_0_0),
    .I0_0_1(other_ops_3_I0_0_1),
    .I0_0_2(other_ops_3_I0_0_2),
    .I0_1_0(other_ops_3_I0_1_0),
    .I0_1_1(other_ops_3_I0_1_1),
    .I0_1_2(other_ops_3_I0_1_2),
    .I1_0(other_ops_3_I1_0),
    .I1_1(other_ops_3_I1_1),
    .I1_2(other_ops_3_I1_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2),
    .O_2_0(other_ops_3_O_2_0),
    .O_2_1(other_ops_3_O_2_1),
    .O_2_2(other_ops_3_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0_0(other_ops_4_I0_0_0),
    .I0_0_1(other_ops_4_I0_0_1),
    .I0_0_2(other_ops_4_I0_0_2),
    .I0_1_0(other_ops_4_I0_1_0),
    .I0_1_1(other_ops_4_I0_1_1),
    .I0_1_2(other_ops_4_I0_1_2),
    .I1_0(other_ops_4_I1_0),
    .I1_1(other_ops_4_I1_1),
    .I1_2(other_ops_4_I1_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2),
    .O_2_0(other_ops_4_O_2_0),
    .O_2_1(other_ops_4_O_2_1),
    .O_2_2(other_ops_4_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0_0(other_ops_5_I0_0_0),
    .I0_0_1(other_ops_5_I0_0_1),
    .I0_0_2(other_ops_5_I0_0_2),
    .I0_1_0(other_ops_5_I0_1_0),
    .I0_1_1(other_ops_5_I0_1_1),
    .I0_1_2(other_ops_5_I0_1_2),
    .I1_0(other_ops_5_I1_0),
    .I1_1(other_ops_5_I1_1),
    .I1_2(other_ops_5_I1_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2),
    .O_2_0(other_ops_5_O_2_0),
    .O_2_1(other_ops_5_O_2_1),
    .O_2_2(other_ops_5_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0_0(other_ops_6_I0_0_0),
    .I0_0_1(other_ops_6_I0_0_1),
    .I0_0_2(other_ops_6_I0_0_2),
    .I0_1_0(other_ops_6_I0_1_0),
    .I0_1_1(other_ops_6_I0_1_1),
    .I0_1_2(other_ops_6_I0_1_2),
    .I1_0(other_ops_6_I1_0),
    .I1_1(other_ops_6_I1_1),
    .I1_2(other_ops_6_I1_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2),
    .O_2_0(other_ops_6_O_2_0),
    .O_2_1(other_ops_6_O_2_1),
    .O_2_2(other_ops_6_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0_0(other_ops_7_I0_0_0),
    .I0_0_1(other_ops_7_I0_0_1),
    .I0_0_2(other_ops_7_I0_0_2),
    .I0_1_0(other_ops_7_I0_1_0),
    .I0_1_1(other_ops_7_I0_1_1),
    .I0_1_2(other_ops_7_I0_1_2),
    .I1_0(other_ops_7_I1_0),
    .I1_1(other_ops_7_I1_1),
    .I1_2(other_ops_7_I1_2),
    .O_0_0(other_ops_7_O_0_0),
    .O_0_1(other_ops_7_O_0_1),
    .O_0_2(other_ops_7_O_0_2),
    .O_1_0(other_ops_7_O_1_0),
    .O_1_1(other_ops_7_O_1_1),
    .O_1_2(other_ops_7_O_1_2),
    .O_2_0(other_ops_7_O_2_0),
    .O_2_1(other_ops_7_O_2_1),
    .O_2_2(other_ops_7_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0_0(other_ops_8_I0_0_0),
    .I0_0_1(other_ops_8_I0_0_1),
    .I0_0_2(other_ops_8_I0_0_2),
    .I0_1_0(other_ops_8_I0_1_0),
    .I0_1_1(other_ops_8_I0_1_1),
    .I0_1_2(other_ops_8_I0_1_2),
    .I1_0(other_ops_8_I1_0),
    .I1_1(other_ops_8_I1_1),
    .I1_2(other_ops_8_I1_2),
    .O_0_0(other_ops_8_O_0_0),
    .O_0_1(other_ops_8_O_0_1),
    .O_0_2(other_ops_8_O_0_2),
    .O_1_0(other_ops_8_O_1_0),
    .O_1_1(other_ops_8_O_1_1),
    .O_1_2(other_ops_8_O_1_2),
    .O_2_0(other_ops_8_O_2_0),
    .O_2_1(other_ops_8_O_2_1),
    .O_2_2(other_ops_8_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0_0(other_ops_9_I0_0_0),
    .I0_0_1(other_ops_9_I0_0_1),
    .I0_0_2(other_ops_9_I0_0_2),
    .I0_1_0(other_ops_9_I0_1_0),
    .I0_1_1(other_ops_9_I0_1_1),
    .I0_1_2(other_ops_9_I0_1_2),
    .I1_0(other_ops_9_I1_0),
    .I1_1(other_ops_9_I1_1),
    .I1_2(other_ops_9_I1_2),
    .O_0_0(other_ops_9_O_0_0),
    .O_0_1(other_ops_9_O_0_1),
    .O_0_2(other_ops_9_O_0_2),
    .O_1_0(other_ops_9_O_1_0),
    .O_1_1(other_ops_9_O_1_1),
    .O_1_2(other_ops_9_O_1_2),
    .O_2_0(other_ops_9_O_2_0),
    .O_2_1(other_ops_9_O_2_1),
    .O_2_2(other_ops_9_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0_0(other_ops_10_I0_0_0),
    .I0_0_1(other_ops_10_I0_0_1),
    .I0_0_2(other_ops_10_I0_0_2),
    .I0_1_0(other_ops_10_I0_1_0),
    .I0_1_1(other_ops_10_I0_1_1),
    .I0_1_2(other_ops_10_I0_1_2),
    .I1_0(other_ops_10_I1_0),
    .I1_1(other_ops_10_I1_1),
    .I1_2(other_ops_10_I1_2),
    .O_0_0(other_ops_10_O_0_0),
    .O_0_1(other_ops_10_O_0_1),
    .O_0_2(other_ops_10_O_0_2),
    .O_1_0(other_ops_10_O_1_0),
    .O_1_1(other_ops_10_O_1_1),
    .O_1_2(other_ops_10_O_1_2),
    .O_2_0(other_ops_10_O_2_0),
    .O_2_1(other_ops_10_O_2_1),
    .O_2_2(other_ops_10_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0_0(other_ops_11_I0_0_0),
    .I0_0_1(other_ops_11_I0_0_1),
    .I0_0_2(other_ops_11_I0_0_2),
    .I0_1_0(other_ops_11_I0_1_0),
    .I0_1_1(other_ops_11_I0_1_1),
    .I0_1_2(other_ops_11_I0_1_2),
    .I1_0(other_ops_11_I1_0),
    .I1_1(other_ops_11_I1_1),
    .I1_2(other_ops_11_I1_2),
    .O_0_0(other_ops_11_O_0_0),
    .O_0_1(other_ops_11_O_0_1),
    .O_0_2(other_ops_11_O_0_2),
    .O_1_0(other_ops_11_O_1_0),
    .O_1_1(other_ops_11_O_1_1),
    .O_1_2(other_ops_11_O_1_2),
    .O_2_0(other_ops_11_O_2_0),
    .O_2_1(other_ops_11_O_2_1),
    .O_2_2(other_ops_11_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0_0(other_ops_12_I0_0_0),
    .I0_0_1(other_ops_12_I0_0_1),
    .I0_0_2(other_ops_12_I0_0_2),
    .I0_1_0(other_ops_12_I0_1_0),
    .I0_1_1(other_ops_12_I0_1_1),
    .I0_1_2(other_ops_12_I0_1_2),
    .I1_0(other_ops_12_I1_0),
    .I1_1(other_ops_12_I1_1),
    .I1_2(other_ops_12_I1_2),
    .O_0_0(other_ops_12_O_0_0),
    .O_0_1(other_ops_12_O_0_1),
    .O_0_2(other_ops_12_O_0_2),
    .O_1_0(other_ops_12_O_1_0),
    .O_1_1(other_ops_12_O_1_1),
    .O_1_2(other_ops_12_O_1_2),
    .O_2_0(other_ops_12_O_2_0),
    .O_2_1(other_ops_12_O_2_1),
    .O_2_2(other_ops_12_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0_0(other_ops_13_I0_0_0),
    .I0_0_1(other_ops_13_I0_0_1),
    .I0_0_2(other_ops_13_I0_0_2),
    .I0_1_0(other_ops_13_I0_1_0),
    .I0_1_1(other_ops_13_I0_1_1),
    .I0_1_2(other_ops_13_I0_1_2),
    .I1_0(other_ops_13_I1_0),
    .I1_1(other_ops_13_I1_1),
    .I1_2(other_ops_13_I1_2),
    .O_0_0(other_ops_13_O_0_0),
    .O_0_1(other_ops_13_O_0_1),
    .O_0_2(other_ops_13_O_0_2),
    .O_1_0(other_ops_13_O_1_0),
    .O_1_1(other_ops_13_O_1_1),
    .O_1_2(other_ops_13_O_1_2),
    .O_2_0(other_ops_13_O_2_0),
    .O_2_1(other_ops_13_O_2_1),
    .O_2_2(other_ops_13_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0_0(other_ops_14_I0_0_0),
    .I0_0_1(other_ops_14_I0_0_1),
    .I0_0_2(other_ops_14_I0_0_2),
    .I0_1_0(other_ops_14_I0_1_0),
    .I0_1_1(other_ops_14_I0_1_1),
    .I0_1_2(other_ops_14_I0_1_2),
    .I1_0(other_ops_14_I1_0),
    .I1_1(other_ops_14_I1_1),
    .I1_2(other_ops_14_I1_2),
    .O_0_0(other_ops_14_O_0_0),
    .O_0_1(other_ops_14_O_0_1),
    .O_0_2(other_ops_14_O_0_2),
    .O_1_0(other_ops_14_O_1_0),
    .O_1_1(other_ops_14_O_1_1),
    .O_1_2(other_ops_14_O_1_2),
    .O_2_0(other_ops_14_O_2_0),
    .O_2_1(other_ops_14_O_2_1),
    .O_2_2(other_ops_14_O_2_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[Map2S.scala 19:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[Map2S.scala 19:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[Map2S.scala 24:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[Map2S.scala 24:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[Map2S.scala 24:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[Map2S.scala 24:12]
  assign O_1_2_0 = other_ops_0_O_2_0; // @[Map2S.scala 24:12]
  assign O_1_2_1 = other_ops_0_O_2_1; // @[Map2S.scala 24:12]
  assign O_1_2_2 = other_ops_0_O_2_2; // @[Map2S.scala 24:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[Map2S.scala 24:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[Map2S.scala 24:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[Map2S.scala 24:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[Map2S.scala 24:12]
  assign O_2_2_0 = other_ops_1_O_2_0; // @[Map2S.scala 24:12]
  assign O_2_2_1 = other_ops_1_O_2_1; // @[Map2S.scala 24:12]
  assign O_2_2_2 = other_ops_1_O_2_2; // @[Map2S.scala 24:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[Map2S.scala 24:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[Map2S.scala 24:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[Map2S.scala 24:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[Map2S.scala 24:12]
  assign O_3_2_0 = other_ops_2_O_2_0; // @[Map2S.scala 24:12]
  assign O_3_2_1 = other_ops_2_O_2_1; // @[Map2S.scala 24:12]
  assign O_3_2_2 = other_ops_2_O_2_2; // @[Map2S.scala 24:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[Map2S.scala 24:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[Map2S.scala 24:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[Map2S.scala 24:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[Map2S.scala 24:12]
  assign O_4_2_0 = other_ops_3_O_2_0; // @[Map2S.scala 24:12]
  assign O_4_2_1 = other_ops_3_O_2_1; // @[Map2S.scala 24:12]
  assign O_4_2_2 = other_ops_3_O_2_2; // @[Map2S.scala 24:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[Map2S.scala 24:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[Map2S.scala 24:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[Map2S.scala 24:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[Map2S.scala 24:12]
  assign O_5_2_0 = other_ops_4_O_2_0; // @[Map2S.scala 24:12]
  assign O_5_2_1 = other_ops_4_O_2_1; // @[Map2S.scala 24:12]
  assign O_5_2_2 = other_ops_4_O_2_2; // @[Map2S.scala 24:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[Map2S.scala 24:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[Map2S.scala 24:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[Map2S.scala 24:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[Map2S.scala 24:12]
  assign O_6_2_0 = other_ops_5_O_2_0; // @[Map2S.scala 24:12]
  assign O_6_2_1 = other_ops_5_O_2_1; // @[Map2S.scala 24:12]
  assign O_6_2_2 = other_ops_5_O_2_2; // @[Map2S.scala 24:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[Map2S.scala 24:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[Map2S.scala 24:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[Map2S.scala 24:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[Map2S.scala 24:12]
  assign O_7_2_0 = other_ops_6_O_2_0; // @[Map2S.scala 24:12]
  assign O_7_2_1 = other_ops_6_O_2_1; // @[Map2S.scala 24:12]
  assign O_7_2_2 = other_ops_6_O_2_2; // @[Map2S.scala 24:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[Map2S.scala 24:12]
  assign O_8_0_1 = other_ops_7_O_0_1; // @[Map2S.scala 24:12]
  assign O_8_0_2 = other_ops_7_O_0_2; // @[Map2S.scala 24:12]
  assign O_8_1_0 = other_ops_7_O_1_0; // @[Map2S.scala 24:12]
  assign O_8_1_1 = other_ops_7_O_1_1; // @[Map2S.scala 24:12]
  assign O_8_1_2 = other_ops_7_O_1_2; // @[Map2S.scala 24:12]
  assign O_8_2_0 = other_ops_7_O_2_0; // @[Map2S.scala 24:12]
  assign O_8_2_1 = other_ops_7_O_2_1; // @[Map2S.scala 24:12]
  assign O_8_2_2 = other_ops_7_O_2_2; // @[Map2S.scala 24:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[Map2S.scala 24:12]
  assign O_9_0_1 = other_ops_8_O_0_1; // @[Map2S.scala 24:12]
  assign O_9_0_2 = other_ops_8_O_0_2; // @[Map2S.scala 24:12]
  assign O_9_1_0 = other_ops_8_O_1_0; // @[Map2S.scala 24:12]
  assign O_9_1_1 = other_ops_8_O_1_1; // @[Map2S.scala 24:12]
  assign O_9_1_2 = other_ops_8_O_1_2; // @[Map2S.scala 24:12]
  assign O_9_2_0 = other_ops_8_O_2_0; // @[Map2S.scala 24:12]
  assign O_9_2_1 = other_ops_8_O_2_1; // @[Map2S.scala 24:12]
  assign O_9_2_2 = other_ops_8_O_2_2; // @[Map2S.scala 24:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[Map2S.scala 24:12]
  assign O_10_0_1 = other_ops_9_O_0_1; // @[Map2S.scala 24:12]
  assign O_10_0_2 = other_ops_9_O_0_2; // @[Map2S.scala 24:12]
  assign O_10_1_0 = other_ops_9_O_1_0; // @[Map2S.scala 24:12]
  assign O_10_1_1 = other_ops_9_O_1_1; // @[Map2S.scala 24:12]
  assign O_10_1_2 = other_ops_9_O_1_2; // @[Map2S.scala 24:12]
  assign O_10_2_0 = other_ops_9_O_2_0; // @[Map2S.scala 24:12]
  assign O_10_2_1 = other_ops_9_O_2_1; // @[Map2S.scala 24:12]
  assign O_10_2_2 = other_ops_9_O_2_2; // @[Map2S.scala 24:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[Map2S.scala 24:12]
  assign O_11_0_1 = other_ops_10_O_0_1; // @[Map2S.scala 24:12]
  assign O_11_0_2 = other_ops_10_O_0_2; // @[Map2S.scala 24:12]
  assign O_11_1_0 = other_ops_10_O_1_0; // @[Map2S.scala 24:12]
  assign O_11_1_1 = other_ops_10_O_1_1; // @[Map2S.scala 24:12]
  assign O_11_1_2 = other_ops_10_O_1_2; // @[Map2S.scala 24:12]
  assign O_11_2_0 = other_ops_10_O_2_0; // @[Map2S.scala 24:12]
  assign O_11_2_1 = other_ops_10_O_2_1; // @[Map2S.scala 24:12]
  assign O_11_2_2 = other_ops_10_O_2_2; // @[Map2S.scala 24:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[Map2S.scala 24:12]
  assign O_12_0_1 = other_ops_11_O_0_1; // @[Map2S.scala 24:12]
  assign O_12_0_2 = other_ops_11_O_0_2; // @[Map2S.scala 24:12]
  assign O_12_1_0 = other_ops_11_O_1_0; // @[Map2S.scala 24:12]
  assign O_12_1_1 = other_ops_11_O_1_1; // @[Map2S.scala 24:12]
  assign O_12_1_2 = other_ops_11_O_1_2; // @[Map2S.scala 24:12]
  assign O_12_2_0 = other_ops_11_O_2_0; // @[Map2S.scala 24:12]
  assign O_12_2_1 = other_ops_11_O_2_1; // @[Map2S.scala 24:12]
  assign O_12_2_2 = other_ops_11_O_2_2; // @[Map2S.scala 24:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[Map2S.scala 24:12]
  assign O_13_0_1 = other_ops_12_O_0_1; // @[Map2S.scala 24:12]
  assign O_13_0_2 = other_ops_12_O_0_2; // @[Map2S.scala 24:12]
  assign O_13_1_0 = other_ops_12_O_1_0; // @[Map2S.scala 24:12]
  assign O_13_1_1 = other_ops_12_O_1_1; // @[Map2S.scala 24:12]
  assign O_13_1_2 = other_ops_12_O_1_2; // @[Map2S.scala 24:12]
  assign O_13_2_0 = other_ops_12_O_2_0; // @[Map2S.scala 24:12]
  assign O_13_2_1 = other_ops_12_O_2_1; // @[Map2S.scala 24:12]
  assign O_13_2_2 = other_ops_12_O_2_2; // @[Map2S.scala 24:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[Map2S.scala 24:12]
  assign O_14_0_1 = other_ops_13_O_0_1; // @[Map2S.scala 24:12]
  assign O_14_0_2 = other_ops_13_O_0_2; // @[Map2S.scala 24:12]
  assign O_14_1_0 = other_ops_13_O_1_0; // @[Map2S.scala 24:12]
  assign O_14_1_1 = other_ops_13_O_1_1; // @[Map2S.scala 24:12]
  assign O_14_1_2 = other_ops_13_O_1_2; // @[Map2S.scala 24:12]
  assign O_14_2_0 = other_ops_13_O_2_0; // @[Map2S.scala 24:12]
  assign O_14_2_1 = other_ops_13_O_2_1; // @[Map2S.scala 24:12]
  assign O_14_2_2 = other_ops_13_O_2_2; // @[Map2S.scala 24:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[Map2S.scala 24:12]
  assign O_15_0_1 = other_ops_14_O_0_1; // @[Map2S.scala 24:12]
  assign O_15_0_2 = other_ops_14_O_0_2; // @[Map2S.scala 24:12]
  assign O_15_1_0 = other_ops_14_O_1_0; // @[Map2S.scala 24:12]
  assign O_15_1_1 = other_ops_14_O_1_1; // @[Map2S.scala 24:12]
  assign O_15_1_2 = other_ops_14_O_1_2; // @[Map2S.scala 24:12]
  assign O_15_2_0 = other_ops_14_O_2_0; // @[Map2S.scala 24:12]
  assign O_15_2_1 = other_ops_14_O_2_1; // @[Map2S.scala 24:12]
  assign O_15_2_2 = other_ops_14_O_2_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_2 = I0_0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_0 = I0_0_1_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_1 = I0_0_1_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_2 = I0_0_1_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0 = I0_1_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_1 = I0_1_0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_2 = I0_1_0_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_0 = I0_1_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_1 = I0_1_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_2 = I0_1_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = I1_1_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = I1_1_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = I1_1_2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0_0 = I0_2_0_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_1 = I0_2_0_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_2 = I0_2_0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_0 = I0_2_1_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_1 = I0_2_1_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_2 = I0_2_1_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = I1_2_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = I1_2_1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = I1_2_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0_0 = I0_3_0_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_1 = I0_3_0_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_2 = I0_3_0_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_0 = I0_3_1_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_1 = I0_3_1_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_2 = I0_3_1_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0 = I1_3_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_1 = I1_3_1; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_2 = I1_3_2; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0_0 = I0_4_0_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_1 = I0_4_0_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_2 = I0_4_0_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_0 = I0_4_1_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_1 = I0_4_1_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_2 = I0_4_1_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0 = I1_4_0; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_1 = I1_4_1; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_2 = I1_4_2; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0_0 = I0_5_0_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_1 = I0_5_0_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_2 = I0_5_0_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_0 = I0_5_1_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_1 = I0_5_1_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_2 = I0_5_1_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0 = I1_5_0; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_1 = I1_5_1; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_2 = I1_5_2; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0_0 = I0_6_0_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_1 = I0_6_0_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_2 = I0_6_0_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_0 = I0_6_1_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_1 = I0_6_1_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_2 = I0_6_1_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0 = I1_6_0; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_1 = I1_6_1; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_2 = I1_6_2; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0_0 = I0_7_0_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_1 = I0_7_0_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_2 = I0_7_0_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_0 = I0_7_1_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_1 = I0_7_1_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_2 = I0_7_1_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0 = I1_7_0; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_1 = I1_7_1; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_2 = I1_7_2; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0_0 = I0_8_0_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_0_1 = I0_8_0_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_0_2 = I0_8_0_2; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1_0 = I0_8_1_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1_1 = I0_8_1_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1_2 = I0_8_1_2; // @[Map2S.scala 22:43]
  assign other_ops_7_I1_0 = I1_8_0; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_1 = I1_8_1; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_2 = I1_8_2; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0_0 = I0_9_0_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_0_1 = I0_9_0_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_0_2 = I0_9_0_2; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1_0 = I0_9_1_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1_1 = I0_9_1_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1_2 = I0_9_1_2; // @[Map2S.scala 22:43]
  assign other_ops_8_I1_0 = I1_9_0; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_1 = I1_9_1; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_2 = I1_9_2; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0_0 = I0_10_0_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_0_1 = I0_10_0_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_0_2 = I0_10_0_2; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1_0 = I0_10_1_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1_1 = I0_10_1_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1_2 = I0_10_1_2; // @[Map2S.scala 22:43]
  assign other_ops_9_I1_0 = I1_10_0; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_1 = I1_10_1; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_2 = I1_10_2; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0_0 = I0_11_0_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_0_1 = I0_11_0_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_0_2 = I0_11_0_2; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1_0 = I0_11_1_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1_1 = I0_11_1_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1_2 = I0_11_1_2; // @[Map2S.scala 22:43]
  assign other_ops_10_I1_0 = I1_11_0; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_1 = I1_11_1; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_2 = I1_11_2; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0_0 = I0_12_0_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_0_1 = I0_12_0_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_0_2 = I0_12_0_2; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1_0 = I0_12_1_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1_1 = I0_12_1_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1_2 = I0_12_1_2; // @[Map2S.scala 22:43]
  assign other_ops_11_I1_0 = I1_12_0; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_1 = I1_12_1; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_2 = I1_12_2; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0_0 = I0_13_0_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_0_1 = I0_13_0_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_0_2 = I0_13_0_2; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1_0 = I0_13_1_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1_1 = I0_13_1_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1_2 = I0_13_1_2; // @[Map2S.scala 22:43]
  assign other_ops_12_I1_0 = I1_13_0; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_1 = I1_13_1; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_2 = I1_13_2; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0_0 = I0_14_0_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_0_1 = I0_14_0_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_0_2 = I0_14_0_2; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1_0 = I0_14_1_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1_1 = I0_14_1_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1_2 = I0_14_1_2; // @[Map2S.scala 22:43]
  assign other_ops_13_I1_0 = I1_14_0; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_1 = I1_14_1; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_2 = I1_14_2; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0_0 = I0_15_0_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_0_1 = I0_15_0_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_0_2 = I0_15_0_2; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1_0 = I0_15_1_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1_1 = I0_15_1_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1_2 = I0_15_1_2; // @[Map2S.scala 22:43]
  assign other_ops_14_I1_0 = I1_15_0; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_1 = I1_15_1; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_2 = I1_15_2; // @[Map2S.scala 23:43]
endmodule
module PartitionS_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  input  [7:0] I_1_1_0,
  input  [7:0] I_1_1_1,
  input  [7:0] I_1_1_2,
  input  [7:0] I_1_2_0,
  input  [7:0] I_1_2_1,
  input  [7:0] I_1_2_2,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_2_0_2,
  input  [7:0] I_2_1_0,
  input  [7:0] I_2_1_1,
  input  [7:0] I_2_1_2,
  input  [7:0] I_2_2_0,
  input  [7:0] I_2_2_1,
  input  [7:0] I_2_2_2,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_3_0_2,
  input  [7:0] I_3_1_0,
  input  [7:0] I_3_1_1,
  input  [7:0] I_3_1_2,
  input  [7:0] I_3_2_0,
  input  [7:0] I_3_2_1,
  input  [7:0] I_3_2_2,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_4_0_2,
  input  [7:0] I_4_1_0,
  input  [7:0] I_4_1_1,
  input  [7:0] I_4_1_2,
  input  [7:0] I_4_2_0,
  input  [7:0] I_4_2_1,
  input  [7:0] I_4_2_2,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_5_0_2,
  input  [7:0] I_5_1_0,
  input  [7:0] I_5_1_1,
  input  [7:0] I_5_1_2,
  input  [7:0] I_5_2_0,
  input  [7:0] I_5_2_1,
  input  [7:0] I_5_2_2,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_6_0_2,
  input  [7:0] I_6_1_0,
  input  [7:0] I_6_1_1,
  input  [7:0] I_6_1_2,
  input  [7:0] I_6_2_0,
  input  [7:0] I_6_2_1,
  input  [7:0] I_6_2_2,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_7_0_2,
  input  [7:0] I_7_1_0,
  input  [7:0] I_7_1_1,
  input  [7:0] I_7_1_2,
  input  [7:0] I_7_2_0,
  input  [7:0] I_7_2_1,
  input  [7:0] I_7_2_2,
  input  [7:0] I_8_0_0,
  input  [7:0] I_8_0_1,
  input  [7:0] I_8_0_2,
  input  [7:0] I_8_1_0,
  input  [7:0] I_8_1_1,
  input  [7:0] I_8_1_2,
  input  [7:0] I_8_2_0,
  input  [7:0] I_8_2_1,
  input  [7:0] I_8_2_2,
  input  [7:0] I_9_0_0,
  input  [7:0] I_9_0_1,
  input  [7:0] I_9_0_2,
  input  [7:0] I_9_1_0,
  input  [7:0] I_9_1_1,
  input  [7:0] I_9_1_2,
  input  [7:0] I_9_2_0,
  input  [7:0] I_9_2_1,
  input  [7:0] I_9_2_2,
  input  [7:0] I_10_0_0,
  input  [7:0] I_10_0_1,
  input  [7:0] I_10_0_2,
  input  [7:0] I_10_1_0,
  input  [7:0] I_10_1_1,
  input  [7:0] I_10_1_2,
  input  [7:0] I_10_2_0,
  input  [7:0] I_10_2_1,
  input  [7:0] I_10_2_2,
  input  [7:0] I_11_0_0,
  input  [7:0] I_11_0_1,
  input  [7:0] I_11_0_2,
  input  [7:0] I_11_1_0,
  input  [7:0] I_11_1_1,
  input  [7:0] I_11_1_2,
  input  [7:0] I_11_2_0,
  input  [7:0] I_11_2_1,
  input  [7:0] I_11_2_2,
  input  [7:0] I_12_0_0,
  input  [7:0] I_12_0_1,
  input  [7:0] I_12_0_2,
  input  [7:0] I_12_1_0,
  input  [7:0] I_12_1_1,
  input  [7:0] I_12_1_2,
  input  [7:0] I_12_2_0,
  input  [7:0] I_12_2_1,
  input  [7:0] I_12_2_2,
  input  [7:0] I_13_0_0,
  input  [7:0] I_13_0_1,
  input  [7:0] I_13_0_2,
  input  [7:0] I_13_1_0,
  input  [7:0] I_13_1_1,
  input  [7:0] I_13_1_2,
  input  [7:0] I_13_2_0,
  input  [7:0] I_13_2_1,
  input  [7:0] I_13_2_2,
  input  [7:0] I_14_0_0,
  input  [7:0] I_14_0_1,
  input  [7:0] I_14_0_2,
  input  [7:0] I_14_1_0,
  input  [7:0] I_14_1_1,
  input  [7:0] I_14_1_2,
  input  [7:0] I_14_2_0,
  input  [7:0] I_14_2_1,
  input  [7:0] I_14_2_2,
  input  [7:0] I_15_0_0,
  input  [7:0] I_15_0_1,
  input  [7:0] I_15_0_2,
  input  [7:0] I_15_1_0,
  input  [7:0] I_15_1_1,
  input  [7:0] I_15_1_2,
  input  [7:0] I_15_2_0,
  input  [7:0] I_15_2_1,
  input  [7:0] I_15_2_2,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_0_2,
  output [7:0] O_0_0_1_0,
  output [7:0] O_0_0_1_1,
  output [7:0] O_0_0_1_2,
  output [7:0] O_0_0_2_0,
  output [7:0] O_0_0_2_1,
  output [7:0] O_0_0_2_2,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_0_2,
  output [7:0] O_1_0_1_0,
  output [7:0] O_1_0_1_1,
  output [7:0] O_1_0_1_2,
  output [7:0] O_1_0_2_0,
  output [7:0] O_1_0_2_1,
  output [7:0] O_1_0_2_2,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_2_0_0_2,
  output [7:0] O_2_0_1_0,
  output [7:0] O_2_0_1_1,
  output [7:0] O_2_0_1_2,
  output [7:0] O_2_0_2_0,
  output [7:0] O_2_0_2_1,
  output [7:0] O_2_0_2_2,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_3_0_0_2,
  output [7:0] O_3_0_1_0,
  output [7:0] O_3_0_1_1,
  output [7:0] O_3_0_1_2,
  output [7:0] O_3_0_2_0,
  output [7:0] O_3_0_2_1,
  output [7:0] O_3_0_2_2,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_4_0_0_2,
  output [7:0] O_4_0_1_0,
  output [7:0] O_4_0_1_1,
  output [7:0] O_4_0_1_2,
  output [7:0] O_4_0_2_0,
  output [7:0] O_4_0_2_1,
  output [7:0] O_4_0_2_2,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_5_0_0_2,
  output [7:0] O_5_0_1_0,
  output [7:0] O_5_0_1_1,
  output [7:0] O_5_0_1_2,
  output [7:0] O_5_0_2_0,
  output [7:0] O_5_0_2_1,
  output [7:0] O_5_0_2_2,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_6_0_0_2,
  output [7:0] O_6_0_1_0,
  output [7:0] O_6_0_1_1,
  output [7:0] O_6_0_1_2,
  output [7:0] O_6_0_2_0,
  output [7:0] O_6_0_2_1,
  output [7:0] O_6_0_2_2,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_7_0_0_2,
  output [7:0] O_7_0_1_0,
  output [7:0] O_7_0_1_1,
  output [7:0] O_7_0_1_2,
  output [7:0] O_7_0_2_0,
  output [7:0] O_7_0_2_1,
  output [7:0] O_7_0_2_2,
  output [7:0] O_8_0_0_0,
  output [7:0] O_8_0_0_1,
  output [7:0] O_8_0_0_2,
  output [7:0] O_8_0_1_0,
  output [7:0] O_8_0_1_1,
  output [7:0] O_8_0_1_2,
  output [7:0] O_8_0_2_0,
  output [7:0] O_8_0_2_1,
  output [7:0] O_8_0_2_2,
  output [7:0] O_9_0_0_0,
  output [7:0] O_9_0_0_1,
  output [7:0] O_9_0_0_2,
  output [7:0] O_9_0_1_0,
  output [7:0] O_9_0_1_1,
  output [7:0] O_9_0_1_2,
  output [7:0] O_9_0_2_0,
  output [7:0] O_9_0_2_1,
  output [7:0] O_9_0_2_2,
  output [7:0] O_10_0_0_0,
  output [7:0] O_10_0_0_1,
  output [7:0] O_10_0_0_2,
  output [7:0] O_10_0_1_0,
  output [7:0] O_10_0_1_1,
  output [7:0] O_10_0_1_2,
  output [7:0] O_10_0_2_0,
  output [7:0] O_10_0_2_1,
  output [7:0] O_10_0_2_2,
  output [7:0] O_11_0_0_0,
  output [7:0] O_11_0_0_1,
  output [7:0] O_11_0_0_2,
  output [7:0] O_11_0_1_0,
  output [7:0] O_11_0_1_1,
  output [7:0] O_11_0_1_2,
  output [7:0] O_11_0_2_0,
  output [7:0] O_11_0_2_1,
  output [7:0] O_11_0_2_2,
  output [7:0] O_12_0_0_0,
  output [7:0] O_12_0_0_1,
  output [7:0] O_12_0_0_2,
  output [7:0] O_12_0_1_0,
  output [7:0] O_12_0_1_1,
  output [7:0] O_12_0_1_2,
  output [7:0] O_12_0_2_0,
  output [7:0] O_12_0_2_1,
  output [7:0] O_12_0_2_2,
  output [7:0] O_13_0_0_0,
  output [7:0] O_13_0_0_1,
  output [7:0] O_13_0_0_2,
  output [7:0] O_13_0_1_0,
  output [7:0] O_13_0_1_1,
  output [7:0] O_13_0_1_2,
  output [7:0] O_13_0_2_0,
  output [7:0] O_13_0_2_1,
  output [7:0] O_13_0_2_2,
  output [7:0] O_14_0_0_0,
  output [7:0] O_14_0_0_1,
  output [7:0] O_14_0_0_2,
  output [7:0] O_14_0_1_0,
  output [7:0] O_14_0_1_1,
  output [7:0] O_14_0_1_2,
  output [7:0] O_14_0_2_0,
  output [7:0] O_14_0_2_1,
  output [7:0] O_14_0_2_2,
  output [7:0] O_15_0_0_0,
  output [7:0] O_15_0_0_1,
  output [7:0] O_15_0_0_2,
  output [7:0] O_15_0_1_0,
  output [7:0] O_15_0_1_1,
  output [7:0] O_15_0_1_2,
  output [7:0] O_15_0_2_0,
  output [7:0] O_15_0_2_1,
  output [7:0] O_15_0_2_2
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0_0 = I_0_0_0; // @[Partition.scala 15:39]
  assign O_0_0_0_1 = I_0_0_1; // @[Partition.scala 15:39]
  assign O_0_0_0_2 = I_0_0_2; // @[Partition.scala 15:39]
  assign O_0_0_1_0 = I_0_1_0; // @[Partition.scala 15:39]
  assign O_0_0_1_1 = I_0_1_1; // @[Partition.scala 15:39]
  assign O_0_0_1_2 = I_0_1_2; // @[Partition.scala 15:39]
  assign O_0_0_2_0 = I_0_2_0; // @[Partition.scala 15:39]
  assign O_0_0_2_1 = I_0_2_1; // @[Partition.scala 15:39]
  assign O_0_0_2_2 = I_0_2_2; // @[Partition.scala 15:39]
  assign O_1_0_0_0 = I_1_0_0; // @[Partition.scala 15:39]
  assign O_1_0_0_1 = I_1_0_1; // @[Partition.scala 15:39]
  assign O_1_0_0_2 = I_1_0_2; // @[Partition.scala 15:39]
  assign O_1_0_1_0 = I_1_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1_1 = I_1_1_1; // @[Partition.scala 15:39]
  assign O_1_0_1_2 = I_1_1_2; // @[Partition.scala 15:39]
  assign O_1_0_2_0 = I_1_2_0; // @[Partition.scala 15:39]
  assign O_1_0_2_1 = I_1_2_1; // @[Partition.scala 15:39]
  assign O_1_0_2_2 = I_1_2_2; // @[Partition.scala 15:39]
  assign O_2_0_0_0 = I_2_0_0; // @[Partition.scala 15:39]
  assign O_2_0_0_1 = I_2_0_1; // @[Partition.scala 15:39]
  assign O_2_0_0_2 = I_2_0_2; // @[Partition.scala 15:39]
  assign O_2_0_1_0 = I_2_1_0; // @[Partition.scala 15:39]
  assign O_2_0_1_1 = I_2_1_1; // @[Partition.scala 15:39]
  assign O_2_0_1_2 = I_2_1_2; // @[Partition.scala 15:39]
  assign O_2_0_2_0 = I_2_2_0; // @[Partition.scala 15:39]
  assign O_2_0_2_1 = I_2_2_1; // @[Partition.scala 15:39]
  assign O_2_0_2_2 = I_2_2_2; // @[Partition.scala 15:39]
  assign O_3_0_0_0 = I_3_0_0; // @[Partition.scala 15:39]
  assign O_3_0_0_1 = I_3_0_1; // @[Partition.scala 15:39]
  assign O_3_0_0_2 = I_3_0_2; // @[Partition.scala 15:39]
  assign O_3_0_1_0 = I_3_1_0; // @[Partition.scala 15:39]
  assign O_3_0_1_1 = I_3_1_1; // @[Partition.scala 15:39]
  assign O_3_0_1_2 = I_3_1_2; // @[Partition.scala 15:39]
  assign O_3_0_2_0 = I_3_2_0; // @[Partition.scala 15:39]
  assign O_3_0_2_1 = I_3_2_1; // @[Partition.scala 15:39]
  assign O_3_0_2_2 = I_3_2_2; // @[Partition.scala 15:39]
  assign O_4_0_0_0 = I_4_0_0; // @[Partition.scala 15:39]
  assign O_4_0_0_1 = I_4_0_1; // @[Partition.scala 15:39]
  assign O_4_0_0_2 = I_4_0_2; // @[Partition.scala 15:39]
  assign O_4_0_1_0 = I_4_1_0; // @[Partition.scala 15:39]
  assign O_4_0_1_1 = I_4_1_1; // @[Partition.scala 15:39]
  assign O_4_0_1_2 = I_4_1_2; // @[Partition.scala 15:39]
  assign O_4_0_2_0 = I_4_2_0; // @[Partition.scala 15:39]
  assign O_4_0_2_1 = I_4_2_1; // @[Partition.scala 15:39]
  assign O_4_0_2_2 = I_4_2_2; // @[Partition.scala 15:39]
  assign O_5_0_0_0 = I_5_0_0; // @[Partition.scala 15:39]
  assign O_5_0_0_1 = I_5_0_1; // @[Partition.scala 15:39]
  assign O_5_0_0_2 = I_5_0_2; // @[Partition.scala 15:39]
  assign O_5_0_1_0 = I_5_1_0; // @[Partition.scala 15:39]
  assign O_5_0_1_1 = I_5_1_1; // @[Partition.scala 15:39]
  assign O_5_0_1_2 = I_5_1_2; // @[Partition.scala 15:39]
  assign O_5_0_2_0 = I_5_2_0; // @[Partition.scala 15:39]
  assign O_5_0_2_1 = I_5_2_1; // @[Partition.scala 15:39]
  assign O_5_0_2_2 = I_5_2_2; // @[Partition.scala 15:39]
  assign O_6_0_0_0 = I_6_0_0; // @[Partition.scala 15:39]
  assign O_6_0_0_1 = I_6_0_1; // @[Partition.scala 15:39]
  assign O_6_0_0_2 = I_6_0_2; // @[Partition.scala 15:39]
  assign O_6_0_1_0 = I_6_1_0; // @[Partition.scala 15:39]
  assign O_6_0_1_1 = I_6_1_1; // @[Partition.scala 15:39]
  assign O_6_0_1_2 = I_6_1_2; // @[Partition.scala 15:39]
  assign O_6_0_2_0 = I_6_2_0; // @[Partition.scala 15:39]
  assign O_6_0_2_1 = I_6_2_1; // @[Partition.scala 15:39]
  assign O_6_0_2_2 = I_6_2_2; // @[Partition.scala 15:39]
  assign O_7_0_0_0 = I_7_0_0; // @[Partition.scala 15:39]
  assign O_7_0_0_1 = I_7_0_1; // @[Partition.scala 15:39]
  assign O_7_0_0_2 = I_7_0_2; // @[Partition.scala 15:39]
  assign O_7_0_1_0 = I_7_1_0; // @[Partition.scala 15:39]
  assign O_7_0_1_1 = I_7_1_1; // @[Partition.scala 15:39]
  assign O_7_0_1_2 = I_7_1_2; // @[Partition.scala 15:39]
  assign O_7_0_2_0 = I_7_2_0; // @[Partition.scala 15:39]
  assign O_7_0_2_1 = I_7_2_1; // @[Partition.scala 15:39]
  assign O_7_0_2_2 = I_7_2_2; // @[Partition.scala 15:39]
  assign O_8_0_0_0 = I_8_0_0; // @[Partition.scala 15:39]
  assign O_8_0_0_1 = I_8_0_1; // @[Partition.scala 15:39]
  assign O_8_0_0_2 = I_8_0_2; // @[Partition.scala 15:39]
  assign O_8_0_1_0 = I_8_1_0; // @[Partition.scala 15:39]
  assign O_8_0_1_1 = I_8_1_1; // @[Partition.scala 15:39]
  assign O_8_0_1_2 = I_8_1_2; // @[Partition.scala 15:39]
  assign O_8_0_2_0 = I_8_2_0; // @[Partition.scala 15:39]
  assign O_8_0_2_1 = I_8_2_1; // @[Partition.scala 15:39]
  assign O_8_0_2_2 = I_8_2_2; // @[Partition.scala 15:39]
  assign O_9_0_0_0 = I_9_0_0; // @[Partition.scala 15:39]
  assign O_9_0_0_1 = I_9_0_1; // @[Partition.scala 15:39]
  assign O_9_0_0_2 = I_9_0_2; // @[Partition.scala 15:39]
  assign O_9_0_1_0 = I_9_1_0; // @[Partition.scala 15:39]
  assign O_9_0_1_1 = I_9_1_1; // @[Partition.scala 15:39]
  assign O_9_0_1_2 = I_9_1_2; // @[Partition.scala 15:39]
  assign O_9_0_2_0 = I_9_2_0; // @[Partition.scala 15:39]
  assign O_9_0_2_1 = I_9_2_1; // @[Partition.scala 15:39]
  assign O_9_0_2_2 = I_9_2_2; // @[Partition.scala 15:39]
  assign O_10_0_0_0 = I_10_0_0; // @[Partition.scala 15:39]
  assign O_10_0_0_1 = I_10_0_1; // @[Partition.scala 15:39]
  assign O_10_0_0_2 = I_10_0_2; // @[Partition.scala 15:39]
  assign O_10_0_1_0 = I_10_1_0; // @[Partition.scala 15:39]
  assign O_10_0_1_1 = I_10_1_1; // @[Partition.scala 15:39]
  assign O_10_0_1_2 = I_10_1_2; // @[Partition.scala 15:39]
  assign O_10_0_2_0 = I_10_2_0; // @[Partition.scala 15:39]
  assign O_10_0_2_1 = I_10_2_1; // @[Partition.scala 15:39]
  assign O_10_0_2_2 = I_10_2_2; // @[Partition.scala 15:39]
  assign O_11_0_0_0 = I_11_0_0; // @[Partition.scala 15:39]
  assign O_11_0_0_1 = I_11_0_1; // @[Partition.scala 15:39]
  assign O_11_0_0_2 = I_11_0_2; // @[Partition.scala 15:39]
  assign O_11_0_1_0 = I_11_1_0; // @[Partition.scala 15:39]
  assign O_11_0_1_1 = I_11_1_1; // @[Partition.scala 15:39]
  assign O_11_0_1_2 = I_11_1_2; // @[Partition.scala 15:39]
  assign O_11_0_2_0 = I_11_2_0; // @[Partition.scala 15:39]
  assign O_11_0_2_1 = I_11_2_1; // @[Partition.scala 15:39]
  assign O_11_0_2_2 = I_11_2_2; // @[Partition.scala 15:39]
  assign O_12_0_0_0 = I_12_0_0; // @[Partition.scala 15:39]
  assign O_12_0_0_1 = I_12_0_1; // @[Partition.scala 15:39]
  assign O_12_0_0_2 = I_12_0_2; // @[Partition.scala 15:39]
  assign O_12_0_1_0 = I_12_1_0; // @[Partition.scala 15:39]
  assign O_12_0_1_1 = I_12_1_1; // @[Partition.scala 15:39]
  assign O_12_0_1_2 = I_12_1_2; // @[Partition.scala 15:39]
  assign O_12_0_2_0 = I_12_2_0; // @[Partition.scala 15:39]
  assign O_12_0_2_1 = I_12_2_1; // @[Partition.scala 15:39]
  assign O_12_0_2_2 = I_12_2_2; // @[Partition.scala 15:39]
  assign O_13_0_0_0 = I_13_0_0; // @[Partition.scala 15:39]
  assign O_13_0_0_1 = I_13_0_1; // @[Partition.scala 15:39]
  assign O_13_0_0_2 = I_13_0_2; // @[Partition.scala 15:39]
  assign O_13_0_1_0 = I_13_1_0; // @[Partition.scala 15:39]
  assign O_13_0_1_1 = I_13_1_1; // @[Partition.scala 15:39]
  assign O_13_0_1_2 = I_13_1_2; // @[Partition.scala 15:39]
  assign O_13_0_2_0 = I_13_2_0; // @[Partition.scala 15:39]
  assign O_13_0_2_1 = I_13_2_1; // @[Partition.scala 15:39]
  assign O_13_0_2_2 = I_13_2_2; // @[Partition.scala 15:39]
  assign O_14_0_0_0 = I_14_0_0; // @[Partition.scala 15:39]
  assign O_14_0_0_1 = I_14_0_1; // @[Partition.scala 15:39]
  assign O_14_0_0_2 = I_14_0_2; // @[Partition.scala 15:39]
  assign O_14_0_1_0 = I_14_1_0; // @[Partition.scala 15:39]
  assign O_14_0_1_1 = I_14_1_1; // @[Partition.scala 15:39]
  assign O_14_0_1_2 = I_14_1_2; // @[Partition.scala 15:39]
  assign O_14_0_2_0 = I_14_2_0; // @[Partition.scala 15:39]
  assign O_14_0_2_1 = I_14_2_1; // @[Partition.scala 15:39]
  assign O_14_0_2_2 = I_14_2_2; // @[Partition.scala 15:39]
  assign O_15_0_0_0 = I_15_0_0; // @[Partition.scala 15:39]
  assign O_15_0_0_1 = I_15_0_1; // @[Partition.scala 15:39]
  assign O_15_0_0_2 = I_15_0_2; // @[Partition.scala 15:39]
  assign O_15_0_1_0 = I_15_1_0; // @[Partition.scala 15:39]
  assign O_15_0_1_1 = I_15_1_1; // @[Partition.scala 15:39]
  assign O_15_0_1_2 = I_15_1_2; // @[Partition.scala 15:39]
  assign O_15_0_2_0 = I_15_2_0; // @[Partition.scala 15:39]
  assign O_15_0_2_1 = I_15_2_1; // @[Partition.scala 15:39]
  assign O_15_0_2_2 = I_15_2_2; // @[Partition.scala 15:39]
endmodule
module SSeqTupleToSSeq_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_2_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0_0 = I_0_0; // @[Tuple.scala 41:5]
  assign O_0_1 = I_0_1; // @[Tuple.scala 41:5]
  assign O_0_2 = I_0_2; // @[Tuple.scala 41:5]
  assign O_1_0 = I_1_0; // @[Tuple.scala 41:5]
  assign O_1_1 = I_1_1; // @[Tuple.scala 41:5]
  assign O_1_2 = I_1_2; // @[Tuple.scala 41:5]
  assign O_2_0 = I_2_0; // @[Tuple.scala 41:5]
  assign O_2_1 = I_2_1; // @[Tuple.scala 41:5]
  assign O_2_2 = I_2_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq_3 op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0_0(op_inst_I_0_0),
    .I_0_1(op_inst_I_0_1),
    .I_0_2(op_inst_I_0_2),
    .I_1_0(op_inst_I_1_0),
    .I_1_1(op_inst_I_1_1),
    .I_1_2(op_inst_I_1_2),
    .I_2_0(op_inst_I_2_0),
    .I_2_1(op_inst_I_2_1),
    .I_2_2(op_inst_I_2_2),
    .O_0_0(op_inst_O_0_0),
    .O_0_1(op_inst_O_0_1),
    .O_0_2(op_inst_O_0_2),
    .O_1_0(op_inst_O_1_0),
    .O_1_1(op_inst_O_1_1),
    .O_1_2(op_inst_O_1_2),
    .O_2_0(op_inst_O_2_0),
    .O_2_1(op_inst_O_2_1),
    .O_2_2(op_inst_O_2_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0_0 = op_inst_O_0_0; // @[Remove1S.scala 14:5]
  assign O_0_1 = op_inst_O_0_1; // @[Remove1S.scala 14:5]
  assign O_0_2 = op_inst_O_0_2; // @[Remove1S.scala 14:5]
  assign O_1_0 = op_inst_O_1_0; // @[Remove1S.scala 14:5]
  assign O_1_1 = op_inst_O_1_1; // @[Remove1S.scala 14:5]
  assign O_1_2 = op_inst_O_1_2; // @[Remove1S.scala 14:5]
  assign O_2_0 = op_inst_O_2_0; // @[Remove1S.scala 14:5]
  assign O_2_1 = op_inst_O_2_1; // @[Remove1S.scala 14:5]
  assign O_2_2 = op_inst_O_2_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0_0 = I_0_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_1 = I_0_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_2 = I_0_0_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_0 = I_0_1_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_1 = I_0_1_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_2 = I_0_1_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_0 = I_0_2_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_1 = I_0_2_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_2 = I_0_2_2; // @[Remove1S.scala 13:13]
endmodule
module MapS_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0_0,
  input  [7:0] I_0_0_0_1,
  input  [7:0] I_0_0_0_2,
  input  [7:0] I_0_0_1_0,
  input  [7:0] I_0_0_1_1,
  input  [7:0] I_0_0_1_2,
  input  [7:0] I_0_0_2_0,
  input  [7:0] I_0_0_2_1,
  input  [7:0] I_0_0_2_2,
  input  [7:0] I_1_0_0_0,
  input  [7:0] I_1_0_0_1,
  input  [7:0] I_1_0_0_2,
  input  [7:0] I_1_0_1_0,
  input  [7:0] I_1_0_1_1,
  input  [7:0] I_1_0_1_2,
  input  [7:0] I_1_0_2_0,
  input  [7:0] I_1_0_2_1,
  input  [7:0] I_1_0_2_2,
  input  [7:0] I_2_0_0_0,
  input  [7:0] I_2_0_0_1,
  input  [7:0] I_2_0_0_2,
  input  [7:0] I_2_0_1_0,
  input  [7:0] I_2_0_1_1,
  input  [7:0] I_2_0_1_2,
  input  [7:0] I_2_0_2_0,
  input  [7:0] I_2_0_2_1,
  input  [7:0] I_2_0_2_2,
  input  [7:0] I_3_0_0_0,
  input  [7:0] I_3_0_0_1,
  input  [7:0] I_3_0_0_2,
  input  [7:0] I_3_0_1_0,
  input  [7:0] I_3_0_1_1,
  input  [7:0] I_3_0_1_2,
  input  [7:0] I_3_0_2_0,
  input  [7:0] I_3_0_2_1,
  input  [7:0] I_3_0_2_2,
  input  [7:0] I_4_0_0_0,
  input  [7:0] I_4_0_0_1,
  input  [7:0] I_4_0_0_2,
  input  [7:0] I_4_0_1_0,
  input  [7:0] I_4_0_1_1,
  input  [7:0] I_4_0_1_2,
  input  [7:0] I_4_0_2_0,
  input  [7:0] I_4_0_2_1,
  input  [7:0] I_4_0_2_2,
  input  [7:0] I_5_0_0_0,
  input  [7:0] I_5_0_0_1,
  input  [7:0] I_5_0_0_2,
  input  [7:0] I_5_0_1_0,
  input  [7:0] I_5_0_1_1,
  input  [7:0] I_5_0_1_2,
  input  [7:0] I_5_0_2_0,
  input  [7:0] I_5_0_2_1,
  input  [7:0] I_5_0_2_2,
  input  [7:0] I_6_0_0_0,
  input  [7:0] I_6_0_0_1,
  input  [7:0] I_6_0_0_2,
  input  [7:0] I_6_0_1_0,
  input  [7:0] I_6_0_1_1,
  input  [7:0] I_6_0_1_2,
  input  [7:0] I_6_0_2_0,
  input  [7:0] I_6_0_2_1,
  input  [7:0] I_6_0_2_2,
  input  [7:0] I_7_0_0_0,
  input  [7:0] I_7_0_0_1,
  input  [7:0] I_7_0_0_2,
  input  [7:0] I_7_0_1_0,
  input  [7:0] I_7_0_1_1,
  input  [7:0] I_7_0_1_2,
  input  [7:0] I_7_0_2_0,
  input  [7:0] I_7_0_2_1,
  input  [7:0] I_7_0_2_2,
  input  [7:0] I_8_0_0_0,
  input  [7:0] I_8_0_0_1,
  input  [7:0] I_8_0_0_2,
  input  [7:0] I_8_0_1_0,
  input  [7:0] I_8_0_1_1,
  input  [7:0] I_8_0_1_2,
  input  [7:0] I_8_0_2_0,
  input  [7:0] I_8_0_2_1,
  input  [7:0] I_8_0_2_2,
  input  [7:0] I_9_0_0_0,
  input  [7:0] I_9_0_0_1,
  input  [7:0] I_9_0_0_2,
  input  [7:0] I_9_0_1_0,
  input  [7:0] I_9_0_1_1,
  input  [7:0] I_9_0_1_2,
  input  [7:0] I_9_0_2_0,
  input  [7:0] I_9_0_2_1,
  input  [7:0] I_9_0_2_2,
  input  [7:0] I_10_0_0_0,
  input  [7:0] I_10_0_0_1,
  input  [7:0] I_10_0_0_2,
  input  [7:0] I_10_0_1_0,
  input  [7:0] I_10_0_1_1,
  input  [7:0] I_10_0_1_2,
  input  [7:0] I_10_0_2_0,
  input  [7:0] I_10_0_2_1,
  input  [7:0] I_10_0_2_2,
  input  [7:0] I_11_0_0_0,
  input  [7:0] I_11_0_0_1,
  input  [7:0] I_11_0_0_2,
  input  [7:0] I_11_0_1_0,
  input  [7:0] I_11_0_1_1,
  input  [7:0] I_11_0_1_2,
  input  [7:0] I_11_0_2_0,
  input  [7:0] I_11_0_2_1,
  input  [7:0] I_11_0_2_2,
  input  [7:0] I_12_0_0_0,
  input  [7:0] I_12_0_0_1,
  input  [7:0] I_12_0_0_2,
  input  [7:0] I_12_0_1_0,
  input  [7:0] I_12_0_1_1,
  input  [7:0] I_12_0_1_2,
  input  [7:0] I_12_0_2_0,
  input  [7:0] I_12_0_2_1,
  input  [7:0] I_12_0_2_2,
  input  [7:0] I_13_0_0_0,
  input  [7:0] I_13_0_0_1,
  input  [7:0] I_13_0_0_2,
  input  [7:0] I_13_0_1_0,
  input  [7:0] I_13_0_1_1,
  input  [7:0] I_13_0_1_2,
  input  [7:0] I_13_0_2_0,
  input  [7:0] I_13_0_2_1,
  input  [7:0] I_13_0_2_2,
  input  [7:0] I_14_0_0_0,
  input  [7:0] I_14_0_0_1,
  input  [7:0] I_14_0_0_2,
  input  [7:0] I_14_0_1_0,
  input  [7:0] I_14_0_1_1,
  input  [7:0] I_14_0_1_2,
  input  [7:0] I_14_0_2_0,
  input  [7:0] I_14_0_2_1,
  input  [7:0] I_14_0_2_2,
  input  [7:0] I_15_0_0_0,
  input  [7:0] I_15_0_0_1,
  input  [7:0] I_15_0_0_2,
  input  [7:0] I_15_0_1_0,
  input  [7:0] I_15_0_1_1,
  input  [7:0] I_15_0_1_2,
  input  [7:0] I_15_0_2_0,
  input  [7:0] I_15_0_2_1,
  input  [7:0] I_15_0_2_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_0_2_0,
  output [7:0] O_0_2_1,
  output [7:0] O_0_2_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2,
  output [7:0] O_1_2_0,
  output [7:0] O_1_2_1,
  output [7:0] O_1_2_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_2_1_0,
  output [7:0] O_2_1_1,
  output [7:0] O_2_1_2,
  output [7:0] O_2_2_0,
  output [7:0] O_2_2_1,
  output [7:0] O_2_2_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_3_1_0,
  output [7:0] O_3_1_1,
  output [7:0] O_3_1_2,
  output [7:0] O_3_2_0,
  output [7:0] O_3_2_1,
  output [7:0] O_3_2_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_4_1_0,
  output [7:0] O_4_1_1,
  output [7:0] O_4_1_2,
  output [7:0] O_4_2_0,
  output [7:0] O_4_2_1,
  output [7:0] O_4_2_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_5_1_0,
  output [7:0] O_5_1_1,
  output [7:0] O_5_1_2,
  output [7:0] O_5_2_0,
  output [7:0] O_5_2_1,
  output [7:0] O_5_2_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_6_1_0,
  output [7:0] O_6_1_1,
  output [7:0] O_6_1_2,
  output [7:0] O_6_2_0,
  output [7:0] O_6_2_1,
  output [7:0] O_6_2_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2,
  output [7:0] O_7_1_0,
  output [7:0] O_7_1_1,
  output [7:0] O_7_1_2,
  output [7:0] O_7_2_0,
  output [7:0] O_7_2_1,
  output [7:0] O_7_2_2,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_0_2,
  output [7:0] O_8_1_0,
  output [7:0] O_8_1_1,
  output [7:0] O_8_1_2,
  output [7:0] O_8_2_0,
  output [7:0] O_8_2_1,
  output [7:0] O_8_2_2,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_0_2,
  output [7:0] O_9_1_0,
  output [7:0] O_9_1_1,
  output [7:0] O_9_1_2,
  output [7:0] O_9_2_0,
  output [7:0] O_9_2_1,
  output [7:0] O_9_2_2,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_0_2,
  output [7:0] O_10_1_0,
  output [7:0] O_10_1_1,
  output [7:0] O_10_1_2,
  output [7:0] O_10_2_0,
  output [7:0] O_10_2_1,
  output [7:0] O_10_2_2,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_0_2,
  output [7:0] O_11_1_0,
  output [7:0] O_11_1_1,
  output [7:0] O_11_1_2,
  output [7:0] O_11_2_0,
  output [7:0] O_11_2_1,
  output [7:0] O_11_2_2,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_0_2,
  output [7:0] O_12_1_0,
  output [7:0] O_12_1_1,
  output [7:0] O_12_1_2,
  output [7:0] O_12_2_0,
  output [7:0] O_12_2_1,
  output [7:0] O_12_2_2,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_0_2,
  output [7:0] O_13_1_0,
  output [7:0] O_13_1_1,
  output [7:0] O_13_1_2,
  output [7:0] O_13_2_0,
  output [7:0] O_13_2_1,
  output [7:0] O_13_2_2,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_0_2,
  output [7:0] O_14_1_0,
  output [7:0] O_14_1_1,
  output [7:0] O_14_1_2,
  output [7:0] O_14_2_0,
  output [7:0] O_14_2_1,
  output [7:0] O_14_2_2,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_0_2,
  output [7:0] O_15_1_0,
  output [7:0] O_15_1_1,
  output [7:0] O_15_1_2,
  output [7:0] O_15_2_0,
  output [7:0] O_15_2_1,
  output [7:0] O_15_2_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_2_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  Remove1S_3 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0_0(fst_op_I_0_0_0),
    .I_0_0_1(fst_op_I_0_0_1),
    .I_0_0_2(fst_op_I_0_0_2),
    .I_0_1_0(fst_op_I_0_1_0),
    .I_0_1_1(fst_op_I_0_1_1),
    .I_0_1_2(fst_op_I_0_1_2),
    .I_0_2_0(fst_op_I_0_2_0),
    .I_0_2_1(fst_op_I_0_2_1),
    .I_0_2_2(fst_op_I_0_2_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  Remove1S_3 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0_0(other_ops_0_I_0_0_0),
    .I_0_0_1(other_ops_0_I_0_0_1),
    .I_0_0_2(other_ops_0_I_0_0_2),
    .I_0_1_0(other_ops_0_I_0_1_0),
    .I_0_1_1(other_ops_0_I_0_1_1),
    .I_0_1_2(other_ops_0_I_0_1_2),
    .I_0_2_0(other_ops_0_I_0_2_0),
    .I_0_2_1(other_ops_0_I_0_2_1),
    .I_0_2_2(other_ops_0_I_0_2_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2),
    .O_2_0(other_ops_0_O_2_0),
    .O_2_1(other_ops_0_O_2_1),
    .O_2_2(other_ops_0_O_2_2)
  );
  Remove1S_3 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0_0(other_ops_1_I_0_0_0),
    .I_0_0_1(other_ops_1_I_0_0_1),
    .I_0_0_2(other_ops_1_I_0_0_2),
    .I_0_1_0(other_ops_1_I_0_1_0),
    .I_0_1_1(other_ops_1_I_0_1_1),
    .I_0_1_2(other_ops_1_I_0_1_2),
    .I_0_2_0(other_ops_1_I_0_2_0),
    .I_0_2_1(other_ops_1_I_0_2_1),
    .I_0_2_2(other_ops_1_I_0_2_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2),
    .O_2_0(other_ops_1_O_2_0),
    .O_2_1(other_ops_1_O_2_1),
    .O_2_2(other_ops_1_O_2_2)
  );
  Remove1S_3 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0_0(other_ops_2_I_0_0_0),
    .I_0_0_1(other_ops_2_I_0_0_1),
    .I_0_0_2(other_ops_2_I_0_0_2),
    .I_0_1_0(other_ops_2_I_0_1_0),
    .I_0_1_1(other_ops_2_I_0_1_1),
    .I_0_1_2(other_ops_2_I_0_1_2),
    .I_0_2_0(other_ops_2_I_0_2_0),
    .I_0_2_1(other_ops_2_I_0_2_1),
    .I_0_2_2(other_ops_2_I_0_2_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2),
    .O_2_0(other_ops_2_O_2_0),
    .O_2_1(other_ops_2_O_2_1),
    .O_2_2(other_ops_2_O_2_2)
  );
  Remove1S_3 other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0_0(other_ops_3_I_0_0_0),
    .I_0_0_1(other_ops_3_I_0_0_1),
    .I_0_0_2(other_ops_3_I_0_0_2),
    .I_0_1_0(other_ops_3_I_0_1_0),
    .I_0_1_1(other_ops_3_I_0_1_1),
    .I_0_1_2(other_ops_3_I_0_1_2),
    .I_0_2_0(other_ops_3_I_0_2_0),
    .I_0_2_1(other_ops_3_I_0_2_1),
    .I_0_2_2(other_ops_3_I_0_2_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2),
    .O_2_0(other_ops_3_O_2_0),
    .O_2_1(other_ops_3_O_2_1),
    .O_2_2(other_ops_3_O_2_2)
  );
  Remove1S_3 other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0_0(other_ops_4_I_0_0_0),
    .I_0_0_1(other_ops_4_I_0_0_1),
    .I_0_0_2(other_ops_4_I_0_0_2),
    .I_0_1_0(other_ops_4_I_0_1_0),
    .I_0_1_1(other_ops_4_I_0_1_1),
    .I_0_1_2(other_ops_4_I_0_1_2),
    .I_0_2_0(other_ops_4_I_0_2_0),
    .I_0_2_1(other_ops_4_I_0_2_1),
    .I_0_2_2(other_ops_4_I_0_2_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2),
    .O_2_0(other_ops_4_O_2_0),
    .O_2_1(other_ops_4_O_2_1),
    .O_2_2(other_ops_4_O_2_2)
  );
  Remove1S_3 other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0_0(other_ops_5_I_0_0_0),
    .I_0_0_1(other_ops_5_I_0_0_1),
    .I_0_0_2(other_ops_5_I_0_0_2),
    .I_0_1_0(other_ops_5_I_0_1_0),
    .I_0_1_1(other_ops_5_I_0_1_1),
    .I_0_1_2(other_ops_5_I_0_1_2),
    .I_0_2_0(other_ops_5_I_0_2_0),
    .I_0_2_1(other_ops_5_I_0_2_1),
    .I_0_2_2(other_ops_5_I_0_2_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2),
    .O_2_0(other_ops_5_O_2_0),
    .O_2_1(other_ops_5_O_2_1),
    .O_2_2(other_ops_5_O_2_2)
  );
  Remove1S_3 other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0_0(other_ops_6_I_0_0_0),
    .I_0_0_1(other_ops_6_I_0_0_1),
    .I_0_0_2(other_ops_6_I_0_0_2),
    .I_0_1_0(other_ops_6_I_0_1_0),
    .I_0_1_1(other_ops_6_I_0_1_1),
    .I_0_1_2(other_ops_6_I_0_1_2),
    .I_0_2_0(other_ops_6_I_0_2_0),
    .I_0_2_1(other_ops_6_I_0_2_1),
    .I_0_2_2(other_ops_6_I_0_2_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2),
    .O_2_0(other_ops_6_O_2_0),
    .O_2_1(other_ops_6_O_2_1),
    .O_2_2(other_ops_6_O_2_2)
  );
  Remove1S_3 other_ops_7 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I_0_0_0(other_ops_7_I_0_0_0),
    .I_0_0_1(other_ops_7_I_0_0_1),
    .I_0_0_2(other_ops_7_I_0_0_2),
    .I_0_1_0(other_ops_7_I_0_1_0),
    .I_0_1_1(other_ops_7_I_0_1_1),
    .I_0_1_2(other_ops_7_I_0_1_2),
    .I_0_2_0(other_ops_7_I_0_2_0),
    .I_0_2_1(other_ops_7_I_0_2_1),
    .I_0_2_2(other_ops_7_I_0_2_2),
    .O_0_0(other_ops_7_O_0_0),
    .O_0_1(other_ops_7_O_0_1),
    .O_0_2(other_ops_7_O_0_2),
    .O_1_0(other_ops_7_O_1_0),
    .O_1_1(other_ops_7_O_1_1),
    .O_1_2(other_ops_7_O_1_2),
    .O_2_0(other_ops_7_O_2_0),
    .O_2_1(other_ops_7_O_2_1),
    .O_2_2(other_ops_7_O_2_2)
  );
  Remove1S_3 other_ops_8 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I_0_0_0(other_ops_8_I_0_0_0),
    .I_0_0_1(other_ops_8_I_0_0_1),
    .I_0_0_2(other_ops_8_I_0_0_2),
    .I_0_1_0(other_ops_8_I_0_1_0),
    .I_0_1_1(other_ops_8_I_0_1_1),
    .I_0_1_2(other_ops_8_I_0_1_2),
    .I_0_2_0(other_ops_8_I_0_2_0),
    .I_0_2_1(other_ops_8_I_0_2_1),
    .I_0_2_2(other_ops_8_I_0_2_2),
    .O_0_0(other_ops_8_O_0_0),
    .O_0_1(other_ops_8_O_0_1),
    .O_0_2(other_ops_8_O_0_2),
    .O_1_0(other_ops_8_O_1_0),
    .O_1_1(other_ops_8_O_1_1),
    .O_1_2(other_ops_8_O_1_2),
    .O_2_0(other_ops_8_O_2_0),
    .O_2_1(other_ops_8_O_2_1),
    .O_2_2(other_ops_8_O_2_2)
  );
  Remove1S_3 other_ops_9 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I_0_0_0(other_ops_9_I_0_0_0),
    .I_0_0_1(other_ops_9_I_0_0_1),
    .I_0_0_2(other_ops_9_I_0_0_2),
    .I_0_1_0(other_ops_9_I_0_1_0),
    .I_0_1_1(other_ops_9_I_0_1_1),
    .I_0_1_2(other_ops_9_I_0_1_2),
    .I_0_2_0(other_ops_9_I_0_2_0),
    .I_0_2_1(other_ops_9_I_0_2_1),
    .I_0_2_2(other_ops_9_I_0_2_2),
    .O_0_0(other_ops_9_O_0_0),
    .O_0_1(other_ops_9_O_0_1),
    .O_0_2(other_ops_9_O_0_2),
    .O_1_0(other_ops_9_O_1_0),
    .O_1_1(other_ops_9_O_1_1),
    .O_1_2(other_ops_9_O_1_2),
    .O_2_0(other_ops_9_O_2_0),
    .O_2_1(other_ops_9_O_2_1),
    .O_2_2(other_ops_9_O_2_2)
  );
  Remove1S_3 other_ops_10 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I_0_0_0(other_ops_10_I_0_0_0),
    .I_0_0_1(other_ops_10_I_0_0_1),
    .I_0_0_2(other_ops_10_I_0_0_2),
    .I_0_1_0(other_ops_10_I_0_1_0),
    .I_0_1_1(other_ops_10_I_0_1_1),
    .I_0_1_2(other_ops_10_I_0_1_2),
    .I_0_2_0(other_ops_10_I_0_2_0),
    .I_0_2_1(other_ops_10_I_0_2_1),
    .I_0_2_2(other_ops_10_I_0_2_2),
    .O_0_0(other_ops_10_O_0_0),
    .O_0_1(other_ops_10_O_0_1),
    .O_0_2(other_ops_10_O_0_2),
    .O_1_0(other_ops_10_O_1_0),
    .O_1_1(other_ops_10_O_1_1),
    .O_1_2(other_ops_10_O_1_2),
    .O_2_0(other_ops_10_O_2_0),
    .O_2_1(other_ops_10_O_2_1),
    .O_2_2(other_ops_10_O_2_2)
  );
  Remove1S_3 other_ops_11 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I_0_0_0(other_ops_11_I_0_0_0),
    .I_0_0_1(other_ops_11_I_0_0_1),
    .I_0_0_2(other_ops_11_I_0_0_2),
    .I_0_1_0(other_ops_11_I_0_1_0),
    .I_0_1_1(other_ops_11_I_0_1_1),
    .I_0_1_2(other_ops_11_I_0_1_2),
    .I_0_2_0(other_ops_11_I_0_2_0),
    .I_0_2_1(other_ops_11_I_0_2_1),
    .I_0_2_2(other_ops_11_I_0_2_2),
    .O_0_0(other_ops_11_O_0_0),
    .O_0_1(other_ops_11_O_0_1),
    .O_0_2(other_ops_11_O_0_2),
    .O_1_0(other_ops_11_O_1_0),
    .O_1_1(other_ops_11_O_1_1),
    .O_1_2(other_ops_11_O_1_2),
    .O_2_0(other_ops_11_O_2_0),
    .O_2_1(other_ops_11_O_2_1),
    .O_2_2(other_ops_11_O_2_2)
  );
  Remove1S_3 other_ops_12 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I_0_0_0(other_ops_12_I_0_0_0),
    .I_0_0_1(other_ops_12_I_0_0_1),
    .I_0_0_2(other_ops_12_I_0_0_2),
    .I_0_1_0(other_ops_12_I_0_1_0),
    .I_0_1_1(other_ops_12_I_0_1_1),
    .I_0_1_2(other_ops_12_I_0_1_2),
    .I_0_2_0(other_ops_12_I_0_2_0),
    .I_0_2_1(other_ops_12_I_0_2_1),
    .I_0_2_2(other_ops_12_I_0_2_2),
    .O_0_0(other_ops_12_O_0_0),
    .O_0_1(other_ops_12_O_0_1),
    .O_0_2(other_ops_12_O_0_2),
    .O_1_0(other_ops_12_O_1_0),
    .O_1_1(other_ops_12_O_1_1),
    .O_1_2(other_ops_12_O_1_2),
    .O_2_0(other_ops_12_O_2_0),
    .O_2_1(other_ops_12_O_2_1),
    .O_2_2(other_ops_12_O_2_2)
  );
  Remove1S_3 other_ops_13 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I_0_0_0(other_ops_13_I_0_0_0),
    .I_0_0_1(other_ops_13_I_0_0_1),
    .I_0_0_2(other_ops_13_I_0_0_2),
    .I_0_1_0(other_ops_13_I_0_1_0),
    .I_0_1_1(other_ops_13_I_0_1_1),
    .I_0_1_2(other_ops_13_I_0_1_2),
    .I_0_2_0(other_ops_13_I_0_2_0),
    .I_0_2_1(other_ops_13_I_0_2_1),
    .I_0_2_2(other_ops_13_I_0_2_2),
    .O_0_0(other_ops_13_O_0_0),
    .O_0_1(other_ops_13_O_0_1),
    .O_0_2(other_ops_13_O_0_2),
    .O_1_0(other_ops_13_O_1_0),
    .O_1_1(other_ops_13_O_1_1),
    .O_1_2(other_ops_13_O_1_2),
    .O_2_0(other_ops_13_O_2_0),
    .O_2_1(other_ops_13_O_2_1),
    .O_2_2(other_ops_13_O_2_2)
  );
  Remove1S_3 other_ops_14 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I_0_0_0(other_ops_14_I_0_0_0),
    .I_0_0_1(other_ops_14_I_0_0_1),
    .I_0_0_2(other_ops_14_I_0_0_2),
    .I_0_1_0(other_ops_14_I_0_1_0),
    .I_0_1_1(other_ops_14_I_0_1_1),
    .I_0_1_2(other_ops_14_I_0_1_2),
    .I_0_2_0(other_ops_14_I_0_2_0),
    .I_0_2_1(other_ops_14_I_0_2_1),
    .I_0_2_2(other_ops_14_I_0_2_2),
    .O_0_0(other_ops_14_O_0_0),
    .O_0_1(other_ops_14_O_0_1),
    .O_0_2(other_ops_14_O_0_2),
    .O_1_0(other_ops_14_O_1_0),
    .O_1_1(other_ops_14_O_1_1),
    .O_1_2(other_ops_14_O_1_2),
    .O_2_0(other_ops_14_O_2_0),
    .O_2_1(other_ops_14_O_2_1),
    .O_2_2(other_ops_14_O_2_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[MapS.scala 17:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[MapS.scala 17:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[MapS.scala 17:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[MapS.scala 17:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[MapS.scala 17:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[MapS.scala 17:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[MapS.scala 17:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[MapS.scala 21:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[MapS.scala 21:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[MapS.scala 21:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[MapS.scala 21:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[MapS.scala 21:12]
  assign O_1_2_0 = other_ops_0_O_2_0; // @[MapS.scala 21:12]
  assign O_1_2_1 = other_ops_0_O_2_1; // @[MapS.scala 21:12]
  assign O_1_2_2 = other_ops_0_O_2_2; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[MapS.scala 21:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[MapS.scala 21:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[MapS.scala 21:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[MapS.scala 21:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[MapS.scala 21:12]
  assign O_2_2_0 = other_ops_1_O_2_0; // @[MapS.scala 21:12]
  assign O_2_2_1 = other_ops_1_O_2_1; // @[MapS.scala 21:12]
  assign O_2_2_2 = other_ops_1_O_2_2; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[MapS.scala 21:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[MapS.scala 21:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[MapS.scala 21:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[MapS.scala 21:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[MapS.scala 21:12]
  assign O_3_2_0 = other_ops_2_O_2_0; // @[MapS.scala 21:12]
  assign O_3_2_1 = other_ops_2_O_2_1; // @[MapS.scala 21:12]
  assign O_3_2_2 = other_ops_2_O_2_2; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[MapS.scala 21:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[MapS.scala 21:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[MapS.scala 21:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[MapS.scala 21:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[MapS.scala 21:12]
  assign O_4_2_0 = other_ops_3_O_2_0; // @[MapS.scala 21:12]
  assign O_4_2_1 = other_ops_3_O_2_1; // @[MapS.scala 21:12]
  assign O_4_2_2 = other_ops_3_O_2_2; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[MapS.scala 21:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[MapS.scala 21:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[MapS.scala 21:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[MapS.scala 21:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[MapS.scala 21:12]
  assign O_5_2_0 = other_ops_4_O_2_0; // @[MapS.scala 21:12]
  assign O_5_2_1 = other_ops_4_O_2_1; // @[MapS.scala 21:12]
  assign O_5_2_2 = other_ops_4_O_2_2; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[MapS.scala 21:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[MapS.scala 21:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[MapS.scala 21:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[MapS.scala 21:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[MapS.scala 21:12]
  assign O_6_2_0 = other_ops_5_O_2_0; // @[MapS.scala 21:12]
  assign O_6_2_1 = other_ops_5_O_2_1; // @[MapS.scala 21:12]
  assign O_6_2_2 = other_ops_5_O_2_2; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[MapS.scala 21:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[MapS.scala 21:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[MapS.scala 21:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[MapS.scala 21:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[MapS.scala 21:12]
  assign O_7_2_0 = other_ops_6_O_2_0; // @[MapS.scala 21:12]
  assign O_7_2_1 = other_ops_6_O_2_1; // @[MapS.scala 21:12]
  assign O_7_2_2 = other_ops_6_O_2_2; // @[MapS.scala 21:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[MapS.scala 21:12]
  assign O_8_0_1 = other_ops_7_O_0_1; // @[MapS.scala 21:12]
  assign O_8_0_2 = other_ops_7_O_0_2; // @[MapS.scala 21:12]
  assign O_8_1_0 = other_ops_7_O_1_0; // @[MapS.scala 21:12]
  assign O_8_1_1 = other_ops_7_O_1_1; // @[MapS.scala 21:12]
  assign O_8_1_2 = other_ops_7_O_1_2; // @[MapS.scala 21:12]
  assign O_8_2_0 = other_ops_7_O_2_0; // @[MapS.scala 21:12]
  assign O_8_2_1 = other_ops_7_O_2_1; // @[MapS.scala 21:12]
  assign O_8_2_2 = other_ops_7_O_2_2; // @[MapS.scala 21:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[MapS.scala 21:12]
  assign O_9_0_1 = other_ops_8_O_0_1; // @[MapS.scala 21:12]
  assign O_9_0_2 = other_ops_8_O_0_2; // @[MapS.scala 21:12]
  assign O_9_1_0 = other_ops_8_O_1_0; // @[MapS.scala 21:12]
  assign O_9_1_1 = other_ops_8_O_1_1; // @[MapS.scala 21:12]
  assign O_9_1_2 = other_ops_8_O_1_2; // @[MapS.scala 21:12]
  assign O_9_2_0 = other_ops_8_O_2_0; // @[MapS.scala 21:12]
  assign O_9_2_1 = other_ops_8_O_2_1; // @[MapS.scala 21:12]
  assign O_9_2_2 = other_ops_8_O_2_2; // @[MapS.scala 21:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[MapS.scala 21:12]
  assign O_10_0_1 = other_ops_9_O_0_1; // @[MapS.scala 21:12]
  assign O_10_0_2 = other_ops_9_O_0_2; // @[MapS.scala 21:12]
  assign O_10_1_0 = other_ops_9_O_1_0; // @[MapS.scala 21:12]
  assign O_10_1_1 = other_ops_9_O_1_1; // @[MapS.scala 21:12]
  assign O_10_1_2 = other_ops_9_O_1_2; // @[MapS.scala 21:12]
  assign O_10_2_0 = other_ops_9_O_2_0; // @[MapS.scala 21:12]
  assign O_10_2_1 = other_ops_9_O_2_1; // @[MapS.scala 21:12]
  assign O_10_2_2 = other_ops_9_O_2_2; // @[MapS.scala 21:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[MapS.scala 21:12]
  assign O_11_0_1 = other_ops_10_O_0_1; // @[MapS.scala 21:12]
  assign O_11_0_2 = other_ops_10_O_0_2; // @[MapS.scala 21:12]
  assign O_11_1_0 = other_ops_10_O_1_0; // @[MapS.scala 21:12]
  assign O_11_1_1 = other_ops_10_O_1_1; // @[MapS.scala 21:12]
  assign O_11_1_2 = other_ops_10_O_1_2; // @[MapS.scala 21:12]
  assign O_11_2_0 = other_ops_10_O_2_0; // @[MapS.scala 21:12]
  assign O_11_2_1 = other_ops_10_O_2_1; // @[MapS.scala 21:12]
  assign O_11_2_2 = other_ops_10_O_2_2; // @[MapS.scala 21:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[MapS.scala 21:12]
  assign O_12_0_1 = other_ops_11_O_0_1; // @[MapS.scala 21:12]
  assign O_12_0_2 = other_ops_11_O_0_2; // @[MapS.scala 21:12]
  assign O_12_1_0 = other_ops_11_O_1_0; // @[MapS.scala 21:12]
  assign O_12_1_1 = other_ops_11_O_1_1; // @[MapS.scala 21:12]
  assign O_12_1_2 = other_ops_11_O_1_2; // @[MapS.scala 21:12]
  assign O_12_2_0 = other_ops_11_O_2_0; // @[MapS.scala 21:12]
  assign O_12_2_1 = other_ops_11_O_2_1; // @[MapS.scala 21:12]
  assign O_12_2_2 = other_ops_11_O_2_2; // @[MapS.scala 21:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[MapS.scala 21:12]
  assign O_13_0_1 = other_ops_12_O_0_1; // @[MapS.scala 21:12]
  assign O_13_0_2 = other_ops_12_O_0_2; // @[MapS.scala 21:12]
  assign O_13_1_0 = other_ops_12_O_1_0; // @[MapS.scala 21:12]
  assign O_13_1_1 = other_ops_12_O_1_1; // @[MapS.scala 21:12]
  assign O_13_1_2 = other_ops_12_O_1_2; // @[MapS.scala 21:12]
  assign O_13_2_0 = other_ops_12_O_2_0; // @[MapS.scala 21:12]
  assign O_13_2_1 = other_ops_12_O_2_1; // @[MapS.scala 21:12]
  assign O_13_2_2 = other_ops_12_O_2_2; // @[MapS.scala 21:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[MapS.scala 21:12]
  assign O_14_0_1 = other_ops_13_O_0_1; // @[MapS.scala 21:12]
  assign O_14_0_2 = other_ops_13_O_0_2; // @[MapS.scala 21:12]
  assign O_14_1_0 = other_ops_13_O_1_0; // @[MapS.scala 21:12]
  assign O_14_1_1 = other_ops_13_O_1_1; // @[MapS.scala 21:12]
  assign O_14_1_2 = other_ops_13_O_1_2; // @[MapS.scala 21:12]
  assign O_14_2_0 = other_ops_13_O_2_0; // @[MapS.scala 21:12]
  assign O_14_2_1 = other_ops_13_O_2_1; // @[MapS.scala 21:12]
  assign O_14_2_2 = other_ops_13_O_2_2; // @[MapS.scala 21:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[MapS.scala 21:12]
  assign O_15_0_1 = other_ops_14_O_0_1; // @[MapS.scala 21:12]
  assign O_15_0_2 = other_ops_14_O_0_2; // @[MapS.scala 21:12]
  assign O_15_1_0 = other_ops_14_O_1_0; // @[MapS.scala 21:12]
  assign O_15_1_1 = other_ops_14_O_1_1; // @[MapS.scala 21:12]
  assign O_15_1_2 = other_ops_14_O_1_2; // @[MapS.scala 21:12]
  assign O_15_2_0 = other_ops_14_O_2_0; // @[MapS.scala 21:12]
  assign O_15_2_1 = other_ops_14_O_2_1; // @[MapS.scala 21:12]
  assign O_15_2_2 = other_ops_14_O_2_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0_0 = I_0_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_1 = I_0_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_2 = I_0_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_0 = I_0_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_1 = I_0_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_2 = I_0_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_0 = I_0_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_1 = I_0_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_2 = I_0_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0_0 = I_1_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_1 = I_1_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_2 = I_1_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_0 = I_1_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_1 = I_1_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_2 = I_1_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_0 = I_1_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_1 = I_1_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_2 = I_1_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0_0 = I_2_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_1 = I_2_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_2 = I_2_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_0 = I_2_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_1 = I_2_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_2 = I_2_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_0 = I_2_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_1 = I_2_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_2 = I_2_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0_0 = I_3_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_1 = I_3_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_2 = I_3_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_0 = I_3_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_1 = I_3_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_2 = I_3_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_0 = I_3_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_1 = I_3_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_2 = I_3_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0_0 = I_4_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_1 = I_4_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_2 = I_4_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_0 = I_4_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_1 = I_4_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_2 = I_4_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_0 = I_4_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_1 = I_4_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_2 = I_4_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0_0 = I_5_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_1 = I_5_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_2 = I_5_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_0 = I_5_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_1 = I_5_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_2 = I_5_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_0 = I_5_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_1 = I_5_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_2 = I_5_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0_0 = I_6_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_1 = I_6_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_2 = I_6_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_0 = I_6_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_1 = I_6_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_2 = I_6_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_0 = I_6_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_1 = I_6_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_2 = I_6_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0_0 = I_7_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_1 = I_7_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_2 = I_7_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_0 = I_7_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_1 = I_7_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_2 = I_7_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_0 = I_7_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_1 = I_7_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_2 = I_7_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I_0_0_0 = I_8_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_0_1 = I_8_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_0_2 = I_8_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1_0 = I_8_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1_1 = I_8_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1_2 = I_8_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2_0 = I_8_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2_1 = I_8_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2_2 = I_8_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I_0_0_0 = I_9_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_0_1 = I_9_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_0_2 = I_9_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1_0 = I_9_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1_1 = I_9_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1_2 = I_9_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2_0 = I_9_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2_1 = I_9_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2_2 = I_9_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I_0_0_0 = I_10_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_0_1 = I_10_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_0_2 = I_10_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1_0 = I_10_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1_1 = I_10_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1_2 = I_10_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2_0 = I_10_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2_1 = I_10_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2_2 = I_10_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I_0_0_0 = I_11_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_0_1 = I_11_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_0_2 = I_11_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1_0 = I_11_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1_1 = I_11_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1_2 = I_11_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2_0 = I_11_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2_1 = I_11_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2_2 = I_11_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I_0_0_0 = I_12_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_0_1 = I_12_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_0_2 = I_12_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1_0 = I_12_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1_1 = I_12_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1_2 = I_12_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2_0 = I_12_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2_1 = I_12_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2_2 = I_12_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I_0_0_0 = I_13_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_0_1 = I_13_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_0_2 = I_13_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1_0 = I_13_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1_1 = I_13_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1_2 = I_13_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2_0 = I_13_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2_1 = I_13_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2_2 = I_13_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I_0_0_0 = I_14_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_0_1 = I_14_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_0_2 = I_14_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1_0 = I_14_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1_1 = I_14_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1_2 = I_14_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2_0 = I_14_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2_1 = I_14_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2_2 = I_14_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I_0_0_0 = I_15_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_0_1 = I_15_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_0_2 = I_15_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1_0 = I_15_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1_1 = I_15_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1_2 = I_15_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2_0 = I_15_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2_1 = I_15_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2_2 = I_15_0_2_2; // @[MapS.scala 20:41]
endmodule
module InitialDelayCounter(
  input   clock,
  input   reset,
  output  valid_down
);
  reg  value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire  _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 1'h1; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 1'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 1'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module AtomTuple(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  input  [7:0] I1,
  output [7:0] O_t0b,
  output [7:0] O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b = I1; // @[Tuple.scala 50:9]
endmodule
module Map2S_8(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I0_2,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  output [7:0] O_0_t0b,
  output [7:0] O_0_t1b,
  output [7:0] O_1_t0b,
  output [7:0] O_1_t1b,
  output [7:0] O_2_t0b,
  output [7:0] O_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  AtomTuple other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_t0b(other_ops_0_O_t0b),
    .O_t1b(other_ops_0_O_t1b)
  );
  AtomTuple other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_t0b(other_ops_1_O_t0b),
    .O_t1b(other_ops_1_O_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign O_1_t0b = other_ops_0_O_t0b; // @[Map2S.scala 24:12]
  assign O_1_t1b = other_ops_0_O_t1b; // @[Map2S.scala 24:12]
  assign O_2_t0b = other_ops_1_O_t0b; // @[Map2S.scala 24:12]
  assign O_2_t1b = other_ops_1_O_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
endmodule
module Map2S_9(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_0_2,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_1_2,
  input  [7:0] I0_2_0,
  input  [7:0] I0_2_1,
  input  [7:0] I0_2_2,
  output [7:0] O_0_0_t0b,
  output [7:0] O_0_0_t1b,
  output [7:0] O_0_1_t0b,
  output [7:0] O_0_1_t1b,
  output [7:0] O_0_2_t0b,
  output [7:0] O_0_2_t1b,
  output [7:0] O_1_0_t0b,
  output [7:0] O_1_0_t1b,
  output [7:0] O_1_1_t0b,
  output [7:0] O_1_1_t1b,
  output [7:0] O_1_2_t0b,
  output [7:0] O_1_2_t1b,
  output [7:0] O_2_0_t0b,
  output [7:0] O_2_0_t1b,
  output [7:0] O_2_1_t0b,
  output [7:0] O_2_1_t1b,
  output [7:0] O_2_2_t0b,
  output [7:0] O_2_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_t1b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  Map2S_8 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b),
    .O_1_t0b(fst_op_O_1_t0b),
    .O_1_t1b(fst_op_O_1_t1b),
    .O_2_t0b(fst_op_O_2_t0b),
    .O_2_t1b(fst_op_O_2_t1b)
  );
  Map2S_8 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I0_2(other_ops_0_I0_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_t0b(other_ops_0_O_0_t0b),
    .O_0_t1b(other_ops_0_O_0_t1b),
    .O_1_t0b(other_ops_0_O_1_t0b),
    .O_1_t1b(other_ops_0_O_1_t1b),
    .O_2_t0b(other_ops_0_O_2_t0b),
    .O_2_t1b(other_ops_0_O_2_t1b)
  );
  Map2S_8 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I0_2(other_ops_1_I0_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_t0b(other_ops_1_O_0_t0b),
    .O_0_t1b(other_ops_1_O_0_t1b),
    .O_1_t0b(other_ops_1_O_1_t0b),
    .O_1_t1b(other_ops_1_O_1_t1b),
    .O_2_t0b(other_ops_1_O_2_t0b),
    .O_2_t1b(other_ops_1_O_2_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign O_0_1_t0b = fst_op_O_1_t0b; // @[Map2S.scala 19:8]
  assign O_0_1_t1b = fst_op_O_1_t1b; // @[Map2S.scala 19:8]
  assign O_0_2_t0b = fst_op_O_2_t0b; // @[Map2S.scala 19:8]
  assign O_0_2_t1b = fst_op_O_2_t1b; // @[Map2S.scala 19:8]
  assign O_1_0_t0b = other_ops_0_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_1_0_t1b = other_ops_0_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_1_1_t0b = other_ops_0_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_1_1_t1b = other_ops_0_O_1_t1b; // @[Map2S.scala 24:12]
  assign O_1_2_t0b = other_ops_0_O_2_t0b; // @[Map2S.scala 24:12]
  assign O_1_2_t1b = other_ops_0_O_2_t1b; // @[Map2S.scala 24:12]
  assign O_2_0_t0b = other_ops_1_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_2_0_t1b = other_ops_1_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_2_1_t0b = other_ops_1_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_2_1_t1b = other_ops_1_O_1_t1b; // @[Map2S.scala 24:12]
  assign O_2_2_t0b = other_ops_1_O_2_t0b; // @[Map2S.scala 24:12]
  assign O_2_2_t1b = other_ops_1_O_2_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = 8'h0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = 8'h1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = 8'h0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2 = I0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = 8'h1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = 8'h2; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = 8'h1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2 = I0_2_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = 8'h0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = 8'h1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = 8'h0; // @[Map2S.scala 23:43]
endmodule
module LShift(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  wire [262:0] _GEN_0; // @[Arithmetic.scala 301:25]
  wire [262:0] _T; // @[Arithmetic.scala 301:25]
  assign _GEN_0 = {{255'd0}, I_t0b}; // @[Arithmetic.scala 301:25]
  assign _T = _GEN_0 << I_t1b; // @[Arithmetic.scala 301:25]
  assign valid_down = valid_up; // @[Arithmetic.scala 303:14]
  assign O = _T[7:0]; // @[Arithmetic.scala 301:7]
endmodule
module MapS_4(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  input  [7:0] I_1_t0b,
  input  [7:0] I_1_t1b,
  input  [7:0] I_2_t0b,
  input  [7:0] I_2_t1b,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  LShift fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  LShift other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_t0b(other_ops_0_I_t0b),
    .I_t1b(other_ops_0_I_t1b),
    .O(other_ops_0_O)
  );
  LShift other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_t0b(other_ops_1_I_t0b),
    .I_t1b(other_ops_1_I_t1b),
    .O(other_ops_1_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_t0b = I_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_t1b = I_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_t0b = I_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_t1b = I_2_t1b; // @[MapS.scala 20:41]
endmodule
module MapS_5(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_t0b,
  input  [7:0] I_0_0_t1b,
  input  [7:0] I_0_1_t0b,
  input  [7:0] I_0_1_t1b,
  input  [7:0] I_0_2_t0b,
  input  [7:0] I_0_2_t1b,
  input  [7:0] I_1_0_t0b,
  input  [7:0] I_1_0_t1b,
  input  [7:0] I_1_1_t0b,
  input  [7:0] I_1_1_t1b,
  input  [7:0] I_1_2_t0b,
  input  [7:0] I_1_2_t1b,
  input  [7:0] I_2_0_t0b,
  input  [7:0] I_2_0_t1b,
  input  [7:0] I_2_1_t0b,
  input  [7:0] I_2_1_t1b,
  input  [7:0] I_2_2_t0b,
  input  [7:0] I_2_2_t1b,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  MapS_4 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .I_1_t0b(fst_op_I_1_t0b),
    .I_1_t1b(fst_op_I_1_t1b),
    .I_2_t0b(fst_op_I_2_t0b),
    .I_2_t1b(fst_op_I_2_t1b),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  MapS_4 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_t0b(other_ops_0_I_0_t0b),
    .I_0_t1b(other_ops_0_I_0_t1b),
    .I_1_t0b(other_ops_0_I_1_t0b),
    .I_1_t1b(other_ops_0_I_1_t1b),
    .I_2_t0b(other_ops_0_I_2_t0b),
    .I_2_t1b(other_ops_0_I_2_t1b),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  MapS_4 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_t0b(other_ops_1_I_0_t0b),
    .I_0_t1b(other_ops_1_I_0_t1b),
    .I_1_t0b(other_ops_1_I_1_t0b),
    .I_1_t1b(other_ops_1_I_1_t1b),
    .I_2_t0b(other_ops_1_I_2_t0b),
    .I_2_t1b(other_ops_1_I_2_t1b),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_1_2 = other_ops_0_O_2; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign O_2_1 = other_ops_1_O_1; // @[MapS.scala 21:12]
  assign O_2_2 = other_ops_1_O_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t0b = I_0_1_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t1b = I_0_1_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_2_t0b = I_0_2_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_2_t1b = I_0_2_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_t0b = I_1_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_t1b = I_1_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t0b = I_1_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t1b = I_1_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_t0b = I_1_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_t1b = I_1_2_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_t0b = I_2_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_t1b = I_2_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_t0b = I_2_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_t1b = I_2_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_t0b = I_2_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_t1b = I_2_2_t1b; // @[MapS.scala 20:41]
endmodule
module AddNoValid(
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  assign O = I_t0b + I_t1b; // @[Arithmetic.scala 122:7]
endmodule
module ReduceS(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  output [7:0] O_0
);
  wire [7:0] AddNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_O; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_1_I_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_1_I_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_1_O; // @[ReduceS.scala 20:43]
  reg [7:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_1;
  AddNoValid AddNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  AddNoValid AddNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_1_I_t0b),
    .I_t1b(AddNoValid_1_I_t1b),
    .O(AddNoValid_1_O)
  );
  assign valid_down = _T_1; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign AddNoValid_I_t0b = I_0; // @[ReduceS.scala 43:18]
  assign AddNoValid_I_t1b = AddNoValid_1_O; // @[ReduceS.scala 36:18]
  assign AddNoValid_1_I_t0b = I_1; // @[ReduceS.scala 43:18]
  assign AddNoValid_1_I_t1b = I_2; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= AddNoValid_O;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module MapS_6(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_2_2,
  output [7:0] O_0_0,
  output [7:0] O_1_0,
  output [7:0] O_2_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  ReduceS fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .I_2(fst_op_I_2),
    .O_0(fst_op_O_0)
  );
  ReduceS other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0(other_ops_0_I_0),
    .I_1(other_ops_0_I_1),
    .I_2(other_ops_0_I_2),
    .O_0(other_ops_0_O_0)
  );
  ReduceS other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0(other_ops_1_I_0),
    .I_1(other_ops_1_I_1),
    .I_2(other_ops_1_I_2),
    .O_0(other_ops_1_O_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_2 = I_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0 = I_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1 = I_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2 = I_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0 = I_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1 = I_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2 = I_2_2; // @[MapS.scala 20:41]
endmodule
module MapSNoValid(
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  output [7:0] O_0
);
  wire [7:0] fst_op_I_t0b; // @[MapS.scala 28:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 28:22]
  wire [7:0] fst_op_O; // @[MapS.scala 28:22]
  AddNoValid fst_op ( // @[MapS.scala 28:22]
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign O_0 = fst_op_O; // @[MapS.scala 35:8]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 34:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 34:12]
endmodule
module ReduceS_1(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_1_0,
  input  [7:0] I_2_0,
  output [7:0] O_0_0
);
  wire [7:0] MapSNoValid_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_O_0; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_1_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_1_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_1_O_0; // @[ReduceS.scala 20:43]
  reg [7:0] _T_0; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_1;
  MapSNoValid MapSNoValid ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_I_0_t0b),
    .I_0_t1b(MapSNoValid_I_0_t1b),
    .O_0(MapSNoValid_O_0)
  );
  MapSNoValid MapSNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_1_I_0_t0b),
    .I_0_t1b(MapSNoValid_1_I_0_t1b),
    .O_0(MapSNoValid_1_O_0)
  );
  assign valid_down = _T_1; // @[ReduceS.scala 47:14]
  assign O_0_0 = _T_0; // @[ReduceS.scala 27:14]
  assign MapSNoValid_I_0_t0b = I_1_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_I_0_t1b = MapSNoValid_1_O_0; // @[ReduceS.scala 36:18]
  assign MapSNoValid_1_I_0_t0b = I_0_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_1_I_0_t1b = I_2_0; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0 <= MapSNoValid_O_0;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module InitialDelayCounter_1(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [1:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [1:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 2'h3; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 2'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 2'h3; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 2'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module Map2S_10(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  output [7:0] O_0_t0b,
  output [7:0] O_0_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = 8'h4; // @[Map2S.scala 18:13]
endmodule
module Map2S_11(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  output [7:0] O_0_0_t0b,
  output [7:0] O_0_0_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  Map2S_10 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
endmodule
module RShift(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 272:14]
  assign O = I_t0b >> I_t1b; // @[Arithmetic.scala 270:7]
endmodule
module MapS_7(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  output [7:0] O_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  RShift fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
endmodule
module MapS_8(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_t0b,
  input  [7:0] I_0_0_t1b,
  output [7:0] O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  MapS_7 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
endmodule
module Module_0(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_2_2,
  output [7:0] O_0_0
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n69_valid_up; // @[Top.scala 16:21]
  wire  n69_valid_down; // @[Top.scala 16:21]
  wire [7:0] n69_I0_0_0; // @[Top.scala 16:21]
  wire [7:0] n69_I0_0_1; // @[Top.scala 16:21]
  wire [7:0] n69_I0_0_2; // @[Top.scala 16:21]
  wire [7:0] n69_I0_1_0; // @[Top.scala 16:21]
  wire [7:0] n69_I0_1_1; // @[Top.scala 16:21]
  wire [7:0] n69_I0_1_2; // @[Top.scala 16:21]
  wire [7:0] n69_I0_2_0; // @[Top.scala 16:21]
  wire [7:0] n69_I0_2_1; // @[Top.scala 16:21]
  wire [7:0] n69_I0_2_2; // @[Top.scala 16:21]
  wire [7:0] n69_O_0_0_t0b; // @[Top.scala 16:21]
  wire [7:0] n69_O_0_0_t1b; // @[Top.scala 16:21]
  wire [7:0] n69_O_0_1_t0b; // @[Top.scala 16:21]
  wire [7:0] n69_O_0_1_t1b; // @[Top.scala 16:21]
  wire [7:0] n69_O_0_2_t0b; // @[Top.scala 16:21]
  wire [7:0] n69_O_0_2_t1b; // @[Top.scala 16:21]
  wire [7:0] n69_O_1_0_t0b; // @[Top.scala 16:21]
  wire [7:0] n69_O_1_0_t1b; // @[Top.scala 16:21]
  wire [7:0] n69_O_1_1_t0b; // @[Top.scala 16:21]
  wire [7:0] n69_O_1_1_t1b; // @[Top.scala 16:21]
  wire [7:0] n69_O_1_2_t0b; // @[Top.scala 16:21]
  wire [7:0] n69_O_1_2_t1b; // @[Top.scala 16:21]
  wire [7:0] n69_O_2_0_t0b; // @[Top.scala 16:21]
  wire [7:0] n69_O_2_0_t1b; // @[Top.scala 16:21]
  wire [7:0] n69_O_2_1_t0b; // @[Top.scala 16:21]
  wire [7:0] n69_O_2_1_t1b; // @[Top.scala 16:21]
  wire [7:0] n69_O_2_2_t0b; // @[Top.scala 16:21]
  wire [7:0] n69_O_2_2_t1b; // @[Top.scala 16:21]
  wire  n80_valid_up; // @[Top.scala 20:21]
  wire  n80_valid_down; // @[Top.scala 20:21]
  wire [7:0] n80_I_0_0_t0b; // @[Top.scala 20:21]
  wire [7:0] n80_I_0_0_t1b; // @[Top.scala 20:21]
  wire [7:0] n80_I_0_1_t0b; // @[Top.scala 20:21]
  wire [7:0] n80_I_0_1_t1b; // @[Top.scala 20:21]
  wire [7:0] n80_I_0_2_t0b; // @[Top.scala 20:21]
  wire [7:0] n80_I_0_2_t1b; // @[Top.scala 20:21]
  wire [7:0] n80_I_1_0_t0b; // @[Top.scala 20:21]
  wire [7:0] n80_I_1_0_t1b; // @[Top.scala 20:21]
  wire [7:0] n80_I_1_1_t0b; // @[Top.scala 20:21]
  wire [7:0] n80_I_1_1_t1b; // @[Top.scala 20:21]
  wire [7:0] n80_I_1_2_t0b; // @[Top.scala 20:21]
  wire [7:0] n80_I_1_2_t1b; // @[Top.scala 20:21]
  wire [7:0] n80_I_2_0_t0b; // @[Top.scala 20:21]
  wire [7:0] n80_I_2_0_t1b; // @[Top.scala 20:21]
  wire [7:0] n80_I_2_1_t0b; // @[Top.scala 20:21]
  wire [7:0] n80_I_2_1_t1b; // @[Top.scala 20:21]
  wire [7:0] n80_I_2_2_t0b; // @[Top.scala 20:21]
  wire [7:0] n80_I_2_2_t1b; // @[Top.scala 20:21]
  wire [7:0] n80_O_0_0; // @[Top.scala 20:21]
  wire [7:0] n80_O_0_1; // @[Top.scala 20:21]
  wire [7:0] n80_O_0_2; // @[Top.scala 20:21]
  wire [7:0] n80_O_1_0; // @[Top.scala 20:21]
  wire [7:0] n80_O_1_1; // @[Top.scala 20:21]
  wire [7:0] n80_O_1_2; // @[Top.scala 20:21]
  wire [7:0] n80_O_2_0; // @[Top.scala 20:21]
  wire [7:0] n80_O_2_1; // @[Top.scala 20:21]
  wire [7:0] n80_O_2_2; // @[Top.scala 20:21]
  wire  n85_clock; // @[Top.scala 23:21]
  wire  n85_reset; // @[Top.scala 23:21]
  wire  n85_valid_up; // @[Top.scala 23:21]
  wire  n85_valid_down; // @[Top.scala 23:21]
  wire [7:0] n85_I_0_0; // @[Top.scala 23:21]
  wire [7:0] n85_I_0_1; // @[Top.scala 23:21]
  wire [7:0] n85_I_0_2; // @[Top.scala 23:21]
  wire [7:0] n85_I_1_0; // @[Top.scala 23:21]
  wire [7:0] n85_I_1_1; // @[Top.scala 23:21]
  wire [7:0] n85_I_1_2; // @[Top.scala 23:21]
  wire [7:0] n85_I_2_0; // @[Top.scala 23:21]
  wire [7:0] n85_I_2_1; // @[Top.scala 23:21]
  wire [7:0] n85_I_2_2; // @[Top.scala 23:21]
  wire [7:0] n85_O_0_0; // @[Top.scala 23:21]
  wire [7:0] n85_O_1_0; // @[Top.scala 23:21]
  wire [7:0] n85_O_2_0; // @[Top.scala 23:21]
  wire  n90_clock; // @[Top.scala 26:21]
  wire  n90_reset; // @[Top.scala 26:21]
  wire  n90_valid_up; // @[Top.scala 26:21]
  wire  n90_valid_down; // @[Top.scala 26:21]
  wire [7:0] n90_I_0_0; // @[Top.scala 26:21]
  wire [7:0] n90_I_1_0; // @[Top.scala 26:21]
  wire [7:0] n90_I_2_0; // @[Top.scala 26:21]
  wire [7:0] n90_O_0_0; // @[Top.scala 26:21]
  wire  InitialDelayCounter_1_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_valid_down; // @[Const.scala 11:33]
  wire  n93_valid_up; // @[Top.scala 30:21]
  wire  n93_valid_down; // @[Top.scala 30:21]
  wire [7:0] n93_I0_0_0; // @[Top.scala 30:21]
  wire [7:0] n93_O_0_0_t0b; // @[Top.scala 30:21]
  wire [7:0] n93_O_0_0_t1b; // @[Top.scala 30:21]
  wire  n104_valid_up; // @[Top.scala 34:22]
  wire  n104_valid_down; // @[Top.scala 34:22]
  wire [7:0] n104_I_0_0_t0b; // @[Top.scala 34:22]
  wire [7:0] n104_I_0_0_t1b; // @[Top.scala 34:22]
  wire [7:0] n104_O_0_0; // @[Top.scala 34:22]
  InitialDelayCounter InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  Map2S_9 n69 ( // @[Top.scala 16:21]
    .valid_up(n69_valid_up),
    .valid_down(n69_valid_down),
    .I0_0_0(n69_I0_0_0),
    .I0_0_1(n69_I0_0_1),
    .I0_0_2(n69_I0_0_2),
    .I0_1_0(n69_I0_1_0),
    .I0_1_1(n69_I0_1_1),
    .I0_1_2(n69_I0_1_2),
    .I0_2_0(n69_I0_2_0),
    .I0_2_1(n69_I0_2_1),
    .I0_2_2(n69_I0_2_2),
    .O_0_0_t0b(n69_O_0_0_t0b),
    .O_0_0_t1b(n69_O_0_0_t1b),
    .O_0_1_t0b(n69_O_0_1_t0b),
    .O_0_1_t1b(n69_O_0_1_t1b),
    .O_0_2_t0b(n69_O_0_2_t0b),
    .O_0_2_t1b(n69_O_0_2_t1b),
    .O_1_0_t0b(n69_O_1_0_t0b),
    .O_1_0_t1b(n69_O_1_0_t1b),
    .O_1_1_t0b(n69_O_1_1_t0b),
    .O_1_1_t1b(n69_O_1_1_t1b),
    .O_1_2_t0b(n69_O_1_2_t0b),
    .O_1_2_t1b(n69_O_1_2_t1b),
    .O_2_0_t0b(n69_O_2_0_t0b),
    .O_2_0_t1b(n69_O_2_0_t1b),
    .O_2_1_t0b(n69_O_2_1_t0b),
    .O_2_1_t1b(n69_O_2_1_t1b),
    .O_2_2_t0b(n69_O_2_2_t0b),
    .O_2_2_t1b(n69_O_2_2_t1b)
  );
  MapS_5 n80 ( // @[Top.scala 20:21]
    .valid_up(n80_valid_up),
    .valid_down(n80_valid_down),
    .I_0_0_t0b(n80_I_0_0_t0b),
    .I_0_0_t1b(n80_I_0_0_t1b),
    .I_0_1_t0b(n80_I_0_1_t0b),
    .I_0_1_t1b(n80_I_0_1_t1b),
    .I_0_2_t0b(n80_I_0_2_t0b),
    .I_0_2_t1b(n80_I_0_2_t1b),
    .I_1_0_t0b(n80_I_1_0_t0b),
    .I_1_0_t1b(n80_I_1_0_t1b),
    .I_1_1_t0b(n80_I_1_1_t0b),
    .I_1_1_t1b(n80_I_1_1_t1b),
    .I_1_2_t0b(n80_I_1_2_t0b),
    .I_1_2_t1b(n80_I_1_2_t1b),
    .I_2_0_t0b(n80_I_2_0_t0b),
    .I_2_0_t1b(n80_I_2_0_t1b),
    .I_2_1_t0b(n80_I_2_1_t0b),
    .I_2_1_t1b(n80_I_2_1_t1b),
    .I_2_2_t0b(n80_I_2_2_t0b),
    .I_2_2_t1b(n80_I_2_2_t1b),
    .O_0_0(n80_O_0_0),
    .O_0_1(n80_O_0_1),
    .O_0_2(n80_O_0_2),
    .O_1_0(n80_O_1_0),
    .O_1_1(n80_O_1_1),
    .O_1_2(n80_O_1_2),
    .O_2_0(n80_O_2_0),
    .O_2_1(n80_O_2_1),
    .O_2_2(n80_O_2_2)
  );
  MapS_6 n85 ( // @[Top.scala 23:21]
    .clock(n85_clock),
    .reset(n85_reset),
    .valid_up(n85_valid_up),
    .valid_down(n85_valid_down),
    .I_0_0(n85_I_0_0),
    .I_0_1(n85_I_0_1),
    .I_0_2(n85_I_0_2),
    .I_1_0(n85_I_1_0),
    .I_1_1(n85_I_1_1),
    .I_1_2(n85_I_1_2),
    .I_2_0(n85_I_2_0),
    .I_2_1(n85_I_2_1),
    .I_2_2(n85_I_2_2),
    .O_0_0(n85_O_0_0),
    .O_1_0(n85_O_1_0),
    .O_2_0(n85_O_2_0)
  );
  ReduceS_1 n90 ( // @[Top.scala 26:21]
    .clock(n90_clock),
    .reset(n90_reset),
    .valid_up(n90_valid_up),
    .valid_down(n90_valid_down),
    .I_0_0(n90_I_0_0),
    .I_1_0(n90_I_1_0),
    .I_2_0(n90_I_2_0),
    .O_0_0(n90_O_0_0)
  );
  InitialDelayCounter_1 InitialDelayCounter_1 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_1_clock),
    .reset(InitialDelayCounter_1_reset),
    .valid_down(InitialDelayCounter_1_valid_down)
  );
  Map2S_11 n93 ( // @[Top.scala 30:21]
    .valid_up(n93_valid_up),
    .valid_down(n93_valid_down),
    .I0_0_0(n93_I0_0_0),
    .O_0_0_t0b(n93_O_0_0_t0b),
    .O_0_0_t1b(n93_O_0_0_t1b)
  );
  MapS_8 n104 ( // @[Top.scala 34:22]
    .valid_up(n104_valid_up),
    .valid_down(n104_valid_down),
    .I_0_0_t0b(n104_I_0_0_t0b),
    .I_0_0_t1b(n104_I_0_0_t1b),
    .O_0_0(n104_O_0_0)
  );
  assign valid_down = n104_valid_down; // @[Top.scala 38:16]
  assign O_0_0 = n104_O_0_0; // @[Top.scala 37:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n69_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 19:18]
  assign n69_I0_0_0 = I_0_0; // @[Top.scala 17:12]
  assign n69_I0_0_1 = I_0_1; // @[Top.scala 17:12]
  assign n69_I0_0_2 = I_0_2; // @[Top.scala 17:12]
  assign n69_I0_1_0 = I_1_0; // @[Top.scala 17:12]
  assign n69_I0_1_1 = I_1_1; // @[Top.scala 17:12]
  assign n69_I0_1_2 = I_1_2; // @[Top.scala 17:12]
  assign n69_I0_2_0 = I_2_0; // @[Top.scala 17:12]
  assign n69_I0_2_1 = I_2_1; // @[Top.scala 17:12]
  assign n69_I0_2_2 = I_2_2; // @[Top.scala 17:12]
  assign n80_valid_up = n69_valid_down; // @[Top.scala 22:18]
  assign n80_I_0_0_t0b = n69_O_0_0_t0b; // @[Top.scala 21:11]
  assign n80_I_0_0_t1b = n69_O_0_0_t1b; // @[Top.scala 21:11]
  assign n80_I_0_1_t0b = n69_O_0_1_t0b; // @[Top.scala 21:11]
  assign n80_I_0_1_t1b = n69_O_0_1_t1b; // @[Top.scala 21:11]
  assign n80_I_0_2_t0b = n69_O_0_2_t0b; // @[Top.scala 21:11]
  assign n80_I_0_2_t1b = n69_O_0_2_t1b; // @[Top.scala 21:11]
  assign n80_I_1_0_t0b = n69_O_1_0_t0b; // @[Top.scala 21:11]
  assign n80_I_1_0_t1b = n69_O_1_0_t1b; // @[Top.scala 21:11]
  assign n80_I_1_1_t0b = n69_O_1_1_t0b; // @[Top.scala 21:11]
  assign n80_I_1_1_t1b = n69_O_1_1_t1b; // @[Top.scala 21:11]
  assign n80_I_1_2_t0b = n69_O_1_2_t0b; // @[Top.scala 21:11]
  assign n80_I_1_2_t1b = n69_O_1_2_t1b; // @[Top.scala 21:11]
  assign n80_I_2_0_t0b = n69_O_2_0_t0b; // @[Top.scala 21:11]
  assign n80_I_2_0_t1b = n69_O_2_0_t1b; // @[Top.scala 21:11]
  assign n80_I_2_1_t0b = n69_O_2_1_t0b; // @[Top.scala 21:11]
  assign n80_I_2_1_t1b = n69_O_2_1_t1b; // @[Top.scala 21:11]
  assign n80_I_2_2_t0b = n69_O_2_2_t0b; // @[Top.scala 21:11]
  assign n80_I_2_2_t1b = n69_O_2_2_t1b; // @[Top.scala 21:11]
  assign n85_clock = clock;
  assign n85_reset = reset;
  assign n85_valid_up = n80_valid_down; // @[Top.scala 25:18]
  assign n85_I_0_0 = n80_O_0_0; // @[Top.scala 24:11]
  assign n85_I_0_1 = n80_O_0_1; // @[Top.scala 24:11]
  assign n85_I_0_2 = n80_O_0_2; // @[Top.scala 24:11]
  assign n85_I_1_0 = n80_O_1_0; // @[Top.scala 24:11]
  assign n85_I_1_1 = n80_O_1_1; // @[Top.scala 24:11]
  assign n85_I_1_2 = n80_O_1_2; // @[Top.scala 24:11]
  assign n85_I_2_0 = n80_O_2_0; // @[Top.scala 24:11]
  assign n85_I_2_1 = n80_O_2_1; // @[Top.scala 24:11]
  assign n85_I_2_2 = n80_O_2_2; // @[Top.scala 24:11]
  assign n90_clock = clock;
  assign n90_reset = reset;
  assign n90_valid_up = n85_valid_down; // @[Top.scala 28:18]
  assign n90_I_0_0 = n85_O_0_0; // @[Top.scala 27:11]
  assign n90_I_1_0 = n85_O_1_0; // @[Top.scala 27:11]
  assign n90_I_2_0 = n85_O_2_0; // @[Top.scala 27:11]
  assign InitialDelayCounter_1_clock = clock;
  assign InitialDelayCounter_1_reset = reset;
  assign n93_valid_up = n90_valid_down & InitialDelayCounter_1_valid_down; // @[Top.scala 33:18]
  assign n93_I0_0_0 = n90_O_0_0; // @[Top.scala 31:12]
  assign n104_valid_up = n93_valid_down; // @[Top.scala 36:19]
  assign n104_I_0_0_t0b = n93_O_0_0_t0b; // @[Top.scala 35:12]
  assign n104_I_0_0_t1b = n93_O_0_0_t1b; // @[Top.scala 35:12]
endmodule
module MapS_9(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  input  [7:0] I_1_1_0,
  input  [7:0] I_1_1_1,
  input  [7:0] I_1_1_2,
  input  [7:0] I_1_2_0,
  input  [7:0] I_1_2_1,
  input  [7:0] I_1_2_2,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_2_0_2,
  input  [7:0] I_2_1_0,
  input  [7:0] I_2_1_1,
  input  [7:0] I_2_1_2,
  input  [7:0] I_2_2_0,
  input  [7:0] I_2_2_1,
  input  [7:0] I_2_2_2,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_3_0_2,
  input  [7:0] I_3_1_0,
  input  [7:0] I_3_1_1,
  input  [7:0] I_3_1_2,
  input  [7:0] I_3_2_0,
  input  [7:0] I_3_2_1,
  input  [7:0] I_3_2_2,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_4_0_2,
  input  [7:0] I_4_1_0,
  input  [7:0] I_4_1_1,
  input  [7:0] I_4_1_2,
  input  [7:0] I_4_2_0,
  input  [7:0] I_4_2_1,
  input  [7:0] I_4_2_2,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_5_0_2,
  input  [7:0] I_5_1_0,
  input  [7:0] I_5_1_1,
  input  [7:0] I_5_1_2,
  input  [7:0] I_5_2_0,
  input  [7:0] I_5_2_1,
  input  [7:0] I_5_2_2,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_6_0_2,
  input  [7:0] I_6_1_0,
  input  [7:0] I_6_1_1,
  input  [7:0] I_6_1_2,
  input  [7:0] I_6_2_0,
  input  [7:0] I_6_2_1,
  input  [7:0] I_6_2_2,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_7_0_2,
  input  [7:0] I_7_1_0,
  input  [7:0] I_7_1_1,
  input  [7:0] I_7_1_2,
  input  [7:0] I_7_2_0,
  input  [7:0] I_7_2_1,
  input  [7:0] I_7_2_2,
  input  [7:0] I_8_0_0,
  input  [7:0] I_8_0_1,
  input  [7:0] I_8_0_2,
  input  [7:0] I_8_1_0,
  input  [7:0] I_8_1_1,
  input  [7:0] I_8_1_2,
  input  [7:0] I_8_2_0,
  input  [7:0] I_8_2_1,
  input  [7:0] I_8_2_2,
  input  [7:0] I_9_0_0,
  input  [7:0] I_9_0_1,
  input  [7:0] I_9_0_2,
  input  [7:0] I_9_1_0,
  input  [7:0] I_9_1_1,
  input  [7:0] I_9_1_2,
  input  [7:0] I_9_2_0,
  input  [7:0] I_9_2_1,
  input  [7:0] I_9_2_2,
  input  [7:0] I_10_0_0,
  input  [7:0] I_10_0_1,
  input  [7:0] I_10_0_2,
  input  [7:0] I_10_1_0,
  input  [7:0] I_10_1_1,
  input  [7:0] I_10_1_2,
  input  [7:0] I_10_2_0,
  input  [7:0] I_10_2_1,
  input  [7:0] I_10_2_2,
  input  [7:0] I_11_0_0,
  input  [7:0] I_11_0_1,
  input  [7:0] I_11_0_2,
  input  [7:0] I_11_1_0,
  input  [7:0] I_11_1_1,
  input  [7:0] I_11_1_2,
  input  [7:0] I_11_2_0,
  input  [7:0] I_11_2_1,
  input  [7:0] I_11_2_2,
  input  [7:0] I_12_0_0,
  input  [7:0] I_12_0_1,
  input  [7:0] I_12_0_2,
  input  [7:0] I_12_1_0,
  input  [7:0] I_12_1_1,
  input  [7:0] I_12_1_2,
  input  [7:0] I_12_2_0,
  input  [7:0] I_12_2_1,
  input  [7:0] I_12_2_2,
  input  [7:0] I_13_0_0,
  input  [7:0] I_13_0_1,
  input  [7:0] I_13_0_2,
  input  [7:0] I_13_1_0,
  input  [7:0] I_13_1_1,
  input  [7:0] I_13_1_2,
  input  [7:0] I_13_2_0,
  input  [7:0] I_13_2_1,
  input  [7:0] I_13_2_2,
  input  [7:0] I_14_0_0,
  input  [7:0] I_14_0_1,
  input  [7:0] I_14_0_2,
  input  [7:0] I_14_1_0,
  input  [7:0] I_14_1_1,
  input  [7:0] I_14_1_2,
  input  [7:0] I_14_2_0,
  input  [7:0] I_14_2_1,
  input  [7:0] I_14_2_2,
  input  [7:0] I_15_0_0,
  input  [7:0] I_15_0_1,
  input  [7:0] I_15_0_2,
  input  [7:0] I_15_1_0,
  input  [7:0] I_15_1_1,
  input  [7:0] I_15_1_2,
  input  [7:0] I_15_2_0,
  input  [7:0] I_15_2_1,
  input  [7:0] I_15_2_2,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0,
  output [7:0] O_8_0_0,
  output [7:0] O_9_0_0,
  output [7:0] O_10_0_0,
  output [7:0] O_11_0_0,
  output [7:0] O_12_0_0,
  output [7:0] O_13_0_0,
  output [7:0] O_14_0_0,
  output [7:0] O_15_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_2_clock; // @[MapS.scala 10:86]
  wire  other_ops_2_reset; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_3_clock; // @[MapS.scala 10:86]
  wire  other_ops_3_reset; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_4_clock; // @[MapS.scala 10:86]
  wire  other_ops_4_reset; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_5_clock; // @[MapS.scala 10:86]
  wire  other_ops_5_reset; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_6_clock; // @[MapS.scala 10:86]
  wire  other_ops_6_reset; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_7_clock; // @[MapS.scala 10:86]
  wire  other_ops_7_reset; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_8_clock; // @[MapS.scala 10:86]
  wire  other_ops_8_reset; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_9_clock; // @[MapS.scala 10:86]
  wire  other_ops_9_reset; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_10_clock; // @[MapS.scala 10:86]
  wire  other_ops_10_reset; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_11_clock; // @[MapS.scala 10:86]
  wire  other_ops_11_reset; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_12_clock; // @[MapS.scala 10:86]
  wire  other_ops_12_reset; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_13_clock; // @[MapS.scala 10:86]
  wire  other_ops_13_reset; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_14_clock; // @[MapS.scala 10:86]
  wire  other_ops_14_reset; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  Module_0 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .I_1_0(fst_op_I_1_0),
    .I_1_1(fst_op_I_1_1),
    .I_1_2(fst_op_I_1_2),
    .I_2_0(fst_op_I_2_0),
    .I_2_1(fst_op_I_2_1),
    .I_2_2(fst_op_I_2_2),
    .O_0_0(fst_op_O_0_0)
  );
  Module_0 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .I_1_0(other_ops_0_I_1_0),
    .I_1_1(other_ops_0_I_1_1),
    .I_1_2(other_ops_0_I_1_2),
    .I_2_0(other_ops_0_I_2_0),
    .I_2_1(other_ops_0_I_2_1),
    .I_2_2(other_ops_0_I_2_2),
    .O_0_0(other_ops_0_O_0_0)
  );
  Module_0 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_0_2(other_ops_1_I_0_2),
    .I_1_0(other_ops_1_I_1_0),
    .I_1_1(other_ops_1_I_1_1),
    .I_1_2(other_ops_1_I_1_2),
    .I_2_0(other_ops_1_I_2_0),
    .I_2_1(other_ops_1_I_2_1),
    .I_2_2(other_ops_1_I_2_2),
    .O_0_0(other_ops_1_O_0_0)
  );
  Module_0 other_ops_2 ( // @[MapS.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_0_2(other_ops_2_I_0_2),
    .I_1_0(other_ops_2_I_1_0),
    .I_1_1(other_ops_2_I_1_1),
    .I_1_2(other_ops_2_I_1_2),
    .I_2_0(other_ops_2_I_2_0),
    .I_2_1(other_ops_2_I_2_1),
    .I_2_2(other_ops_2_I_2_2),
    .O_0_0(other_ops_2_O_0_0)
  );
  Module_0 other_ops_3 ( // @[MapS.scala 10:86]
    .clock(other_ops_3_clock),
    .reset(other_ops_3_reset),
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0(other_ops_3_I_0_0),
    .I_0_1(other_ops_3_I_0_1),
    .I_0_2(other_ops_3_I_0_2),
    .I_1_0(other_ops_3_I_1_0),
    .I_1_1(other_ops_3_I_1_1),
    .I_1_2(other_ops_3_I_1_2),
    .I_2_0(other_ops_3_I_2_0),
    .I_2_1(other_ops_3_I_2_1),
    .I_2_2(other_ops_3_I_2_2),
    .O_0_0(other_ops_3_O_0_0)
  );
  Module_0 other_ops_4 ( // @[MapS.scala 10:86]
    .clock(other_ops_4_clock),
    .reset(other_ops_4_reset),
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0(other_ops_4_I_0_0),
    .I_0_1(other_ops_4_I_0_1),
    .I_0_2(other_ops_4_I_0_2),
    .I_1_0(other_ops_4_I_1_0),
    .I_1_1(other_ops_4_I_1_1),
    .I_1_2(other_ops_4_I_1_2),
    .I_2_0(other_ops_4_I_2_0),
    .I_2_1(other_ops_4_I_2_1),
    .I_2_2(other_ops_4_I_2_2),
    .O_0_0(other_ops_4_O_0_0)
  );
  Module_0 other_ops_5 ( // @[MapS.scala 10:86]
    .clock(other_ops_5_clock),
    .reset(other_ops_5_reset),
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0(other_ops_5_I_0_0),
    .I_0_1(other_ops_5_I_0_1),
    .I_0_2(other_ops_5_I_0_2),
    .I_1_0(other_ops_5_I_1_0),
    .I_1_1(other_ops_5_I_1_1),
    .I_1_2(other_ops_5_I_1_2),
    .I_2_0(other_ops_5_I_2_0),
    .I_2_1(other_ops_5_I_2_1),
    .I_2_2(other_ops_5_I_2_2),
    .O_0_0(other_ops_5_O_0_0)
  );
  Module_0 other_ops_6 ( // @[MapS.scala 10:86]
    .clock(other_ops_6_clock),
    .reset(other_ops_6_reset),
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0(other_ops_6_I_0_0),
    .I_0_1(other_ops_6_I_0_1),
    .I_0_2(other_ops_6_I_0_2),
    .I_1_0(other_ops_6_I_1_0),
    .I_1_1(other_ops_6_I_1_1),
    .I_1_2(other_ops_6_I_1_2),
    .I_2_0(other_ops_6_I_2_0),
    .I_2_1(other_ops_6_I_2_1),
    .I_2_2(other_ops_6_I_2_2),
    .O_0_0(other_ops_6_O_0_0)
  );
  Module_0 other_ops_7 ( // @[MapS.scala 10:86]
    .clock(other_ops_7_clock),
    .reset(other_ops_7_reset),
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I_0_0(other_ops_7_I_0_0),
    .I_0_1(other_ops_7_I_0_1),
    .I_0_2(other_ops_7_I_0_2),
    .I_1_0(other_ops_7_I_1_0),
    .I_1_1(other_ops_7_I_1_1),
    .I_1_2(other_ops_7_I_1_2),
    .I_2_0(other_ops_7_I_2_0),
    .I_2_1(other_ops_7_I_2_1),
    .I_2_2(other_ops_7_I_2_2),
    .O_0_0(other_ops_7_O_0_0)
  );
  Module_0 other_ops_8 ( // @[MapS.scala 10:86]
    .clock(other_ops_8_clock),
    .reset(other_ops_8_reset),
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I_0_0(other_ops_8_I_0_0),
    .I_0_1(other_ops_8_I_0_1),
    .I_0_2(other_ops_8_I_0_2),
    .I_1_0(other_ops_8_I_1_0),
    .I_1_1(other_ops_8_I_1_1),
    .I_1_2(other_ops_8_I_1_2),
    .I_2_0(other_ops_8_I_2_0),
    .I_2_1(other_ops_8_I_2_1),
    .I_2_2(other_ops_8_I_2_2),
    .O_0_0(other_ops_8_O_0_0)
  );
  Module_0 other_ops_9 ( // @[MapS.scala 10:86]
    .clock(other_ops_9_clock),
    .reset(other_ops_9_reset),
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I_0_0(other_ops_9_I_0_0),
    .I_0_1(other_ops_9_I_0_1),
    .I_0_2(other_ops_9_I_0_2),
    .I_1_0(other_ops_9_I_1_0),
    .I_1_1(other_ops_9_I_1_1),
    .I_1_2(other_ops_9_I_1_2),
    .I_2_0(other_ops_9_I_2_0),
    .I_2_1(other_ops_9_I_2_1),
    .I_2_2(other_ops_9_I_2_2),
    .O_0_0(other_ops_9_O_0_0)
  );
  Module_0 other_ops_10 ( // @[MapS.scala 10:86]
    .clock(other_ops_10_clock),
    .reset(other_ops_10_reset),
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I_0_0(other_ops_10_I_0_0),
    .I_0_1(other_ops_10_I_0_1),
    .I_0_2(other_ops_10_I_0_2),
    .I_1_0(other_ops_10_I_1_0),
    .I_1_1(other_ops_10_I_1_1),
    .I_1_2(other_ops_10_I_1_2),
    .I_2_0(other_ops_10_I_2_0),
    .I_2_1(other_ops_10_I_2_1),
    .I_2_2(other_ops_10_I_2_2),
    .O_0_0(other_ops_10_O_0_0)
  );
  Module_0 other_ops_11 ( // @[MapS.scala 10:86]
    .clock(other_ops_11_clock),
    .reset(other_ops_11_reset),
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I_0_0(other_ops_11_I_0_0),
    .I_0_1(other_ops_11_I_0_1),
    .I_0_2(other_ops_11_I_0_2),
    .I_1_0(other_ops_11_I_1_0),
    .I_1_1(other_ops_11_I_1_1),
    .I_1_2(other_ops_11_I_1_2),
    .I_2_0(other_ops_11_I_2_0),
    .I_2_1(other_ops_11_I_2_1),
    .I_2_2(other_ops_11_I_2_2),
    .O_0_0(other_ops_11_O_0_0)
  );
  Module_0 other_ops_12 ( // @[MapS.scala 10:86]
    .clock(other_ops_12_clock),
    .reset(other_ops_12_reset),
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I_0_0(other_ops_12_I_0_0),
    .I_0_1(other_ops_12_I_0_1),
    .I_0_2(other_ops_12_I_0_2),
    .I_1_0(other_ops_12_I_1_0),
    .I_1_1(other_ops_12_I_1_1),
    .I_1_2(other_ops_12_I_1_2),
    .I_2_0(other_ops_12_I_2_0),
    .I_2_1(other_ops_12_I_2_1),
    .I_2_2(other_ops_12_I_2_2),
    .O_0_0(other_ops_12_O_0_0)
  );
  Module_0 other_ops_13 ( // @[MapS.scala 10:86]
    .clock(other_ops_13_clock),
    .reset(other_ops_13_reset),
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I_0_0(other_ops_13_I_0_0),
    .I_0_1(other_ops_13_I_0_1),
    .I_0_2(other_ops_13_I_0_2),
    .I_1_0(other_ops_13_I_1_0),
    .I_1_1(other_ops_13_I_1_1),
    .I_1_2(other_ops_13_I_1_2),
    .I_2_0(other_ops_13_I_2_0),
    .I_2_1(other_ops_13_I_2_1),
    .I_2_2(other_ops_13_I_2_2),
    .O_0_0(other_ops_13_O_0_0)
  );
  Module_0 other_ops_14 ( // @[MapS.scala 10:86]
    .clock(other_ops_14_clock),
    .reset(other_ops_14_reset),
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I_0_0(other_ops_14_I_0_0),
    .I_0_1(other_ops_14_I_0_1),
    .I_0_2(other_ops_14_I_0_2),
    .I_1_0(other_ops_14_I_1_0),
    .I_1_1(other_ops_14_I_1_1),
    .I_1_2(other_ops_14_I_1_2),
    .I_2_0(other_ops_14_I_2_0),
    .I_2_1(other_ops_14_I_2_1),
    .I_2_2(other_ops_14_I_2_2),
    .O_0_0(other_ops_14_O_0_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[MapS.scala 21:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[MapS.scala 21:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[MapS.scala 21:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[MapS.scala 21:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[MapS.scala 21:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[MapS.scala 21:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[MapS.scala 21:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_1_0 = I_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_1_1 = I_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_1_2 = I_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_2_0 = I_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_2_1 = I_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_2_2 = I_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_0 = I_1_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_1 = I_1_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_2 = I_1_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_0 = I_1_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_1 = I_1_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_2 = I_1_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2 = I_2_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_0 = I_2_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_1 = I_2_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_2 = I_2_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_0 = I_2_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_1 = I_2_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_2 = I_2_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_2_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2 = I_3_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_0 = I_3_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_1 = I_3_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_2 = I_3_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_0 = I_3_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_1 = I_3_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_2 = I_3_2_2; // @[MapS.scala 20:41]
  assign other_ops_3_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_3_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0 = I_4_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1 = I_4_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2 = I_4_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_0 = I_4_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_1 = I_4_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_2 = I_4_1_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_0 = I_4_2_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_1 = I_4_2_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_2 = I_4_2_2; // @[MapS.scala 20:41]
  assign other_ops_4_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_4_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0 = I_5_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1 = I_5_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2 = I_5_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_0 = I_5_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_1 = I_5_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_2 = I_5_1_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_0 = I_5_2_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_1 = I_5_2_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_2 = I_5_2_2; // @[MapS.scala 20:41]
  assign other_ops_5_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_5_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0 = I_6_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1 = I_6_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2 = I_6_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_0 = I_6_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_1 = I_6_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_2 = I_6_1_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_0 = I_6_2_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_1 = I_6_2_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_2 = I_6_2_2; // @[MapS.scala 20:41]
  assign other_ops_6_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_6_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0 = I_7_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1 = I_7_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2 = I_7_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_0 = I_7_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_1 = I_7_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_2 = I_7_1_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_0 = I_7_2_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_1 = I_7_2_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_2 = I_7_2_2; // @[MapS.scala 20:41]
  assign other_ops_7_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_7_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I_0_0 = I_8_0_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1 = I_8_0_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2 = I_8_0_2; // @[MapS.scala 20:41]
  assign other_ops_7_I_1_0 = I_8_1_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_1_1 = I_8_1_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_1_2 = I_8_1_2; // @[MapS.scala 20:41]
  assign other_ops_7_I_2_0 = I_8_2_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_2_1 = I_8_2_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_2_2 = I_8_2_2; // @[MapS.scala 20:41]
  assign other_ops_8_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_8_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I_0_0 = I_9_0_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1 = I_9_0_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2 = I_9_0_2; // @[MapS.scala 20:41]
  assign other_ops_8_I_1_0 = I_9_1_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_1_1 = I_9_1_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_1_2 = I_9_1_2; // @[MapS.scala 20:41]
  assign other_ops_8_I_2_0 = I_9_2_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_2_1 = I_9_2_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_2_2 = I_9_2_2; // @[MapS.scala 20:41]
  assign other_ops_9_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_9_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I_0_0 = I_10_0_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1 = I_10_0_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2 = I_10_0_2; // @[MapS.scala 20:41]
  assign other_ops_9_I_1_0 = I_10_1_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_1_1 = I_10_1_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_1_2 = I_10_1_2; // @[MapS.scala 20:41]
  assign other_ops_9_I_2_0 = I_10_2_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_2_1 = I_10_2_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_2_2 = I_10_2_2; // @[MapS.scala 20:41]
  assign other_ops_10_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_10_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I_0_0 = I_11_0_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1 = I_11_0_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2 = I_11_0_2; // @[MapS.scala 20:41]
  assign other_ops_10_I_1_0 = I_11_1_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_1_1 = I_11_1_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_1_2 = I_11_1_2; // @[MapS.scala 20:41]
  assign other_ops_10_I_2_0 = I_11_2_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_2_1 = I_11_2_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_2_2 = I_11_2_2; // @[MapS.scala 20:41]
  assign other_ops_11_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_11_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I_0_0 = I_12_0_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1 = I_12_0_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2 = I_12_0_2; // @[MapS.scala 20:41]
  assign other_ops_11_I_1_0 = I_12_1_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_1_1 = I_12_1_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_1_2 = I_12_1_2; // @[MapS.scala 20:41]
  assign other_ops_11_I_2_0 = I_12_2_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_2_1 = I_12_2_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_2_2 = I_12_2_2; // @[MapS.scala 20:41]
  assign other_ops_12_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_12_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I_0_0 = I_13_0_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1 = I_13_0_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2 = I_13_0_2; // @[MapS.scala 20:41]
  assign other_ops_12_I_1_0 = I_13_1_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_1_1 = I_13_1_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_1_2 = I_13_1_2; // @[MapS.scala 20:41]
  assign other_ops_12_I_2_0 = I_13_2_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_2_1 = I_13_2_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_2_2 = I_13_2_2; // @[MapS.scala 20:41]
  assign other_ops_13_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_13_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I_0_0 = I_14_0_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1 = I_14_0_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2 = I_14_0_2; // @[MapS.scala 20:41]
  assign other_ops_13_I_1_0 = I_14_1_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_1_1 = I_14_1_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_1_2 = I_14_1_2; // @[MapS.scala 20:41]
  assign other_ops_13_I_2_0 = I_14_2_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_2_1 = I_14_2_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_2_2 = I_14_2_2; // @[MapS.scala 20:41]
  assign other_ops_14_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_14_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I_0_0 = I_15_0_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1 = I_15_0_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2 = I_15_0_2; // @[MapS.scala 20:41]
  assign other_ops_14_I_1_0 = I_15_1_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_1_1 = I_15_1_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_1_2 = I_15_1_2; // @[MapS.scala 20:41]
  assign other_ops_14_I_2_0 = I_15_2_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_2_1 = I_15_2_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_2_2 = I_15_2_2; // @[MapS.scala 20:41]
endmodule
module UnpartitionS(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_1_0_0,
  input  [7:0] I_2_0_0,
  input  [7:0] I_3_0_0,
  input  [7:0] I_4_0_0,
  input  [7:0] I_5_0_0,
  input  [7:0] I_6_0_0,
  input  [7:0] I_7_0_0,
  input  [7:0] I_8_0_0,
  input  [7:0] I_9_0_0,
  input  [7:0] I_10_0_0,
  input  [7:0] I_11_0_0,
  input  [7:0] I_12_0_0,
  input  [7:0] I_13_0_0,
  input  [7:0] I_14_0_0,
  input  [7:0] I_15_0_0,
  output [7:0] O_0_0,
  output [7:0] O_1_0,
  output [7:0] O_2_0,
  output [7:0] O_3_0,
  output [7:0] O_4_0,
  output [7:0] O_5_0,
  output [7:0] O_6_0,
  output [7:0] O_7_0,
  output [7:0] O_8_0,
  output [7:0] O_9_0,
  output [7:0] O_10_0,
  output [7:0] O_11_0,
  output [7:0] O_12_0,
  output [7:0] O_13_0,
  output [7:0] O_14_0,
  output [7:0] O_15_0
);
  assign valid_down = valid_up; // @[Partition.scala 31:14]
  assign O_0_0 = I_0_0_0; // @[Partition.scala 28:19]
  assign O_1_0 = I_1_0_0; // @[Partition.scala 28:19]
  assign O_2_0 = I_2_0_0; // @[Partition.scala 28:19]
  assign O_3_0 = I_3_0_0; // @[Partition.scala 28:19]
  assign O_4_0 = I_4_0_0; // @[Partition.scala 28:19]
  assign O_5_0 = I_5_0_0; // @[Partition.scala 28:19]
  assign O_6_0 = I_6_0_0; // @[Partition.scala 28:19]
  assign O_7_0 = I_7_0_0; // @[Partition.scala 28:19]
  assign O_8_0 = I_8_0_0; // @[Partition.scala 28:19]
  assign O_9_0 = I_9_0_0; // @[Partition.scala 28:19]
  assign O_10_0 = I_10_0_0; // @[Partition.scala 28:19]
  assign O_11_0 = I_11_0_0; // @[Partition.scala 28:19]
  assign O_12_0 = I_12_0_0; // @[Partition.scala 28:19]
  assign O_13_0 = I_13_0_0; // @[Partition.scala 28:19]
  assign O_14_0 = I_14_0_0; // @[Partition.scala 28:19]
  assign O_15_0 = I_15_0_0; // @[Partition.scala 28:19]
endmodule
module UnpartitionS_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_1_0,
  input  [7:0] I_2_0,
  input  [7:0] I_3_0,
  input  [7:0] I_4_0,
  input  [7:0] I_5_0,
  input  [7:0] I_6_0,
  input  [7:0] I_7_0,
  input  [7:0] I_8_0,
  input  [7:0] I_9_0,
  input  [7:0] I_10_0,
  input  [7:0] I_11_0,
  input  [7:0] I_12_0,
  input  [7:0] I_13_0,
  input  [7:0] I_14_0,
  input  [7:0] I_15_0,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15
);
  assign valid_down = valid_up; // @[Partition.scala 31:14]
  assign O_0 = I_0_0; // @[Partition.scala 28:19]
  assign O_1 = I_1_0; // @[Partition.scala 28:19]
  assign O_2 = I_2_0; // @[Partition.scala 28:19]
  assign O_3 = I_3_0; // @[Partition.scala 28:19]
  assign O_4 = I_4_0; // @[Partition.scala 28:19]
  assign O_5 = I_5_0; // @[Partition.scala 28:19]
  assign O_6 = I_6_0; // @[Partition.scala 28:19]
  assign O_7 = I_7_0; // @[Partition.scala 28:19]
  assign O_8 = I_8_0; // @[Partition.scala 28:19]
  assign O_9 = I_9_0; // @[Partition.scala 28:19]
  assign O_10 = I_10_0; // @[Partition.scala 28:19]
  assign O_11 = I_11_0; // @[Partition.scala 28:19]
  assign O_12 = I_12_0; // @[Partition.scala 28:19]
  assign O_13 = I_13_0; // @[Partition.scala 28:19]
  assign O_14 = I_14_0; // @[Partition.scala 28:19]
  assign O_15 = I_15_0; // @[Partition.scala 28:19]
endmodule
module FIFO_1(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  input  [7:0] I_4,
  input  [7:0] I_5,
  input  [7:0] I_6,
  input  [7:0] I_7,
  input  [7:0] I_8,
  input  [7:0] I_9,
  input  [7:0] I_10,
  input  [7:0] I_11,
  input  [7:0] I_12,
  input  [7:0] I_13,
  input  [7:0] I_14,
  input  [7:0] I_15,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15
);
  reg [7:0] _T__0 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_0;
  wire [7:0] _T__0__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__0__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_1;
  wire [7:0] _T__0__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__0__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__0__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__0__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__0__T_17_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [1:0] _T__0__T_17_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg [7:0] _T__1 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_4;
  wire [7:0] _T__1__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__1__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_5;
  wire [7:0] _T__1__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__1__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__1__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__1__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__1__T_17_en_pipe_0;
  reg [31:0] _RAND_6;
  reg [1:0] _T__1__T_17_addr_pipe_0;
  reg [31:0] _RAND_7;
  reg [7:0] _T__2 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_8;
  wire [7:0] _T__2__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__2__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_9;
  wire [7:0] _T__2__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__2__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__2__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__2__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__2__T_17_en_pipe_0;
  reg [31:0] _RAND_10;
  reg [1:0] _T__2__T_17_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [7:0] _T__3 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_12;
  wire [7:0] _T__3__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__3__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_13;
  wire [7:0] _T__3__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__3__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__3__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__3__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__3__T_17_en_pipe_0;
  reg [31:0] _RAND_14;
  reg [1:0] _T__3__T_17_addr_pipe_0;
  reg [31:0] _RAND_15;
  reg [7:0] _T__4 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_16;
  wire [7:0] _T__4__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__4__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_17;
  wire [7:0] _T__4__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__4__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__4__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__4__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__4__T_17_en_pipe_0;
  reg [31:0] _RAND_18;
  reg [1:0] _T__4__T_17_addr_pipe_0;
  reg [31:0] _RAND_19;
  reg [7:0] _T__5 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_20;
  wire [7:0] _T__5__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__5__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_21;
  wire [7:0] _T__5__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__5__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__5__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__5__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__5__T_17_en_pipe_0;
  reg [31:0] _RAND_22;
  reg [1:0] _T__5__T_17_addr_pipe_0;
  reg [31:0] _RAND_23;
  reg [7:0] _T__6 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_24;
  wire [7:0] _T__6__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__6__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_25;
  wire [7:0] _T__6__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__6__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__6__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__6__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__6__T_17_en_pipe_0;
  reg [31:0] _RAND_26;
  reg [1:0] _T__6__T_17_addr_pipe_0;
  reg [31:0] _RAND_27;
  reg [7:0] _T__7 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_28;
  wire [7:0] _T__7__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__7__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_29;
  wire [7:0] _T__7__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__7__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__7__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__7__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__7__T_17_en_pipe_0;
  reg [31:0] _RAND_30;
  reg [1:0] _T__7__T_17_addr_pipe_0;
  reg [31:0] _RAND_31;
  reg [7:0] _T__8 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_32;
  wire [7:0] _T__8__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__8__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_33;
  wire [7:0] _T__8__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__8__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__8__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__8__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__8__T_17_en_pipe_0;
  reg [31:0] _RAND_34;
  reg [1:0] _T__8__T_17_addr_pipe_0;
  reg [31:0] _RAND_35;
  reg [7:0] _T__9 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_36;
  wire [7:0] _T__9__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__9__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_37;
  wire [7:0] _T__9__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__9__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__9__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__9__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__9__T_17_en_pipe_0;
  reg [31:0] _RAND_38;
  reg [1:0] _T__9__T_17_addr_pipe_0;
  reg [31:0] _RAND_39;
  reg [7:0] _T__10 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_40;
  wire [7:0] _T__10__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__10__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_41;
  wire [7:0] _T__10__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__10__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__10__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__10__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__10__T_17_en_pipe_0;
  reg [31:0] _RAND_42;
  reg [1:0] _T__10__T_17_addr_pipe_0;
  reg [31:0] _RAND_43;
  reg [7:0] _T__11 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_44;
  wire [7:0] _T__11__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__11__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_45;
  wire [7:0] _T__11__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__11__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__11__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__11__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__11__T_17_en_pipe_0;
  reg [31:0] _RAND_46;
  reg [1:0] _T__11__T_17_addr_pipe_0;
  reg [31:0] _RAND_47;
  reg [7:0] _T__12 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_48;
  wire [7:0] _T__12__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__12__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_49;
  wire [7:0] _T__12__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__12__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__12__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__12__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__12__T_17_en_pipe_0;
  reg [31:0] _RAND_50;
  reg [1:0] _T__12__T_17_addr_pipe_0;
  reg [31:0] _RAND_51;
  reg [7:0] _T__13 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_52;
  wire [7:0] _T__13__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__13__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_53;
  wire [7:0] _T__13__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__13__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__13__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__13__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__13__T_17_en_pipe_0;
  reg [31:0] _RAND_54;
  reg [1:0] _T__13__T_17_addr_pipe_0;
  reg [31:0] _RAND_55;
  reg [7:0] _T__14 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_56;
  wire [7:0] _T__14__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__14__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_57;
  wire [7:0] _T__14__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__14__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__14__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__14__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__14__T_17_en_pipe_0;
  reg [31:0] _RAND_58;
  reg [1:0] _T__14__T_17_addr_pipe_0;
  reg [31:0] _RAND_59;
  reg [7:0] _T__15 [0:2]; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_60;
  wire [7:0] _T__15__T_17_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__15__T_17_addr; // @[FIFO.scala 23:33]
  reg [31:0] _RAND_61;
  wire [7:0] _T__15__T_5_data; // @[FIFO.scala 23:33]
  wire [1:0] _T__15__T_5_addr; // @[FIFO.scala 23:33]
  wire  _T__15__T_5_mask; // @[FIFO.scala 23:33]
  wire  _T__15__T_5_en; // @[FIFO.scala 23:33]
  reg  _T__15__T_17_en_pipe_0;
  reg [31:0] _RAND_62;
  reg [1:0] _T__15__T_17_addr_pipe_0;
  reg [31:0] _RAND_63;
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_64;
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg [31:0] _RAND_65;
  reg [1:0] value_2; // @[Counter.scala 29:33]
  reg [31:0] _RAND_66;
  wire  _T_1; // @[FIFO.scala 33:46]
  wire  _T_2; // @[Counter.scala 37:24]
  wire [1:0] _T_4; // @[Counter.scala 38:22]
  wire  _T_6; // @[FIFO.scala 38:39]
  wire [1:0] _T_11; // @[Counter.scala 38:22]
  wire  _T_12; // @[FIFO.scala 42:39]
  wire  _T_18; // @[Counter.scala 37:24]
  wire [1:0] _T_20; // @[Counter.scala 38:22]
  wire  _GEN_8; // @[FIFO.scala 42:57]
  wire  _GEN_70; // @[FIFO.scala 39:15]
  assign _T__0__T_17_addr = _T__0__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__0__T_17_data = _T__0[_T__0__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__0__T_17_data = _T__0__T_17_addr >= 2'h3 ? _RAND_1[7:0] : _T__0[_T__0__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__0__T_5_data = I_0;
  assign _T__0__T_5_addr = value_2;
  assign _T__0__T_5_mask = 1'h1;
  assign _T__0__T_5_en = valid_up;
  assign _T__1__T_17_addr = _T__1__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__1__T_17_data = _T__1[_T__1__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__1__T_17_data = _T__1__T_17_addr >= 2'h3 ? _RAND_5[7:0] : _T__1[_T__1__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__1__T_5_data = I_1;
  assign _T__1__T_5_addr = value_2;
  assign _T__1__T_5_mask = 1'h1;
  assign _T__1__T_5_en = valid_up;
  assign _T__2__T_17_addr = _T__2__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__2__T_17_data = _T__2[_T__2__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__2__T_17_data = _T__2__T_17_addr >= 2'h3 ? _RAND_9[7:0] : _T__2[_T__2__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__2__T_5_data = I_2;
  assign _T__2__T_5_addr = value_2;
  assign _T__2__T_5_mask = 1'h1;
  assign _T__2__T_5_en = valid_up;
  assign _T__3__T_17_addr = _T__3__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__3__T_17_data = _T__3[_T__3__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__3__T_17_data = _T__3__T_17_addr >= 2'h3 ? _RAND_13[7:0] : _T__3[_T__3__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__3__T_5_data = I_3;
  assign _T__3__T_5_addr = value_2;
  assign _T__3__T_5_mask = 1'h1;
  assign _T__3__T_5_en = valid_up;
  assign _T__4__T_17_addr = _T__4__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__4__T_17_data = _T__4[_T__4__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__4__T_17_data = _T__4__T_17_addr >= 2'h3 ? _RAND_17[7:0] : _T__4[_T__4__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__4__T_5_data = I_4;
  assign _T__4__T_5_addr = value_2;
  assign _T__4__T_5_mask = 1'h1;
  assign _T__4__T_5_en = valid_up;
  assign _T__5__T_17_addr = _T__5__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__5__T_17_data = _T__5[_T__5__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__5__T_17_data = _T__5__T_17_addr >= 2'h3 ? _RAND_21[7:0] : _T__5[_T__5__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__5__T_5_data = I_5;
  assign _T__5__T_5_addr = value_2;
  assign _T__5__T_5_mask = 1'h1;
  assign _T__5__T_5_en = valid_up;
  assign _T__6__T_17_addr = _T__6__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__6__T_17_data = _T__6[_T__6__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__6__T_17_data = _T__6__T_17_addr >= 2'h3 ? _RAND_25[7:0] : _T__6[_T__6__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__6__T_5_data = I_6;
  assign _T__6__T_5_addr = value_2;
  assign _T__6__T_5_mask = 1'h1;
  assign _T__6__T_5_en = valid_up;
  assign _T__7__T_17_addr = _T__7__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__7__T_17_data = _T__7[_T__7__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__7__T_17_data = _T__7__T_17_addr >= 2'h3 ? _RAND_29[7:0] : _T__7[_T__7__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__7__T_5_data = I_7;
  assign _T__7__T_5_addr = value_2;
  assign _T__7__T_5_mask = 1'h1;
  assign _T__7__T_5_en = valid_up;
  assign _T__8__T_17_addr = _T__8__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__8__T_17_data = _T__8[_T__8__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__8__T_17_data = _T__8__T_17_addr >= 2'h3 ? _RAND_33[7:0] : _T__8[_T__8__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__8__T_5_data = I_8;
  assign _T__8__T_5_addr = value_2;
  assign _T__8__T_5_mask = 1'h1;
  assign _T__8__T_5_en = valid_up;
  assign _T__9__T_17_addr = _T__9__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__9__T_17_data = _T__9[_T__9__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__9__T_17_data = _T__9__T_17_addr >= 2'h3 ? _RAND_37[7:0] : _T__9[_T__9__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__9__T_5_data = I_9;
  assign _T__9__T_5_addr = value_2;
  assign _T__9__T_5_mask = 1'h1;
  assign _T__9__T_5_en = valid_up;
  assign _T__10__T_17_addr = _T__10__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__10__T_17_data = _T__10[_T__10__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__10__T_17_data = _T__10__T_17_addr >= 2'h3 ? _RAND_41[7:0] : _T__10[_T__10__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__10__T_5_data = I_10;
  assign _T__10__T_5_addr = value_2;
  assign _T__10__T_5_mask = 1'h1;
  assign _T__10__T_5_en = valid_up;
  assign _T__11__T_17_addr = _T__11__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__11__T_17_data = _T__11[_T__11__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__11__T_17_data = _T__11__T_17_addr >= 2'h3 ? _RAND_45[7:0] : _T__11[_T__11__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__11__T_5_data = I_11;
  assign _T__11__T_5_addr = value_2;
  assign _T__11__T_5_mask = 1'h1;
  assign _T__11__T_5_en = valid_up;
  assign _T__12__T_17_addr = _T__12__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__12__T_17_data = _T__12[_T__12__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__12__T_17_data = _T__12__T_17_addr >= 2'h3 ? _RAND_49[7:0] : _T__12[_T__12__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__12__T_5_data = I_12;
  assign _T__12__T_5_addr = value_2;
  assign _T__12__T_5_mask = 1'h1;
  assign _T__12__T_5_en = valid_up;
  assign _T__13__T_17_addr = _T__13__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__13__T_17_data = _T__13[_T__13__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__13__T_17_data = _T__13__T_17_addr >= 2'h3 ? _RAND_53[7:0] : _T__13[_T__13__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__13__T_5_data = I_13;
  assign _T__13__T_5_addr = value_2;
  assign _T__13__T_5_mask = 1'h1;
  assign _T__13__T_5_en = valid_up;
  assign _T__14__T_17_addr = _T__14__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__14__T_17_data = _T__14[_T__14__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__14__T_17_data = _T__14__T_17_addr >= 2'h3 ? _RAND_57[7:0] : _T__14[_T__14__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__14__T_5_data = I_14;
  assign _T__14__T_5_addr = value_2;
  assign _T__14__T_5_mask = 1'h1;
  assign _T__14__T_5_en = valid_up;
  assign _T__15__T_17_addr = _T__15__T_17_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__15__T_17_data = _T__15[_T__15__T_17_addr]; // @[FIFO.scala 23:33]
  `else
  assign _T__15__T_17_data = _T__15__T_17_addr >= 2'h3 ? _RAND_61[7:0] : _T__15[_T__15__T_17_addr]; // @[FIFO.scala 23:33]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__15__T_5_data = I_15;
  assign _T__15__T_5_addr = value_2;
  assign _T__15__T_5_mask = 1'h1;
  assign _T__15__T_5_en = valid_up;
  assign _T_1 = value == 2'h2; // @[FIFO.scala 33:46]
  assign _T_2 = value_2 == 2'h2; // @[Counter.scala 37:24]
  assign _T_4 = value_2 + 2'h1; // @[Counter.scala 38:22]
  assign _T_6 = value < 2'h2; // @[FIFO.scala 38:39]
  assign _T_11 = value + 2'h1; // @[Counter.scala 38:22]
  assign _T_12 = value >= 2'h1; // @[FIFO.scala 42:39]
  assign _T_18 = value_1 == 2'h2; // @[Counter.scala 37:24]
  assign _T_20 = value_1 + 2'h1; // @[Counter.scala 38:22]
  assign _GEN_8 = _T_12 & _T_12; // @[FIFO.scala 42:57]
  assign valid_down = value == 2'h2; // @[FIFO.scala 33:16]
  assign O_0 = _T__0__T_17_data; // @[FIFO.scala 43:11]
  assign O_1 = _T__1__T_17_data; // @[FIFO.scala 43:11]
  assign O_2 = _T__2__T_17_data; // @[FIFO.scala 43:11]
  assign O_3 = _T__3__T_17_data; // @[FIFO.scala 43:11]
  assign O_4 = _T__4__T_17_data; // @[FIFO.scala 43:11]
  assign O_5 = _T__5__T_17_data; // @[FIFO.scala 43:11]
  assign O_6 = _T__6__T_17_data; // @[FIFO.scala 43:11]
  assign O_7 = _T__7__T_17_data; // @[FIFO.scala 43:11]
  assign O_8 = _T__8__T_17_data; // @[FIFO.scala 43:11]
  assign O_9 = _T__9__T_17_data; // @[FIFO.scala 43:11]
  assign O_10 = _T__10__T_17_data; // @[FIFO.scala 43:11]
  assign O_11 = _T__11__T_17_data; // @[FIFO.scala 43:11]
  assign O_12 = _T__12__T_17_data; // @[FIFO.scala 43:11]
  assign O_13 = _T__13__T_17_data; // @[FIFO.scala 43:11]
  assign O_14 = _T__14__T_17_data; // @[FIFO.scala 43:11]
  assign O_15 = _T__15__T_17_data; // @[FIFO.scala 43:11]
  assign _GEN_70 = valid_up & _T_6; // @[FIFO.scala 39:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__0[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__0__T_17_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__0__T_17_addr_pipe_0 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__1[initvar] = _RAND_4[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__1__T_17_en_pipe_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__1__T_17_addr_pipe_0 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__2[initvar] = _RAND_8[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T__2__T_17_en_pipe_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T__2__T_17_addr_pipe_0 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__3[initvar] = _RAND_12[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_13 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T__3__T_17_en_pipe_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T__3__T_17_addr_pipe_0 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__4[initvar] = _RAND_16[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_17 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T__4__T_17_en_pipe_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T__4__T_17_addr_pipe_0 = _RAND_19[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__5[initvar] = _RAND_20[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_21 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T__5__T_17_en_pipe_0 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T__5__T_17_addr_pipe_0 = _RAND_23[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__6[initvar] = _RAND_24[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_25 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T__6__T_17_en_pipe_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T__6__T_17_addr_pipe_0 = _RAND_27[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__7[initvar] = _RAND_28[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_29 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T__7__T_17_en_pipe_0 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T__7__T_17_addr_pipe_0 = _RAND_31[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__8[initvar] = _RAND_32[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_33 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T__8__T_17_en_pipe_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T__8__T_17_addr_pipe_0 = _RAND_35[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__9[initvar] = _RAND_36[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_37 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T__9__T_17_en_pipe_0 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T__9__T_17_addr_pipe_0 = _RAND_39[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__10[initvar] = _RAND_40[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_41 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T__10__T_17_en_pipe_0 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T__10__T_17_addr_pipe_0 = _RAND_43[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__11[initvar] = _RAND_44[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_45 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T__11__T_17_en_pipe_0 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T__11__T_17_addr_pipe_0 = _RAND_47[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__12[initvar] = _RAND_48[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_49 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T__12__T_17_en_pipe_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T__12__T_17_addr_pipe_0 = _RAND_51[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__13[initvar] = _RAND_52[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_53 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T__13__T_17_en_pipe_0 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T__13__T_17_addr_pipe_0 = _RAND_55[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__14[initvar] = _RAND_56[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_57 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T__14__T_17_en_pipe_0 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T__14__T_17_addr_pipe_0 = _RAND_59[1:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    _T__15[initvar] = _RAND_60[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_61 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T__15__T_17_en_pipe_0 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T__15__T_17_addr_pipe_0 = _RAND_63[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  value = _RAND_64[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  value_1 = _RAND_65[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  value_2 = _RAND_66[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__0__T_5_en & _T__0__T_5_mask) begin
      _T__0[_T__0__T_5_addr] <= _T__0__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__0__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__0__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__1__T_5_en & _T__1__T_5_mask) begin
      _T__1[_T__1__T_5_addr] <= _T__1__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__1__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__1__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__2__T_5_en & _T__2__T_5_mask) begin
      _T__2[_T__2__T_5_addr] <= _T__2__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__2__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__2__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__3__T_5_en & _T__3__T_5_mask) begin
      _T__3[_T__3__T_5_addr] <= _T__3__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__3__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__3__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__4__T_5_en & _T__4__T_5_mask) begin
      _T__4[_T__4__T_5_addr] <= _T__4__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__4__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__4__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__5__T_5_en & _T__5__T_5_mask) begin
      _T__5[_T__5__T_5_addr] <= _T__5__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__5__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__5__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__6__T_5_en & _T__6__T_5_mask) begin
      _T__6[_T__6__T_5_addr] <= _T__6__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__6__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__6__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__7__T_5_en & _T__7__T_5_mask) begin
      _T__7[_T__7__T_5_addr] <= _T__7__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__7__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__7__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__8__T_5_en & _T__8__T_5_mask) begin
      _T__8[_T__8__T_5_addr] <= _T__8__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__8__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__8__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__9__T_5_en & _T__9__T_5_mask) begin
      _T__9[_T__9__T_5_addr] <= _T__9__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__9__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__9__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__10__T_5_en & _T__10__T_5_mask) begin
      _T__10[_T__10__T_5_addr] <= _T__10__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__10__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__10__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__11__T_5_en & _T__11__T_5_mask) begin
      _T__11[_T__11__T_5_addr] <= _T__11__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__11__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__11__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__12__T_5_en & _T__12__T_5_mask) begin
      _T__12[_T__12__T_5_addr] <= _T__12__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__12__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__12__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__13__T_5_en & _T__13__T_5_mask) begin
      _T__13[_T__13__T_5_addr] <= _T__13__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__13__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__13__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__14__T_5_en & _T__14__T_5_mask) begin
      _T__14[_T__14__T_5_addr] <= _T__14__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__14__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__14__T_17_addr_pipe_0 <= value_1;
    end
    if(_T__15__T_5_en & _T__15__T_5_mask) begin
      _T__15[_T__15__T_5_addr] <= _T__15__T_5_data; // @[FIFO.scala 23:33]
    end
    _T__15__T_17_en_pipe_0 <= valid_up & _GEN_8;
    if (valid_up & _GEN_8) begin
      _T__15__T_17_addr_pipe_0 <= value_1;
    end
    if (reset) begin
      value <= 2'h0;
    end else if (valid_up) begin
      if (_T_6) begin
        if (_T_1) begin
          value <= 2'h0;
        end else begin
          value <= _T_11;
        end
      end
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (valid_up) begin
      if (_T_12) begin
        if (_T_18) begin
          value_1 <= 2'h0;
        end else begin
          value_1 <= _T_20;
        end
      end
    end
    if (reset) begin
      value_2 <= 2'h0;
    end else if (valid_up) begin
      if (_T_2) begin
        value_2 <= 2'h0;
      end else begin
        value_2 <= _T_4;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_70 & ~reset) begin
          $fwrite(32'h80000002,"idc inc\n"); // @[FIFO.scala 39:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Sub(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 139:14]
  assign O = I_t0b - I_t1b; // @[Arithmetic.scala 137:7]
endmodule
module Lt(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  wire  _T; // @[Arithmetic.scala 332:25]
  assign _T = I_t0b < I_t1b; // @[Arithmetic.scala 332:25]
  assign valid_down = valid_up; // @[Arithmetic.scala 334:14]
  assign O = {{7'd0}, _T}; // @[Arithmetic.scala 332:7]
endmodule
module AtomTuple_6(
  input   valid_up,
  output  valid_down,
  input   I0,
  input   I1,
  output  O_t0b,
  output  O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b = I1; // @[Tuple.scala 50:9]
endmodule
module Or(
  input   valid_up,
  output  valid_down,
  input   I_t0b,
  input   I_t1b,
  output  O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 83:14]
  assign O = I_t0b | I_t1b; // @[Arithmetic.scala 82:5]
endmodule
module AtomTuple_8(
  input        valid_up,
  output       valid_down,
  input        I0,
  input  [7:0] I1_t0b,
  input  [7:0] I1_t1b,
  output       O_t0b,
  output [7:0] O_t1b_t0b,
  output [7:0] O_t1b_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b_t0b = I1_t0b; // @[Tuple.scala 50:9]
  assign O_t1b_t1b = I1_t1b; // @[Tuple.scala 50:9]
endmodule
module If(
  input        valid_up,
  output       valid_down,
  input        I_t0b,
  input  [7:0] I_t1b_t0b,
  input  [7:0] I_t1b_t1b,
  output [7:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 395:14]
  assign O = I_t0b ? I_t1b_t0b : I_t1b_t1b; // @[Arithmetic.scala 393:9 Arithmetic.scala 394:20]
endmodule
module Add(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 108:14]
  assign O = I_t0b + I_t1b; // @[Arithmetic.scala 106:7]
endmodule
module Module_1(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  input  [7:0] I1,
  output [7:0] O
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n113_valid_up; // @[Top.scala 46:22]
  wire  n113_valid_down; // @[Top.scala 46:22]
  wire [7:0] n113_I0; // @[Top.scala 46:22]
  wire [7:0] n113_I1; // @[Top.scala 46:22]
  wire [7:0] n113_O_t0b; // @[Top.scala 46:22]
  wire [7:0] n113_O_t1b; // @[Top.scala 46:22]
  wire  n114_valid_up; // @[Top.scala 50:22]
  wire  n114_valid_down; // @[Top.scala 50:22]
  wire [7:0] n114_I_t0b; // @[Top.scala 50:22]
  wire [7:0] n114_I_t1b; // @[Top.scala 50:22]
  wire [7:0] n114_O; // @[Top.scala 50:22]
  wire  n116_valid_up; // @[Top.scala 53:22]
  wire  n116_valid_down; // @[Top.scala 53:22]
  wire [7:0] n116_I0; // @[Top.scala 53:22]
  wire [7:0] n116_I1; // @[Top.scala 53:22]
  wire [7:0] n116_O_t0b; // @[Top.scala 53:22]
  wire [7:0] n116_O_t1b; // @[Top.scala 53:22]
  wire  n117_valid_up; // @[Top.scala 57:22]
  wire  n117_valid_down; // @[Top.scala 57:22]
  wire [7:0] n117_I_t0b; // @[Top.scala 57:22]
  wire [7:0] n117_I_t1b; // @[Top.scala 57:22]
  wire [7:0] n117_O; // @[Top.scala 57:22]
  wire  InitialDelayCounter_1_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_valid_down; // @[Const.scala 11:33]
  wire  n118_valid_up; // @[Top.scala 61:22]
  wire  n118_valid_down; // @[Top.scala 61:22]
  wire [7:0] n118_I0; // @[Top.scala 61:22]
  wire [7:0] n118_I1; // @[Top.scala 61:22]
  wire [7:0] n118_O_t0b; // @[Top.scala 61:22]
  wire [7:0] n118_O_t1b; // @[Top.scala 61:22]
  wire  n119_valid_up; // @[Top.scala 65:22]
  wire  n119_valid_down; // @[Top.scala 65:22]
  wire [7:0] n119_I_t0b; // @[Top.scala 65:22]
  wire [7:0] n119_I_t1b; // @[Top.scala 65:22]
  wire [7:0] n119_O; // @[Top.scala 65:22]
  wire  n121_valid_up; // @[Top.scala 68:22]
  wire  n121_valid_down; // @[Top.scala 68:22]
  wire [7:0] n121_I0; // @[Top.scala 68:22]
  wire [7:0] n121_I1; // @[Top.scala 68:22]
  wire [7:0] n121_O_t0b; // @[Top.scala 68:22]
  wire [7:0] n121_O_t1b; // @[Top.scala 68:22]
  wire  n122_valid_up; // @[Top.scala 72:22]
  wire  n122_valid_down; // @[Top.scala 72:22]
  wire [7:0] n122_I_t0b; // @[Top.scala 72:22]
  wire [7:0] n122_I_t1b; // @[Top.scala 72:22]
  wire [7:0] n122_O; // @[Top.scala 72:22]
  wire  n123_valid_up; // @[Top.scala 75:22]
  wire  n123_valid_down; // @[Top.scala 75:22]
  wire  n123_I0; // @[Top.scala 75:22]
  wire  n123_I1; // @[Top.scala 75:22]
  wire  n123_O_t0b; // @[Top.scala 75:22]
  wire  n123_O_t1b; // @[Top.scala 75:22]
  wire  n124_valid_up; // @[Top.scala 79:22]
  wire  n124_valid_down; // @[Top.scala 79:22]
  wire  n124_I_t0b; // @[Top.scala 79:22]
  wire  n124_I_t1b; // @[Top.scala 79:22]
  wire  n124_O; // @[Top.scala 79:22]
  wire  InitialDelayCounter_2_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_2_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_2_valid_down; // @[Const.scala 11:33]
  wire  n127_valid_up; // @[Top.scala 83:22]
  wire  n127_valid_down; // @[Top.scala 83:22]
  wire [7:0] n127_I0; // @[Top.scala 83:22]
  wire [7:0] n127_I1; // @[Top.scala 83:22]
  wire [7:0] n127_O_t0b; // @[Top.scala 83:22]
  wire [7:0] n127_O_t1b; // @[Top.scala 83:22]
  wire  n128_valid_up; // @[Top.scala 87:22]
  wire  n128_valid_down; // @[Top.scala 87:22]
  wire  n128_I0; // @[Top.scala 87:22]
  wire [7:0] n128_I1_t0b; // @[Top.scala 87:22]
  wire [7:0] n128_I1_t1b; // @[Top.scala 87:22]
  wire  n128_O_t0b; // @[Top.scala 87:22]
  wire [7:0] n128_O_t1b_t0b; // @[Top.scala 87:22]
  wire [7:0] n128_O_t1b_t1b; // @[Top.scala 87:22]
  wire  n129_valid_up; // @[Top.scala 91:22]
  wire  n129_valid_down; // @[Top.scala 91:22]
  wire  n129_I_t0b; // @[Top.scala 91:22]
  wire [7:0] n129_I_t1b_t0b; // @[Top.scala 91:22]
  wire [7:0] n129_I_t1b_t1b; // @[Top.scala 91:22]
  wire [7:0] n129_O; // @[Top.scala 91:22]
  wire  InitialDelayCounter_3_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_3_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_3_valid_down; // @[Const.scala 11:33]
  wire  n132_valid_up; // @[Top.scala 95:22]
  wire  n132_valid_down; // @[Top.scala 95:22]
  wire [7:0] n132_I0; // @[Top.scala 95:22]
  wire [7:0] n132_I1; // @[Top.scala 95:22]
  wire [7:0] n132_O_t0b; // @[Top.scala 95:22]
  wire [7:0] n132_O_t1b; // @[Top.scala 95:22]
  wire  n133_valid_up; // @[Top.scala 99:22]
  wire  n133_valid_down; // @[Top.scala 99:22]
  wire [7:0] n133_I_t0b; // @[Top.scala 99:22]
  wire [7:0] n133_I_t1b; // @[Top.scala 99:22]
  wire [7:0] n133_O; // @[Top.scala 99:22]
  wire  n134_valid_up; // @[Top.scala 102:22]
  wire  n134_valid_down; // @[Top.scala 102:22]
  wire [7:0] n134_I0; // @[Top.scala 102:22]
  wire [7:0] n134_I1; // @[Top.scala 102:22]
  wire [7:0] n134_O_t0b; // @[Top.scala 102:22]
  wire [7:0] n134_O_t1b; // @[Top.scala 102:22]
  wire  n135_valid_up; // @[Top.scala 106:22]
  wire  n135_valid_down; // @[Top.scala 106:22]
  wire [7:0] n135_I_t0b; // @[Top.scala 106:22]
  wire [7:0] n135_I_t1b; // @[Top.scala 106:22]
  wire [7:0] n135_O; // @[Top.scala 106:22]
  InitialDelayCounter_1 InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  AtomTuple n113 ( // @[Top.scala 46:22]
    .valid_up(n113_valid_up),
    .valid_down(n113_valid_down),
    .I0(n113_I0),
    .I1(n113_I1),
    .O_t0b(n113_O_t0b),
    .O_t1b(n113_O_t1b)
  );
  Sub n114 ( // @[Top.scala 50:22]
    .valid_up(n114_valid_up),
    .valid_down(n114_valid_down),
    .I_t0b(n114_I_t0b),
    .I_t1b(n114_I_t1b),
    .O(n114_O)
  );
  AtomTuple n116 ( // @[Top.scala 53:22]
    .valid_up(n116_valid_up),
    .valid_down(n116_valid_down),
    .I0(n116_I0),
    .I1(n116_I1),
    .O_t0b(n116_O_t0b),
    .O_t1b(n116_O_t1b)
  );
  Lt n117 ( // @[Top.scala 57:22]
    .valid_up(n117_valid_up),
    .valid_down(n117_valid_down),
    .I_t0b(n117_I_t0b),
    .I_t1b(n117_I_t1b),
    .O(n117_O)
  );
  InitialDelayCounter_1 InitialDelayCounter_1 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_1_clock),
    .reset(InitialDelayCounter_1_reset),
    .valid_down(InitialDelayCounter_1_valid_down)
  );
  AtomTuple n118 ( // @[Top.scala 61:22]
    .valid_up(n118_valid_up),
    .valid_down(n118_valid_down),
    .I0(n118_I0),
    .I1(n118_I1),
    .O_t0b(n118_O_t0b),
    .O_t1b(n118_O_t1b)
  );
  Sub n119 ( // @[Top.scala 65:22]
    .valid_up(n119_valid_up),
    .valid_down(n119_valid_down),
    .I_t0b(n119_I_t0b),
    .I_t1b(n119_I_t1b),
    .O(n119_O)
  );
  AtomTuple n121 ( // @[Top.scala 68:22]
    .valid_up(n121_valid_up),
    .valid_down(n121_valid_down),
    .I0(n121_I0),
    .I1(n121_I1),
    .O_t0b(n121_O_t0b),
    .O_t1b(n121_O_t1b)
  );
  Lt n122 ( // @[Top.scala 72:22]
    .valid_up(n122_valid_up),
    .valid_down(n122_valid_down),
    .I_t0b(n122_I_t0b),
    .I_t1b(n122_I_t1b),
    .O(n122_O)
  );
  AtomTuple_6 n123 ( // @[Top.scala 75:22]
    .valid_up(n123_valid_up),
    .valid_down(n123_valid_down),
    .I0(n123_I0),
    .I1(n123_I1),
    .O_t0b(n123_O_t0b),
    .O_t1b(n123_O_t1b)
  );
  Or n124 ( // @[Top.scala 79:22]
    .valid_up(n124_valid_up),
    .valid_down(n124_valid_down),
    .I_t0b(n124_I_t0b),
    .I_t1b(n124_I_t1b),
    .O(n124_O)
  );
  InitialDelayCounter_1 InitialDelayCounter_2 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_2_clock),
    .reset(InitialDelayCounter_2_reset),
    .valid_down(InitialDelayCounter_2_valid_down)
  );
  AtomTuple n127 ( // @[Top.scala 83:22]
    .valid_up(n127_valid_up),
    .valid_down(n127_valid_down),
    .I0(n127_I0),
    .I1(n127_I1),
    .O_t0b(n127_O_t0b),
    .O_t1b(n127_O_t1b)
  );
  AtomTuple_8 n128 ( // @[Top.scala 87:22]
    .valid_up(n128_valid_up),
    .valid_down(n128_valid_down),
    .I0(n128_I0),
    .I1_t0b(n128_I1_t0b),
    .I1_t1b(n128_I1_t1b),
    .O_t0b(n128_O_t0b),
    .O_t1b_t0b(n128_O_t1b_t0b),
    .O_t1b_t1b(n128_O_t1b_t1b)
  );
  If n129 ( // @[Top.scala 91:22]
    .valid_up(n129_valid_up),
    .valid_down(n129_valid_down),
    .I_t0b(n129_I_t0b),
    .I_t1b_t0b(n129_I_t1b_t0b),
    .I_t1b_t1b(n129_I_t1b_t1b),
    .O(n129_O)
  );
  InitialDelayCounter_1 InitialDelayCounter_3 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_3_clock),
    .reset(InitialDelayCounter_3_reset),
    .valid_down(InitialDelayCounter_3_valid_down)
  );
  AtomTuple n132 ( // @[Top.scala 95:22]
    .valid_up(n132_valid_up),
    .valid_down(n132_valid_down),
    .I0(n132_I0),
    .I1(n132_I1),
    .O_t0b(n132_O_t0b),
    .O_t1b(n132_O_t1b)
  );
  RShift n133 ( // @[Top.scala 99:22]
    .valid_up(n133_valid_up),
    .valid_down(n133_valid_down),
    .I_t0b(n133_I_t0b),
    .I_t1b(n133_I_t1b),
    .O(n133_O)
  );
  AtomTuple n134 ( // @[Top.scala 102:22]
    .valid_up(n134_valid_up),
    .valid_down(n134_valid_down),
    .I0(n134_I0),
    .I1(n134_I1),
    .O_t0b(n134_O_t0b),
    .O_t1b(n134_O_t1b)
  );
  Add n135 ( // @[Top.scala 106:22]
    .valid_up(n135_valid_up),
    .valid_down(n135_valid_down),
    .I_t0b(n135_I_t0b),
    .I_t1b(n135_I_t1b),
    .O(n135_O)
  );
  assign valid_down = n135_valid_down; // @[Top.scala 110:16]
  assign O = n135_O; // @[Top.scala 109:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n113_valid_up = valid_up; // @[Top.scala 49:19]
  assign n113_I0 = I0; // @[Top.scala 47:13]
  assign n113_I1 = I1; // @[Top.scala 48:13]
  assign n114_valid_up = n113_valid_down; // @[Top.scala 52:19]
  assign n114_I_t0b = n113_O_t0b; // @[Top.scala 51:12]
  assign n114_I_t1b = n113_O_t1b; // @[Top.scala 51:12]
  assign n116_valid_up = InitialDelayCounter_valid_down & n114_valid_down; // @[Top.scala 56:19]
  assign n116_I0 = 8'hf; // @[Top.scala 54:13]
  assign n116_I1 = n114_O; // @[Top.scala 55:13]
  assign n117_valid_up = n116_valid_down; // @[Top.scala 59:19]
  assign n117_I_t0b = n116_O_t0b; // @[Top.scala 58:12]
  assign n117_I_t1b = n116_O_t1b; // @[Top.scala 58:12]
  assign InitialDelayCounter_1_clock = clock;
  assign InitialDelayCounter_1_reset = reset;
  assign n118_valid_up = valid_up; // @[Top.scala 64:19]
  assign n118_I0 = I1; // @[Top.scala 62:13]
  assign n118_I1 = I0; // @[Top.scala 63:13]
  assign n119_valid_up = n118_valid_down; // @[Top.scala 67:19]
  assign n119_I_t0b = n118_O_t0b; // @[Top.scala 66:12]
  assign n119_I_t1b = n118_O_t1b; // @[Top.scala 66:12]
  assign n121_valid_up = InitialDelayCounter_1_valid_down & n119_valid_down; // @[Top.scala 71:19]
  assign n121_I0 = 8'hf; // @[Top.scala 69:13]
  assign n121_I1 = n119_O; // @[Top.scala 70:13]
  assign n122_valid_up = n121_valid_down; // @[Top.scala 74:19]
  assign n122_I_t0b = n121_O_t0b; // @[Top.scala 73:12]
  assign n122_I_t1b = n121_O_t1b; // @[Top.scala 73:12]
  assign n123_valid_up = n117_valid_down & n122_valid_down; // @[Top.scala 78:19]
  assign n123_I0 = n117_O[0]; // @[Top.scala 76:13]
  assign n123_I1 = n122_O[0]; // @[Top.scala 77:13]
  assign n124_valid_up = n123_valid_down; // @[Top.scala 81:19]
  assign n124_I_t0b = n123_O_t0b; // @[Top.scala 80:12]
  assign n124_I_t1b = n123_O_t1b; // @[Top.scala 80:12]
  assign InitialDelayCounter_2_clock = clock;
  assign InitialDelayCounter_2_reset = reset;
  assign n127_valid_up = n119_valid_down & InitialDelayCounter_2_valid_down; // @[Top.scala 86:19]
  assign n127_I0 = n119_O; // @[Top.scala 84:13]
  assign n127_I1 = 8'h0; // @[Top.scala 85:13]
  assign n128_valid_up = n124_valid_down & n127_valid_down; // @[Top.scala 90:19]
  assign n128_I0 = n124_O; // @[Top.scala 88:13]
  assign n128_I1_t0b = n127_O_t0b; // @[Top.scala 89:13]
  assign n128_I1_t1b = n127_O_t1b; // @[Top.scala 89:13]
  assign n129_valid_up = n128_valid_down; // @[Top.scala 93:19]
  assign n129_I_t0b = n128_O_t0b; // @[Top.scala 92:12]
  assign n129_I_t1b_t0b = n128_O_t1b_t0b; // @[Top.scala 92:12]
  assign n129_I_t1b_t1b = n128_O_t1b_t1b; // @[Top.scala 92:12]
  assign InitialDelayCounter_3_clock = clock;
  assign InitialDelayCounter_3_reset = reset;
  assign n132_valid_up = n129_valid_down & InitialDelayCounter_3_valid_down; // @[Top.scala 98:19]
  assign n132_I0 = n129_O; // @[Top.scala 96:13]
  assign n132_I1 = 8'h2; // @[Top.scala 97:13]
  assign n133_valid_up = n132_valid_down; // @[Top.scala 101:19]
  assign n133_I_t0b = n132_O_t0b; // @[Top.scala 100:12]
  assign n133_I_t1b = n132_O_t1b; // @[Top.scala 100:12]
  assign n134_valid_up = valid_up & n133_valid_down; // @[Top.scala 105:19]
  assign n134_I0 = I1; // @[Top.scala 103:13]
  assign n134_I1 = n133_O; // @[Top.scala 104:13]
  assign n135_valid_up = n134_valid_down; // @[Top.scala 108:19]
  assign n135_I_t0b = n134_O_t0b; // @[Top.scala 107:12]
  assign n135_I_t1b = n134_O_t1b; // @[Top.scala 107:12]
endmodule
module Map2S_12(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I0_2,
  input  [7:0] I0_3,
  input  [7:0] I0_4,
  input  [7:0] I0_5,
  input  [7:0] I0_6,
  input  [7:0] I0_7,
  input  [7:0] I0_8,
  input  [7:0] I0_9,
  input  [7:0] I0_10,
  input  [7:0] I0_11,
  input  [7:0] I0_12,
  input  [7:0] I0_13,
  input  [7:0] I0_14,
  input  [7:0] I0_15,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  input  [7:0] I1_3,
  input  [7:0] I1_4,
  input  [7:0] I1_5,
  input  [7:0] I1_6,
  input  [7:0] I1_7,
  input  [7:0] I1_8,
  input  [7:0] I1_9,
  input  [7:0] I1_10,
  input  [7:0] I1_11,
  input  [7:0] I1_12,
  input  [7:0] I1_13,
  input  [7:0] I1_14,
  input  [7:0] I1_15,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15
);
  wire  fst_op_clock; // @[Map2S.scala 9:22]
  wire  fst_op_reset; // @[Map2S.scala 9:22]
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O; // @[Map2S.scala 9:22]
  wire  other_ops_0_clock; // @[Map2S.scala 10:86]
  wire  other_ops_0_reset; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O; // @[Map2S.scala 10:86]
  wire  other_ops_1_clock; // @[Map2S.scala 10:86]
  wire  other_ops_1_reset; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O; // @[Map2S.scala 10:86]
  wire  other_ops_2_clock; // @[Map2S.scala 10:86]
  wire  other_ops_2_reset; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O; // @[Map2S.scala 10:86]
  wire  other_ops_3_clock; // @[Map2S.scala 10:86]
  wire  other_ops_3_reset; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O; // @[Map2S.scala 10:86]
  wire  other_ops_4_clock; // @[Map2S.scala 10:86]
  wire  other_ops_4_reset; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O; // @[Map2S.scala 10:86]
  wire  other_ops_5_clock; // @[Map2S.scala 10:86]
  wire  other_ops_5_reset; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O; // @[Map2S.scala 10:86]
  wire  other_ops_6_clock; // @[Map2S.scala 10:86]
  wire  other_ops_6_reset; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O; // @[Map2S.scala 10:86]
  wire  other_ops_7_clock; // @[Map2S.scala 10:86]
  wire  other_ops_7_reset; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O; // @[Map2S.scala 10:86]
  wire  other_ops_8_clock; // @[Map2S.scala 10:86]
  wire  other_ops_8_reset; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O; // @[Map2S.scala 10:86]
  wire  other_ops_9_clock; // @[Map2S.scala 10:86]
  wire  other_ops_9_reset; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O; // @[Map2S.scala 10:86]
  wire  other_ops_10_clock; // @[Map2S.scala 10:86]
  wire  other_ops_10_reset; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O; // @[Map2S.scala 10:86]
  wire  other_ops_11_clock; // @[Map2S.scala 10:86]
  wire  other_ops_11_reset; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O; // @[Map2S.scala 10:86]
  wire  other_ops_12_clock; // @[Map2S.scala 10:86]
  wire  other_ops_12_reset; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O; // @[Map2S.scala 10:86]
  wire  other_ops_13_clock; // @[Map2S.scala 10:86]
  wire  other_ops_13_reset; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O; // @[Map2S.scala 10:86]
  wire  other_ops_14_clock; // @[Map2S.scala 10:86]
  wire  other_ops_14_reset; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  Module_1 fst_op ( // @[Map2S.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O(fst_op_O)
  );
  Module_1 other_ops_0 ( // @[Map2S.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O(other_ops_0_O)
  );
  Module_1 other_ops_1 ( // @[Map2S.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O(other_ops_1_O)
  );
  Module_1 other_ops_2 ( // @[Map2S.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0(other_ops_2_I0),
    .I1(other_ops_2_I1),
    .O(other_ops_2_O)
  );
  Module_1 other_ops_3 ( // @[Map2S.scala 10:86]
    .clock(other_ops_3_clock),
    .reset(other_ops_3_reset),
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0(other_ops_3_I0),
    .I1(other_ops_3_I1),
    .O(other_ops_3_O)
  );
  Module_1 other_ops_4 ( // @[Map2S.scala 10:86]
    .clock(other_ops_4_clock),
    .reset(other_ops_4_reset),
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0(other_ops_4_I0),
    .I1(other_ops_4_I1),
    .O(other_ops_4_O)
  );
  Module_1 other_ops_5 ( // @[Map2S.scala 10:86]
    .clock(other_ops_5_clock),
    .reset(other_ops_5_reset),
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0(other_ops_5_I0),
    .I1(other_ops_5_I1),
    .O(other_ops_5_O)
  );
  Module_1 other_ops_6 ( // @[Map2S.scala 10:86]
    .clock(other_ops_6_clock),
    .reset(other_ops_6_reset),
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0(other_ops_6_I0),
    .I1(other_ops_6_I1),
    .O(other_ops_6_O)
  );
  Module_1 other_ops_7 ( // @[Map2S.scala 10:86]
    .clock(other_ops_7_clock),
    .reset(other_ops_7_reset),
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0(other_ops_7_I0),
    .I1(other_ops_7_I1),
    .O(other_ops_7_O)
  );
  Module_1 other_ops_8 ( // @[Map2S.scala 10:86]
    .clock(other_ops_8_clock),
    .reset(other_ops_8_reset),
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0(other_ops_8_I0),
    .I1(other_ops_8_I1),
    .O(other_ops_8_O)
  );
  Module_1 other_ops_9 ( // @[Map2S.scala 10:86]
    .clock(other_ops_9_clock),
    .reset(other_ops_9_reset),
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0(other_ops_9_I0),
    .I1(other_ops_9_I1),
    .O(other_ops_9_O)
  );
  Module_1 other_ops_10 ( // @[Map2S.scala 10:86]
    .clock(other_ops_10_clock),
    .reset(other_ops_10_reset),
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0(other_ops_10_I0),
    .I1(other_ops_10_I1),
    .O(other_ops_10_O)
  );
  Module_1 other_ops_11 ( // @[Map2S.scala 10:86]
    .clock(other_ops_11_clock),
    .reset(other_ops_11_reset),
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0(other_ops_11_I0),
    .I1(other_ops_11_I1),
    .O(other_ops_11_O)
  );
  Module_1 other_ops_12 ( // @[Map2S.scala 10:86]
    .clock(other_ops_12_clock),
    .reset(other_ops_12_reset),
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0(other_ops_12_I0),
    .I1(other_ops_12_I1),
    .O(other_ops_12_O)
  );
  Module_1 other_ops_13 ( // @[Map2S.scala 10:86]
    .clock(other_ops_13_clock),
    .reset(other_ops_13_reset),
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0(other_ops_13_I0),
    .I1(other_ops_13_I1),
    .O(other_ops_13_O)
  );
  Module_1 other_ops_14 ( // @[Map2S.scala 10:86]
    .clock(other_ops_14_clock),
    .reset(other_ops_14_reset),
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0(other_ops_14_I0),
    .I1(other_ops_14_I1),
    .O(other_ops_14_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0 = fst_op_O; // @[Map2S.scala 19:8]
  assign O_1 = other_ops_0_O; // @[Map2S.scala 24:12]
  assign O_2 = other_ops_1_O; // @[Map2S.scala 24:12]
  assign O_3 = other_ops_2_O; // @[Map2S.scala 24:12]
  assign O_4 = other_ops_3_O; // @[Map2S.scala 24:12]
  assign O_5 = other_ops_4_O; // @[Map2S.scala 24:12]
  assign O_6 = other_ops_5_O; // @[Map2S.scala 24:12]
  assign O_7 = other_ops_6_O; // @[Map2S.scala 24:12]
  assign O_8 = other_ops_7_O; // @[Map2S.scala 24:12]
  assign O_9 = other_ops_8_O; // @[Map2S.scala 24:12]
  assign O_10 = other_ops_9_O; // @[Map2S.scala 24:12]
  assign O_11 = other_ops_10_O; // @[Map2S.scala 24:12]
  assign O_12 = other_ops_11_O; // @[Map2S.scala 24:12]
  assign O_13 = other_ops_12_O; // @[Map2S.scala 24:12]
  assign O_14 = other_ops_13_O; // @[Map2S.scala 24:12]
  assign O_15 = other_ops_14_O; // @[Map2S.scala 24:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_0_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_1_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_2_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0 = I0_3; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
  assign other_ops_3_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_3_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0 = I0_4; // @[Map2S.scala 22:43]
  assign other_ops_3_I1 = I1_4; // @[Map2S.scala 23:43]
  assign other_ops_4_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_4_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0 = I0_5; // @[Map2S.scala 22:43]
  assign other_ops_4_I1 = I1_5; // @[Map2S.scala 23:43]
  assign other_ops_5_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_5_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0 = I0_6; // @[Map2S.scala 22:43]
  assign other_ops_5_I1 = I1_6; // @[Map2S.scala 23:43]
  assign other_ops_6_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_6_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0 = I0_7; // @[Map2S.scala 22:43]
  assign other_ops_6_I1 = I1_7; // @[Map2S.scala 23:43]
  assign other_ops_7_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_7_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0 = I0_8; // @[Map2S.scala 22:43]
  assign other_ops_7_I1 = I1_8; // @[Map2S.scala 23:43]
  assign other_ops_8_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_8_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0 = I0_9; // @[Map2S.scala 22:43]
  assign other_ops_8_I1 = I1_9; // @[Map2S.scala 23:43]
  assign other_ops_9_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_9_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0 = I0_10; // @[Map2S.scala 22:43]
  assign other_ops_9_I1 = I1_10; // @[Map2S.scala 23:43]
  assign other_ops_10_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_10_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0 = I0_11; // @[Map2S.scala 22:43]
  assign other_ops_10_I1 = I1_11; // @[Map2S.scala 23:43]
  assign other_ops_11_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_11_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0 = I0_12; // @[Map2S.scala 22:43]
  assign other_ops_11_I1 = I1_12; // @[Map2S.scala 23:43]
  assign other_ops_12_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_12_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0 = I0_13; // @[Map2S.scala 22:43]
  assign other_ops_12_I1 = I1_13; // @[Map2S.scala 23:43]
  assign other_ops_13_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_13_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0 = I0_14; // @[Map2S.scala 22:43]
  assign other_ops_13_I1 = I1_14; // @[Map2S.scala 23:43]
  assign other_ops_14_clock = clock; // @[Map2S.scala 10:86]
  assign other_ops_14_reset = reset; // @[Map2S.scala 10:86]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0 = I0_15; // @[Map2S.scala 22:43]
  assign other_ops_14_I1 = I1_15; // @[Map2S.scala 23:43]
endmodule
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  input  [7:0] I_4,
  input  [7:0] I_5,
  input  [7:0] I_6,
  input  [7:0] I_7,
  input  [7:0] I_8,
  input  [7:0] I_9,
  input  [7:0] I_10,
  input  [7:0] I_11,
  input  [7:0] I_12,
  input  [7:0] I_13,
  input  [7:0] I_14,
  input  [7:0] I_15,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15
);
  wire  n1_clock; // @[Top.scala 116:20]
  wire  n1_reset; // @[Top.scala 116:20]
  wire  n1_valid_up; // @[Top.scala 116:20]
  wire  n1_valid_down; // @[Top.scala 116:20]
  wire [7:0] n1_I_0; // @[Top.scala 116:20]
  wire [7:0] n1_I_1; // @[Top.scala 116:20]
  wire [7:0] n1_I_2; // @[Top.scala 116:20]
  wire [7:0] n1_I_3; // @[Top.scala 116:20]
  wire [7:0] n1_I_4; // @[Top.scala 116:20]
  wire [7:0] n1_I_5; // @[Top.scala 116:20]
  wire [7:0] n1_I_6; // @[Top.scala 116:20]
  wire [7:0] n1_I_7; // @[Top.scala 116:20]
  wire [7:0] n1_I_8; // @[Top.scala 116:20]
  wire [7:0] n1_I_9; // @[Top.scala 116:20]
  wire [7:0] n1_I_10; // @[Top.scala 116:20]
  wire [7:0] n1_I_11; // @[Top.scala 116:20]
  wire [7:0] n1_I_12; // @[Top.scala 116:20]
  wire [7:0] n1_I_13; // @[Top.scala 116:20]
  wire [7:0] n1_I_14; // @[Top.scala 116:20]
  wire [7:0] n1_I_15; // @[Top.scala 116:20]
  wire [7:0] n1_O_0; // @[Top.scala 116:20]
  wire [7:0] n1_O_1; // @[Top.scala 116:20]
  wire [7:0] n1_O_2; // @[Top.scala 116:20]
  wire [7:0] n1_O_3; // @[Top.scala 116:20]
  wire [7:0] n1_O_4; // @[Top.scala 116:20]
  wire [7:0] n1_O_5; // @[Top.scala 116:20]
  wire [7:0] n1_O_6; // @[Top.scala 116:20]
  wire [7:0] n1_O_7; // @[Top.scala 116:20]
  wire [7:0] n1_O_8; // @[Top.scala 116:20]
  wire [7:0] n1_O_9; // @[Top.scala 116:20]
  wire [7:0] n1_O_10; // @[Top.scala 116:20]
  wire [7:0] n1_O_11; // @[Top.scala 116:20]
  wire [7:0] n1_O_12; // @[Top.scala 116:20]
  wire [7:0] n1_O_13; // @[Top.scala 116:20]
  wire [7:0] n1_O_14; // @[Top.scala 116:20]
  wire [7:0] n1_O_15; // @[Top.scala 116:20]
  wire  n2_valid_up; // @[Top.scala 119:20]
  wire  n2_valid_down; // @[Top.scala 119:20]
  wire [7:0] n2_I_0; // @[Top.scala 119:20]
  wire [7:0] n2_I_1; // @[Top.scala 119:20]
  wire [7:0] n2_I_2; // @[Top.scala 119:20]
  wire [7:0] n2_I_3; // @[Top.scala 119:20]
  wire [7:0] n2_I_4; // @[Top.scala 119:20]
  wire [7:0] n2_I_5; // @[Top.scala 119:20]
  wire [7:0] n2_I_6; // @[Top.scala 119:20]
  wire [7:0] n2_I_7; // @[Top.scala 119:20]
  wire [7:0] n2_I_8; // @[Top.scala 119:20]
  wire [7:0] n2_I_9; // @[Top.scala 119:20]
  wire [7:0] n2_I_10; // @[Top.scala 119:20]
  wire [7:0] n2_I_11; // @[Top.scala 119:20]
  wire [7:0] n2_I_12; // @[Top.scala 119:20]
  wire [7:0] n2_I_13; // @[Top.scala 119:20]
  wire [7:0] n2_I_14; // @[Top.scala 119:20]
  wire [7:0] n2_I_15; // @[Top.scala 119:20]
  wire [7:0] n2_O_0; // @[Top.scala 119:20]
  wire [7:0] n2_O_1; // @[Top.scala 119:20]
  wire [7:0] n2_O_2; // @[Top.scala 119:20]
  wire [7:0] n2_O_3; // @[Top.scala 119:20]
  wire [7:0] n2_O_4; // @[Top.scala 119:20]
  wire [7:0] n2_O_5; // @[Top.scala 119:20]
  wire [7:0] n2_O_6; // @[Top.scala 119:20]
  wire [7:0] n2_O_7; // @[Top.scala 119:20]
  wire [7:0] n2_O_8; // @[Top.scala 119:20]
  wire [7:0] n2_O_9; // @[Top.scala 119:20]
  wire [7:0] n2_O_10; // @[Top.scala 119:20]
  wire [7:0] n2_O_11; // @[Top.scala 119:20]
  wire [7:0] n2_O_12; // @[Top.scala 119:20]
  wire [7:0] n2_O_13; // @[Top.scala 119:20]
  wire [7:0] n2_O_14; // @[Top.scala 119:20]
  wire [7:0] n2_O_15; // @[Top.scala 119:20]
  wire  n3_valid_up; // @[Top.scala 122:20]
  wire  n3_valid_down; // @[Top.scala 122:20]
  wire [7:0] n3_I_0; // @[Top.scala 122:20]
  wire [7:0] n3_I_1; // @[Top.scala 122:20]
  wire [7:0] n3_I_2; // @[Top.scala 122:20]
  wire [7:0] n3_I_3; // @[Top.scala 122:20]
  wire [7:0] n3_I_4; // @[Top.scala 122:20]
  wire [7:0] n3_I_5; // @[Top.scala 122:20]
  wire [7:0] n3_I_6; // @[Top.scala 122:20]
  wire [7:0] n3_I_7; // @[Top.scala 122:20]
  wire [7:0] n3_I_8; // @[Top.scala 122:20]
  wire [7:0] n3_I_9; // @[Top.scala 122:20]
  wire [7:0] n3_I_10; // @[Top.scala 122:20]
  wire [7:0] n3_I_11; // @[Top.scala 122:20]
  wire [7:0] n3_I_12; // @[Top.scala 122:20]
  wire [7:0] n3_I_13; // @[Top.scala 122:20]
  wire [7:0] n3_I_14; // @[Top.scala 122:20]
  wire [7:0] n3_I_15; // @[Top.scala 122:20]
  wire [7:0] n3_O_0; // @[Top.scala 122:20]
  wire [7:0] n3_O_1; // @[Top.scala 122:20]
  wire [7:0] n3_O_2; // @[Top.scala 122:20]
  wire [7:0] n3_O_3; // @[Top.scala 122:20]
  wire [7:0] n3_O_4; // @[Top.scala 122:20]
  wire [7:0] n3_O_5; // @[Top.scala 122:20]
  wire [7:0] n3_O_6; // @[Top.scala 122:20]
  wire [7:0] n3_O_7; // @[Top.scala 122:20]
  wire [7:0] n3_O_8; // @[Top.scala 122:20]
  wire [7:0] n3_O_9; // @[Top.scala 122:20]
  wire [7:0] n3_O_10; // @[Top.scala 122:20]
  wire [7:0] n3_O_11; // @[Top.scala 122:20]
  wire [7:0] n3_O_12; // @[Top.scala 122:20]
  wire [7:0] n3_O_13; // @[Top.scala 122:20]
  wire [7:0] n3_O_14; // @[Top.scala 122:20]
  wire [7:0] n3_O_15; // @[Top.scala 122:20]
  wire  n4_valid_up; // @[Top.scala 125:20]
  wire  n4_valid_down; // @[Top.scala 125:20]
  wire [7:0] n4_I_0; // @[Top.scala 125:20]
  wire [7:0] n4_I_1; // @[Top.scala 125:20]
  wire [7:0] n4_I_2; // @[Top.scala 125:20]
  wire [7:0] n4_I_3; // @[Top.scala 125:20]
  wire [7:0] n4_I_4; // @[Top.scala 125:20]
  wire [7:0] n4_I_5; // @[Top.scala 125:20]
  wire [7:0] n4_I_6; // @[Top.scala 125:20]
  wire [7:0] n4_I_7; // @[Top.scala 125:20]
  wire [7:0] n4_I_8; // @[Top.scala 125:20]
  wire [7:0] n4_I_9; // @[Top.scala 125:20]
  wire [7:0] n4_I_10; // @[Top.scala 125:20]
  wire [7:0] n4_I_11; // @[Top.scala 125:20]
  wire [7:0] n4_I_12; // @[Top.scala 125:20]
  wire [7:0] n4_I_13; // @[Top.scala 125:20]
  wire [7:0] n4_I_14; // @[Top.scala 125:20]
  wire [7:0] n4_I_15; // @[Top.scala 125:20]
  wire [7:0] n4_O_0; // @[Top.scala 125:20]
  wire [7:0] n4_O_1; // @[Top.scala 125:20]
  wire [7:0] n4_O_2; // @[Top.scala 125:20]
  wire [7:0] n4_O_3; // @[Top.scala 125:20]
  wire [7:0] n4_O_4; // @[Top.scala 125:20]
  wire [7:0] n4_O_5; // @[Top.scala 125:20]
  wire [7:0] n4_O_6; // @[Top.scala 125:20]
  wire [7:0] n4_O_7; // @[Top.scala 125:20]
  wire [7:0] n4_O_8; // @[Top.scala 125:20]
  wire [7:0] n4_O_9; // @[Top.scala 125:20]
  wire [7:0] n4_O_10; // @[Top.scala 125:20]
  wire [7:0] n4_O_11; // @[Top.scala 125:20]
  wire [7:0] n4_O_12; // @[Top.scala 125:20]
  wire [7:0] n4_O_13; // @[Top.scala 125:20]
  wire [7:0] n4_O_14; // @[Top.scala 125:20]
  wire [7:0] n4_O_15; // @[Top.scala 125:20]
  wire  n5_valid_up; // @[Top.scala 128:20]
  wire  n5_valid_down; // @[Top.scala 128:20]
  wire [7:0] n5_I_0; // @[Top.scala 128:20]
  wire [7:0] n5_I_1; // @[Top.scala 128:20]
  wire [7:0] n5_I_2; // @[Top.scala 128:20]
  wire [7:0] n5_I_3; // @[Top.scala 128:20]
  wire [7:0] n5_I_4; // @[Top.scala 128:20]
  wire [7:0] n5_I_5; // @[Top.scala 128:20]
  wire [7:0] n5_I_6; // @[Top.scala 128:20]
  wire [7:0] n5_I_7; // @[Top.scala 128:20]
  wire [7:0] n5_I_8; // @[Top.scala 128:20]
  wire [7:0] n5_I_9; // @[Top.scala 128:20]
  wire [7:0] n5_I_10; // @[Top.scala 128:20]
  wire [7:0] n5_I_11; // @[Top.scala 128:20]
  wire [7:0] n5_I_12; // @[Top.scala 128:20]
  wire [7:0] n5_I_13; // @[Top.scala 128:20]
  wire [7:0] n5_I_14; // @[Top.scala 128:20]
  wire [7:0] n5_I_15; // @[Top.scala 128:20]
  wire [7:0] n5_O_0; // @[Top.scala 128:20]
  wire [7:0] n5_O_1; // @[Top.scala 128:20]
  wire [7:0] n5_O_2; // @[Top.scala 128:20]
  wire [7:0] n5_O_3; // @[Top.scala 128:20]
  wire [7:0] n5_O_4; // @[Top.scala 128:20]
  wire [7:0] n5_O_5; // @[Top.scala 128:20]
  wire [7:0] n5_O_6; // @[Top.scala 128:20]
  wire [7:0] n5_O_7; // @[Top.scala 128:20]
  wire [7:0] n5_O_8; // @[Top.scala 128:20]
  wire [7:0] n5_O_9; // @[Top.scala 128:20]
  wire [7:0] n5_O_10; // @[Top.scala 128:20]
  wire [7:0] n5_O_11; // @[Top.scala 128:20]
  wire [7:0] n5_O_12; // @[Top.scala 128:20]
  wire [7:0] n5_O_13; // @[Top.scala 128:20]
  wire [7:0] n5_O_14; // @[Top.scala 128:20]
  wire [7:0] n5_O_15; // @[Top.scala 128:20]
  wire  n6_valid_up; // @[Top.scala 131:20]
  wire  n6_valid_down; // @[Top.scala 131:20]
  wire [7:0] n6_I0_0; // @[Top.scala 131:20]
  wire [7:0] n6_I0_1; // @[Top.scala 131:20]
  wire [7:0] n6_I0_2; // @[Top.scala 131:20]
  wire [7:0] n6_I0_3; // @[Top.scala 131:20]
  wire [7:0] n6_I0_4; // @[Top.scala 131:20]
  wire [7:0] n6_I0_5; // @[Top.scala 131:20]
  wire [7:0] n6_I0_6; // @[Top.scala 131:20]
  wire [7:0] n6_I0_7; // @[Top.scala 131:20]
  wire [7:0] n6_I0_8; // @[Top.scala 131:20]
  wire [7:0] n6_I0_9; // @[Top.scala 131:20]
  wire [7:0] n6_I0_10; // @[Top.scala 131:20]
  wire [7:0] n6_I0_11; // @[Top.scala 131:20]
  wire [7:0] n6_I0_12; // @[Top.scala 131:20]
  wire [7:0] n6_I0_13; // @[Top.scala 131:20]
  wire [7:0] n6_I0_14; // @[Top.scala 131:20]
  wire [7:0] n6_I0_15; // @[Top.scala 131:20]
  wire [7:0] n6_I1_0; // @[Top.scala 131:20]
  wire [7:0] n6_I1_1; // @[Top.scala 131:20]
  wire [7:0] n6_I1_2; // @[Top.scala 131:20]
  wire [7:0] n6_I1_3; // @[Top.scala 131:20]
  wire [7:0] n6_I1_4; // @[Top.scala 131:20]
  wire [7:0] n6_I1_5; // @[Top.scala 131:20]
  wire [7:0] n6_I1_6; // @[Top.scala 131:20]
  wire [7:0] n6_I1_7; // @[Top.scala 131:20]
  wire [7:0] n6_I1_8; // @[Top.scala 131:20]
  wire [7:0] n6_I1_9; // @[Top.scala 131:20]
  wire [7:0] n6_I1_10; // @[Top.scala 131:20]
  wire [7:0] n6_I1_11; // @[Top.scala 131:20]
  wire [7:0] n6_I1_12; // @[Top.scala 131:20]
  wire [7:0] n6_I1_13; // @[Top.scala 131:20]
  wire [7:0] n6_I1_14; // @[Top.scala 131:20]
  wire [7:0] n6_I1_15; // @[Top.scala 131:20]
  wire [7:0] n6_O_0_0; // @[Top.scala 131:20]
  wire [7:0] n6_O_0_1; // @[Top.scala 131:20]
  wire [7:0] n6_O_1_0; // @[Top.scala 131:20]
  wire [7:0] n6_O_1_1; // @[Top.scala 131:20]
  wire [7:0] n6_O_2_0; // @[Top.scala 131:20]
  wire [7:0] n6_O_2_1; // @[Top.scala 131:20]
  wire [7:0] n6_O_3_0; // @[Top.scala 131:20]
  wire [7:0] n6_O_3_1; // @[Top.scala 131:20]
  wire [7:0] n6_O_4_0; // @[Top.scala 131:20]
  wire [7:0] n6_O_4_1; // @[Top.scala 131:20]
  wire [7:0] n6_O_5_0; // @[Top.scala 131:20]
  wire [7:0] n6_O_5_1; // @[Top.scala 131:20]
  wire [7:0] n6_O_6_0; // @[Top.scala 131:20]
  wire [7:0] n6_O_6_1; // @[Top.scala 131:20]
  wire [7:0] n6_O_7_0; // @[Top.scala 131:20]
  wire [7:0] n6_O_7_1; // @[Top.scala 131:20]
  wire [7:0] n6_O_8_0; // @[Top.scala 131:20]
  wire [7:0] n6_O_8_1; // @[Top.scala 131:20]
  wire [7:0] n6_O_9_0; // @[Top.scala 131:20]
  wire [7:0] n6_O_9_1; // @[Top.scala 131:20]
  wire [7:0] n6_O_10_0; // @[Top.scala 131:20]
  wire [7:0] n6_O_10_1; // @[Top.scala 131:20]
  wire [7:0] n6_O_11_0; // @[Top.scala 131:20]
  wire [7:0] n6_O_11_1; // @[Top.scala 131:20]
  wire [7:0] n6_O_12_0; // @[Top.scala 131:20]
  wire [7:0] n6_O_12_1; // @[Top.scala 131:20]
  wire [7:0] n6_O_13_0; // @[Top.scala 131:20]
  wire [7:0] n6_O_13_1; // @[Top.scala 131:20]
  wire [7:0] n6_O_14_0; // @[Top.scala 131:20]
  wire [7:0] n6_O_14_1; // @[Top.scala 131:20]
  wire [7:0] n6_O_15_0; // @[Top.scala 131:20]
  wire [7:0] n6_O_15_1; // @[Top.scala 131:20]
  wire  n10_valid_up; // @[Top.scala 135:21]
  wire  n10_valid_down; // @[Top.scala 135:21]
  wire [7:0] n10_I0_0_0; // @[Top.scala 135:21]
  wire [7:0] n10_I0_0_1; // @[Top.scala 135:21]
  wire [7:0] n10_I0_1_0; // @[Top.scala 135:21]
  wire [7:0] n10_I0_1_1; // @[Top.scala 135:21]
  wire [7:0] n10_I0_2_0; // @[Top.scala 135:21]
  wire [7:0] n10_I0_2_1; // @[Top.scala 135:21]
  wire [7:0] n10_I0_3_0; // @[Top.scala 135:21]
  wire [7:0] n10_I0_3_1; // @[Top.scala 135:21]
  wire [7:0] n10_I0_4_0; // @[Top.scala 135:21]
  wire [7:0] n10_I0_4_1; // @[Top.scala 135:21]
  wire [7:0] n10_I0_5_0; // @[Top.scala 135:21]
  wire [7:0] n10_I0_5_1; // @[Top.scala 135:21]
  wire [7:0] n10_I0_6_0; // @[Top.scala 135:21]
  wire [7:0] n10_I0_6_1; // @[Top.scala 135:21]
  wire [7:0] n10_I0_7_0; // @[Top.scala 135:21]
  wire [7:0] n10_I0_7_1; // @[Top.scala 135:21]
  wire [7:0] n10_I0_8_0; // @[Top.scala 135:21]
  wire [7:0] n10_I0_8_1; // @[Top.scala 135:21]
  wire [7:0] n10_I0_9_0; // @[Top.scala 135:21]
  wire [7:0] n10_I0_9_1; // @[Top.scala 135:21]
  wire [7:0] n10_I0_10_0; // @[Top.scala 135:21]
  wire [7:0] n10_I0_10_1; // @[Top.scala 135:21]
  wire [7:0] n10_I0_11_0; // @[Top.scala 135:21]
  wire [7:0] n10_I0_11_1; // @[Top.scala 135:21]
  wire [7:0] n10_I0_12_0; // @[Top.scala 135:21]
  wire [7:0] n10_I0_12_1; // @[Top.scala 135:21]
  wire [7:0] n10_I0_13_0; // @[Top.scala 135:21]
  wire [7:0] n10_I0_13_1; // @[Top.scala 135:21]
  wire [7:0] n10_I0_14_0; // @[Top.scala 135:21]
  wire [7:0] n10_I0_14_1; // @[Top.scala 135:21]
  wire [7:0] n10_I0_15_0; // @[Top.scala 135:21]
  wire [7:0] n10_I0_15_1; // @[Top.scala 135:21]
  wire [7:0] n10_I1_0; // @[Top.scala 135:21]
  wire [7:0] n10_I1_1; // @[Top.scala 135:21]
  wire [7:0] n10_I1_2; // @[Top.scala 135:21]
  wire [7:0] n10_I1_3; // @[Top.scala 135:21]
  wire [7:0] n10_I1_4; // @[Top.scala 135:21]
  wire [7:0] n10_I1_5; // @[Top.scala 135:21]
  wire [7:0] n10_I1_6; // @[Top.scala 135:21]
  wire [7:0] n10_I1_7; // @[Top.scala 135:21]
  wire [7:0] n10_I1_8; // @[Top.scala 135:21]
  wire [7:0] n10_I1_9; // @[Top.scala 135:21]
  wire [7:0] n10_I1_10; // @[Top.scala 135:21]
  wire [7:0] n10_I1_11; // @[Top.scala 135:21]
  wire [7:0] n10_I1_12; // @[Top.scala 135:21]
  wire [7:0] n10_I1_13; // @[Top.scala 135:21]
  wire [7:0] n10_I1_14; // @[Top.scala 135:21]
  wire [7:0] n10_I1_15; // @[Top.scala 135:21]
  wire [7:0] n10_O_0_0; // @[Top.scala 135:21]
  wire [7:0] n10_O_0_1; // @[Top.scala 135:21]
  wire [7:0] n10_O_0_2; // @[Top.scala 135:21]
  wire [7:0] n10_O_1_0; // @[Top.scala 135:21]
  wire [7:0] n10_O_1_1; // @[Top.scala 135:21]
  wire [7:0] n10_O_1_2; // @[Top.scala 135:21]
  wire [7:0] n10_O_2_0; // @[Top.scala 135:21]
  wire [7:0] n10_O_2_1; // @[Top.scala 135:21]
  wire [7:0] n10_O_2_2; // @[Top.scala 135:21]
  wire [7:0] n10_O_3_0; // @[Top.scala 135:21]
  wire [7:0] n10_O_3_1; // @[Top.scala 135:21]
  wire [7:0] n10_O_3_2; // @[Top.scala 135:21]
  wire [7:0] n10_O_4_0; // @[Top.scala 135:21]
  wire [7:0] n10_O_4_1; // @[Top.scala 135:21]
  wire [7:0] n10_O_4_2; // @[Top.scala 135:21]
  wire [7:0] n10_O_5_0; // @[Top.scala 135:21]
  wire [7:0] n10_O_5_1; // @[Top.scala 135:21]
  wire [7:0] n10_O_5_2; // @[Top.scala 135:21]
  wire [7:0] n10_O_6_0; // @[Top.scala 135:21]
  wire [7:0] n10_O_6_1; // @[Top.scala 135:21]
  wire [7:0] n10_O_6_2; // @[Top.scala 135:21]
  wire [7:0] n10_O_7_0; // @[Top.scala 135:21]
  wire [7:0] n10_O_7_1; // @[Top.scala 135:21]
  wire [7:0] n10_O_7_2; // @[Top.scala 135:21]
  wire [7:0] n10_O_8_0; // @[Top.scala 135:21]
  wire [7:0] n10_O_8_1; // @[Top.scala 135:21]
  wire [7:0] n10_O_8_2; // @[Top.scala 135:21]
  wire [7:0] n10_O_9_0; // @[Top.scala 135:21]
  wire [7:0] n10_O_9_1; // @[Top.scala 135:21]
  wire [7:0] n10_O_9_2; // @[Top.scala 135:21]
  wire [7:0] n10_O_10_0; // @[Top.scala 135:21]
  wire [7:0] n10_O_10_1; // @[Top.scala 135:21]
  wire [7:0] n10_O_10_2; // @[Top.scala 135:21]
  wire [7:0] n10_O_11_0; // @[Top.scala 135:21]
  wire [7:0] n10_O_11_1; // @[Top.scala 135:21]
  wire [7:0] n10_O_11_2; // @[Top.scala 135:21]
  wire [7:0] n10_O_12_0; // @[Top.scala 135:21]
  wire [7:0] n10_O_12_1; // @[Top.scala 135:21]
  wire [7:0] n10_O_12_2; // @[Top.scala 135:21]
  wire [7:0] n10_O_13_0; // @[Top.scala 135:21]
  wire [7:0] n10_O_13_1; // @[Top.scala 135:21]
  wire [7:0] n10_O_13_2; // @[Top.scala 135:21]
  wire [7:0] n10_O_14_0; // @[Top.scala 135:21]
  wire [7:0] n10_O_14_1; // @[Top.scala 135:21]
  wire [7:0] n10_O_14_2; // @[Top.scala 135:21]
  wire [7:0] n10_O_15_0; // @[Top.scala 135:21]
  wire [7:0] n10_O_15_1; // @[Top.scala 135:21]
  wire [7:0] n10_O_15_2; // @[Top.scala 135:21]
  wire  n14_valid_up; // @[Top.scala 139:21]
  wire  n14_valid_down; // @[Top.scala 139:21]
  wire [7:0] n14_I_0_0; // @[Top.scala 139:21]
  wire [7:0] n14_I_0_1; // @[Top.scala 139:21]
  wire [7:0] n14_I_0_2; // @[Top.scala 139:21]
  wire [7:0] n14_I_1_0; // @[Top.scala 139:21]
  wire [7:0] n14_I_1_1; // @[Top.scala 139:21]
  wire [7:0] n14_I_1_2; // @[Top.scala 139:21]
  wire [7:0] n14_I_2_0; // @[Top.scala 139:21]
  wire [7:0] n14_I_2_1; // @[Top.scala 139:21]
  wire [7:0] n14_I_2_2; // @[Top.scala 139:21]
  wire [7:0] n14_I_3_0; // @[Top.scala 139:21]
  wire [7:0] n14_I_3_1; // @[Top.scala 139:21]
  wire [7:0] n14_I_3_2; // @[Top.scala 139:21]
  wire [7:0] n14_I_4_0; // @[Top.scala 139:21]
  wire [7:0] n14_I_4_1; // @[Top.scala 139:21]
  wire [7:0] n14_I_4_2; // @[Top.scala 139:21]
  wire [7:0] n14_I_5_0; // @[Top.scala 139:21]
  wire [7:0] n14_I_5_1; // @[Top.scala 139:21]
  wire [7:0] n14_I_5_2; // @[Top.scala 139:21]
  wire [7:0] n14_I_6_0; // @[Top.scala 139:21]
  wire [7:0] n14_I_6_1; // @[Top.scala 139:21]
  wire [7:0] n14_I_6_2; // @[Top.scala 139:21]
  wire [7:0] n14_I_7_0; // @[Top.scala 139:21]
  wire [7:0] n14_I_7_1; // @[Top.scala 139:21]
  wire [7:0] n14_I_7_2; // @[Top.scala 139:21]
  wire [7:0] n14_I_8_0; // @[Top.scala 139:21]
  wire [7:0] n14_I_8_1; // @[Top.scala 139:21]
  wire [7:0] n14_I_8_2; // @[Top.scala 139:21]
  wire [7:0] n14_I_9_0; // @[Top.scala 139:21]
  wire [7:0] n14_I_9_1; // @[Top.scala 139:21]
  wire [7:0] n14_I_9_2; // @[Top.scala 139:21]
  wire [7:0] n14_I_10_0; // @[Top.scala 139:21]
  wire [7:0] n14_I_10_1; // @[Top.scala 139:21]
  wire [7:0] n14_I_10_2; // @[Top.scala 139:21]
  wire [7:0] n14_I_11_0; // @[Top.scala 139:21]
  wire [7:0] n14_I_11_1; // @[Top.scala 139:21]
  wire [7:0] n14_I_11_2; // @[Top.scala 139:21]
  wire [7:0] n14_I_12_0; // @[Top.scala 139:21]
  wire [7:0] n14_I_12_1; // @[Top.scala 139:21]
  wire [7:0] n14_I_12_2; // @[Top.scala 139:21]
  wire [7:0] n14_I_13_0; // @[Top.scala 139:21]
  wire [7:0] n14_I_13_1; // @[Top.scala 139:21]
  wire [7:0] n14_I_13_2; // @[Top.scala 139:21]
  wire [7:0] n14_I_14_0; // @[Top.scala 139:21]
  wire [7:0] n14_I_14_1; // @[Top.scala 139:21]
  wire [7:0] n14_I_14_2; // @[Top.scala 139:21]
  wire [7:0] n14_I_15_0; // @[Top.scala 139:21]
  wire [7:0] n14_I_15_1; // @[Top.scala 139:21]
  wire [7:0] n14_I_15_2; // @[Top.scala 139:21]
  wire [7:0] n14_O_0_0_0; // @[Top.scala 139:21]
  wire [7:0] n14_O_0_0_1; // @[Top.scala 139:21]
  wire [7:0] n14_O_0_0_2; // @[Top.scala 139:21]
  wire [7:0] n14_O_1_0_0; // @[Top.scala 139:21]
  wire [7:0] n14_O_1_0_1; // @[Top.scala 139:21]
  wire [7:0] n14_O_1_0_2; // @[Top.scala 139:21]
  wire [7:0] n14_O_2_0_0; // @[Top.scala 139:21]
  wire [7:0] n14_O_2_0_1; // @[Top.scala 139:21]
  wire [7:0] n14_O_2_0_2; // @[Top.scala 139:21]
  wire [7:0] n14_O_3_0_0; // @[Top.scala 139:21]
  wire [7:0] n14_O_3_0_1; // @[Top.scala 139:21]
  wire [7:0] n14_O_3_0_2; // @[Top.scala 139:21]
  wire [7:0] n14_O_4_0_0; // @[Top.scala 139:21]
  wire [7:0] n14_O_4_0_1; // @[Top.scala 139:21]
  wire [7:0] n14_O_4_0_2; // @[Top.scala 139:21]
  wire [7:0] n14_O_5_0_0; // @[Top.scala 139:21]
  wire [7:0] n14_O_5_0_1; // @[Top.scala 139:21]
  wire [7:0] n14_O_5_0_2; // @[Top.scala 139:21]
  wire [7:0] n14_O_6_0_0; // @[Top.scala 139:21]
  wire [7:0] n14_O_6_0_1; // @[Top.scala 139:21]
  wire [7:0] n14_O_6_0_2; // @[Top.scala 139:21]
  wire [7:0] n14_O_7_0_0; // @[Top.scala 139:21]
  wire [7:0] n14_O_7_0_1; // @[Top.scala 139:21]
  wire [7:0] n14_O_7_0_2; // @[Top.scala 139:21]
  wire [7:0] n14_O_8_0_0; // @[Top.scala 139:21]
  wire [7:0] n14_O_8_0_1; // @[Top.scala 139:21]
  wire [7:0] n14_O_8_0_2; // @[Top.scala 139:21]
  wire [7:0] n14_O_9_0_0; // @[Top.scala 139:21]
  wire [7:0] n14_O_9_0_1; // @[Top.scala 139:21]
  wire [7:0] n14_O_9_0_2; // @[Top.scala 139:21]
  wire [7:0] n14_O_10_0_0; // @[Top.scala 139:21]
  wire [7:0] n14_O_10_0_1; // @[Top.scala 139:21]
  wire [7:0] n14_O_10_0_2; // @[Top.scala 139:21]
  wire [7:0] n14_O_11_0_0; // @[Top.scala 139:21]
  wire [7:0] n14_O_11_0_1; // @[Top.scala 139:21]
  wire [7:0] n14_O_11_0_2; // @[Top.scala 139:21]
  wire [7:0] n14_O_12_0_0; // @[Top.scala 139:21]
  wire [7:0] n14_O_12_0_1; // @[Top.scala 139:21]
  wire [7:0] n14_O_12_0_2; // @[Top.scala 139:21]
  wire [7:0] n14_O_13_0_0; // @[Top.scala 139:21]
  wire [7:0] n14_O_13_0_1; // @[Top.scala 139:21]
  wire [7:0] n14_O_13_0_2; // @[Top.scala 139:21]
  wire [7:0] n14_O_14_0_0; // @[Top.scala 139:21]
  wire [7:0] n14_O_14_0_1; // @[Top.scala 139:21]
  wire [7:0] n14_O_14_0_2; // @[Top.scala 139:21]
  wire [7:0] n14_O_15_0_0; // @[Top.scala 139:21]
  wire [7:0] n14_O_15_0_1; // @[Top.scala 139:21]
  wire [7:0] n14_O_15_0_2; // @[Top.scala 139:21]
  wire  n19_valid_up; // @[Top.scala 142:21]
  wire  n19_valid_down; // @[Top.scala 142:21]
  wire [7:0] n19_I_0_0_0; // @[Top.scala 142:21]
  wire [7:0] n19_I_0_0_1; // @[Top.scala 142:21]
  wire [7:0] n19_I_0_0_2; // @[Top.scala 142:21]
  wire [7:0] n19_I_1_0_0; // @[Top.scala 142:21]
  wire [7:0] n19_I_1_0_1; // @[Top.scala 142:21]
  wire [7:0] n19_I_1_0_2; // @[Top.scala 142:21]
  wire [7:0] n19_I_2_0_0; // @[Top.scala 142:21]
  wire [7:0] n19_I_2_0_1; // @[Top.scala 142:21]
  wire [7:0] n19_I_2_0_2; // @[Top.scala 142:21]
  wire [7:0] n19_I_3_0_0; // @[Top.scala 142:21]
  wire [7:0] n19_I_3_0_1; // @[Top.scala 142:21]
  wire [7:0] n19_I_3_0_2; // @[Top.scala 142:21]
  wire [7:0] n19_I_4_0_0; // @[Top.scala 142:21]
  wire [7:0] n19_I_4_0_1; // @[Top.scala 142:21]
  wire [7:0] n19_I_4_0_2; // @[Top.scala 142:21]
  wire [7:0] n19_I_5_0_0; // @[Top.scala 142:21]
  wire [7:0] n19_I_5_0_1; // @[Top.scala 142:21]
  wire [7:0] n19_I_5_0_2; // @[Top.scala 142:21]
  wire [7:0] n19_I_6_0_0; // @[Top.scala 142:21]
  wire [7:0] n19_I_6_0_1; // @[Top.scala 142:21]
  wire [7:0] n19_I_6_0_2; // @[Top.scala 142:21]
  wire [7:0] n19_I_7_0_0; // @[Top.scala 142:21]
  wire [7:0] n19_I_7_0_1; // @[Top.scala 142:21]
  wire [7:0] n19_I_7_0_2; // @[Top.scala 142:21]
  wire [7:0] n19_I_8_0_0; // @[Top.scala 142:21]
  wire [7:0] n19_I_8_0_1; // @[Top.scala 142:21]
  wire [7:0] n19_I_8_0_2; // @[Top.scala 142:21]
  wire [7:0] n19_I_9_0_0; // @[Top.scala 142:21]
  wire [7:0] n19_I_9_0_1; // @[Top.scala 142:21]
  wire [7:0] n19_I_9_0_2; // @[Top.scala 142:21]
  wire [7:0] n19_I_10_0_0; // @[Top.scala 142:21]
  wire [7:0] n19_I_10_0_1; // @[Top.scala 142:21]
  wire [7:0] n19_I_10_0_2; // @[Top.scala 142:21]
  wire [7:0] n19_I_11_0_0; // @[Top.scala 142:21]
  wire [7:0] n19_I_11_0_1; // @[Top.scala 142:21]
  wire [7:0] n19_I_11_0_2; // @[Top.scala 142:21]
  wire [7:0] n19_I_12_0_0; // @[Top.scala 142:21]
  wire [7:0] n19_I_12_0_1; // @[Top.scala 142:21]
  wire [7:0] n19_I_12_0_2; // @[Top.scala 142:21]
  wire [7:0] n19_I_13_0_0; // @[Top.scala 142:21]
  wire [7:0] n19_I_13_0_1; // @[Top.scala 142:21]
  wire [7:0] n19_I_13_0_2; // @[Top.scala 142:21]
  wire [7:0] n19_I_14_0_0; // @[Top.scala 142:21]
  wire [7:0] n19_I_14_0_1; // @[Top.scala 142:21]
  wire [7:0] n19_I_14_0_2; // @[Top.scala 142:21]
  wire [7:0] n19_I_15_0_0; // @[Top.scala 142:21]
  wire [7:0] n19_I_15_0_1; // @[Top.scala 142:21]
  wire [7:0] n19_I_15_0_2; // @[Top.scala 142:21]
  wire [7:0] n19_O_0_0; // @[Top.scala 142:21]
  wire [7:0] n19_O_0_1; // @[Top.scala 142:21]
  wire [7:0] n19_O_0_2; // @[Top.scala 142:21]
  wire [7:0] n19_O_1_0; // @[Top.scala 142:21]
  wire [7:0] n19_O_1_1; // @[Top.scala 142:21]
  wire [7:0] n19_O_1_2; // @[Top.scala 142:21]
  wire [7:0] n19_O_2_0; // @[Top.scala 142:21]
  wire [7:0] n19_O_2_1; // @[Top.scala 142:21]
  wire [7:0] n19_O_2_2; // @[Top.scala 142:21]
  wire [7:0] n19_O_3_0; // @[Top.scala 142:21]
  wire [7:0] n19_O_3_1; // @[Top.scala 142:21]
  wire [7:0] n19_O_3_2; // @[Top.scala 142:21]
  wire [7:0] n19_O_4_0; // @[Top.scala 142:21]
  wire [7:0] n19_O_4_1; // @[Top.scala 142:21]
  wire [7:0] n19_O_4_2; // @[Top.scala 142:21]
  wire [7:0] n19_O_5_0; // @[Top.scala 142:21]
  wire [7:0] n19_O_5_1; // @[Top.scala 142:21]
  wire [7:0] n19_O_5_2; // @[Top.scala 142:21]
  wire [7:0] n19_O_6_0; // @[Top.scala 142:21]
  wire [7:0] n19_O_6_1; // @[Top.scala 142:21]
  wire [7:0] n19_O_6_2; // @[Top.scala 142:21]
  wire [7:0] n19_O_7_0; // @[Top.scala 142:21]
  wire [7:0] n19_O_7_1; // @[Top.scala 142:21]
  wire [7:0] n19_O_7_2; // @[Top.scala 142:21]
  wire [7:0] n19_O_8_0; // @[Top.scala 142:21]
  wire [7:0] n19_O_8_1; // @[Top.scala 142:21]
  wire [7:0] n19_O_8_2; // @[Top.scala 142:21]
  wire [7:0] n19_O_9_0; // @[Top.scala 142:21]
  wire [7:0] n19_O_9_1; // @[Top.scala 142:21]
  wire [7:0] n19_O_9_2; // @[Top.scala 142:21]
  wire [7:0] n19_O_10_0; // @[Top.scala 142:21]
  wire [7:0] n19_O_10_1; // @[Top.scala 142:21]
  wire [7:0] n19_O_10_2; // @[Top.scala 142:21]
  wire [7:0] n19_O_11_0; // @[Top.scala 142:21]
  wire [7:0] n19_O_11_1; // @[Top.scala 142:21]
  wire [7:0] n19_O_11_2; // @[Top.scala 142:21]
  wire [7:0] n19_O_12_0; // @[Top.scala 142:21]
  wire [7:0] n19_O_12_1; // @[Top.scala 142:21]
  wire [7:0] n19_O_12_2; // @[Top.scala 142:21]
  wire [7:0] n19_O_13_0; // @[Top.scala 142:21]
  wire [7:0] n19_O_13_1; // @[Top.scala 142:21]
  wire [7:0] n19_O_13_2; // @[Top.scala 142:21]
  wire [7:0] n19_O_14_0; // @[Top.scala 142:21]
  wire [7:0] n19_O_14_1; // @[Top.scala 142:21]
  wire [7:0] n19_O_14_2; // @[Top.scala 142:21]
  wire [7:0] n19_O_15_0; // @[Top.scala 142:21]
  wire [7:0] n19_O_15_1; // @[Top.scala 142:21]
  wire [7:0] n19_O_15_2; // @[Top.scala 142:21]
  wire  n20_valid_up; // @[Top.scala 145:21]
  wire  n20_valid_down; // @[Top.scala 145:21]
  wire [7:0] n20_I_0; // @[Top.scala 145:21]
  wire [7:0] n20_I_1; // @[Top.scala 145:21]
  wire [7:0] n20_I_2; // @[Top.scala 145:21]
  wire [7:0] n20_I_3; // @[Top.scala 145:21]
  wire [7:0] n20_I_4; // @[Top.scala 145:21]
  wire [7:0] n20_I_5; // @[Top.scala 145:21]
  wire [7:0] n20_I_6; // @[Top.scala 145:21]
  wire [7:0] n20_I_7; // @[Top.scala 145:21]
  wire [7:0] n20_I_8; // @[Top.scala 145:21]
  wire [7:0] n20_I_9; // @[Top.scala 145:21]
  wire [7:0] n20_I_10; // @[Top.scala 145:21]
  wire [7:0] n20_I_11; // @[Top.scala 145:21]
  wire [7:0] n20_I_12; // @[Top.scala 145:21]
  wire [7:0] n20_I_13; // @[Top.scala 145:21]
  wire [7:0] n20_I_14; // @[Top.scala 145:21]
  wire [7:0] n20_I_15; // @[Top.scala 145:21]
  wire [7:0] n20_O_0; // @[Top.scala 145:21]
  wire [7:0] n20_O_1; // @[Top.scala 145:21]
  wire [7:0] n20_O_2; // @[Top.scala 145:21]
  wire [7:0] n20_O_3; // @[Top.scala 145:21]
  wire [7:0] n20_O_4; // @[Top.scala 145:21]
  wire [7:0] n20_O_5; // @[Top.scala 145:21]
  wire [7:0] n20_O_6; // @[Top.scala 145:21]
  wire [7:0] n20_O_7; // @[Top.scala 145:21]
  wire [7:0] n20_O_8; // @[Top.scala 145:21]
  wire [7:0] n20_O_9; // @[Top.scala 145:21]
  wire [7:0] n20_O_10; // @[Top.scala 145:21]
  wire [7:0] n20_O_11; // @[Top.scala 145:21]
  wire [7:0] n20_O_12; // @[Top.scala 145:21]
  wire [7:0] n20_O_13; // @[Top.scala 145:21]
  wire [7:0] n20_O_14; // @[Top.scala 145:21]
  wire [7:0] n20_O_15; // @[Top.scala 145:21]
  wire  n21_valid_up; // @[Top.scala 148:21]
  wire  n21_valid_down; // @[Top.scala 148:21]
  wire [7:0] n21_I_0; // @[Top.scala 148:21]
  wire [7:0] n21_I_1; // @[Top.scala 148:21]
  wire [7:0] n21_I_2; // @[Top.scala 148:21]
  wire [7:0] n21_I_3; // @[Top.scala 148:21]
  wire [7:0] n21_I_4; // @[Top.scala 148:21]
  wire [7:0] n21_I_5; // @[Top.scala 148:21]
  wire [7:0] n21_I_6; // @[Top.scala 148:21]
  wire [7:0] n21_I_7; // @[Top.scala 148:21]
  wire [7:0] n21_I_8; // @[Top.scala 148:21]
  wire [7:0] n21_I_9; // @[Top.scala 148:21]
  wire [7:0] n21_I_10; // @[Top.scala 148:21]
  wire [7:0] n21_I_11; // @[Top.scala 148:21]
  wire [7:0] n21_I_12; // @[Top.scala 148:21]
  wire [7:0] n21_I_13; // @[Top.scala 148:21]
  wire [7:0] n21_I_14; // @[Top.scala 148:21]
  wire [7:0] n21_I_15; // @[Top.scala 148:21]
  wire [7:0] n21_O_0; // @[Top.scala 148:21]
  wire [7:0] n21_O_1; // @[Top.scala 148:21]
  wire [7:0] n21_O_2; // @[Top.scala 148:21]
  wire [7:0] n21_O_3; // @[Top.scala 148:21]
  wire [7:0] n21_O_4; // @[Top.scala 148:21]
  wire [7:0] n21_O_5; // @[Top.scala 148:21]
  wire [7:0] n21_O_6; // @[Top.scala 148:21]
  wire [7:0] n21_O_7; // @[Top.scala 148:21]
  wire [7:0] n21_O_8; // @[Top.scala 148:21]
  wire [7:0] n21_O_9; // @[Top.scala 148:21]
  wire [7:0] n21_O_10; // @[Top.scala 148:21]
  wire [7:0] n21_O_11; // @[Top.scala 148:21]
  wire [7:0] n21_O_12; // @[Top.scala 148:21]
  wire [7:0] n21_O_13; // @[Top.scala 148:21]
  wire [7:0] n21_O_14; // @[Top.scala 148:21]
  wire [7:0] n21_O_15; // @[Top.scala 148:21]
  wire  n22_valid_up; // @[Top.scala 151:21]
  wire  n22_valid_down; // @[Top.scala 151:21]
  wire [7:0] n22_I0_0; // @[Top.scala 151:21]
  wire [7:0] n22_I0_1; // @[Top.scala 151:21]
  wire [7:0] n22_I0_2; // @[Top.scala 151:21]
  wire [7:0] n22_I0_3; // @[Top.scala 151:21]
  wire [7:0] n22_I0_4; // @[Top.scala 151:21]
  wire [7:0] n22_I0_5; // @[Top.scala 151:21]
  wire [7:0] n22_I0_6; // @[Top.scala 151:21]
  wire [7:0] n22_I0_7; // @[Top.scala 151:21]
  wire [7:0] n22_I0_8; // @[Top.scala 151:21]
  wire [7:0] n22_I0_9; // @[Top.scala 151:21]
  wire [7:0] n22_I0_10; // @[Top.scala 151:21]
  wire [7:0] n22_I0_11; // @[Top.scala 151:21]
  wire [7:0] n22_I0_12; // @[Top.scala 151:21]
  wire [7:0] n22_I0_13; // @[Top.scala 151:21]
  wire [7:0] n22_I0_14; // @[Top.scala 151:21]
  wire [7:0] n22_I0_15; // @[Top.scala 151:21]
  wire [7:0] n22_I1_0; // @[Top.scala 151:21]
  wire [7:0] n22_I1_1; // @[Top.scala 151:21]
  wire [7:0] n22_I1_2; // @[Top.scala 151:21]
  wire [7:0] n22_I1_3; // @[Top.scala 151:21]
  wire [7:0] n22_I1_4; // @[Top.scala 151:21]
  wire [7:0] n22_I1_5; // @[Top.scala 151:21]
  wire [7:0] n22_I1_6; // @[Top.scala 151:21]
  wire [7:0] n22_I1_7; // @[Top.scala 151:21]
  wire [7:0] n22_I1_8; // @[Top.scala 151:21]
  wire [7:0] n22_I1_9; // @[Top.scala 151:21]
  wire [7:0] n22_I1_10; // @[Top.scala 151:21]
  wire [7:0] n22_I1_11; // @[Top.scala 151:21]
  wire [7:0] n22_I1_12; // @[Top.scala 151:21]
  wire [7:0] n22_I1_13; // @[Top.scala 151:21]
  wire [7:0] n22_I1_14; // @[Top.scala 151:21]
  wire [7:0] n22_I1_15; // @[Top.scala 151:21]
  wire [7:0] n22_O_0_0; // @[Top.scala 151:21]
  wire [7:0] n22_O_0_1; // @[Top.scala 151:21]
  wire [7:0] n22_O_1_0; // @[Top.scala 151:21]
  wire [7:0] n22_O_1_1; // @[Top.scala 151:21]
  wire [7:0] n22_O_2_0; // @[Top.scala 151:21]
  wire [7:0] n22_O_2_1; // @[Top.scala 151:21]
  wire [7:0] n22_O_3_0; // @[Top.scala 151:21]
  wire [7:0] n22_O_3_1; // @[Top.scala 151:21]
  wire [7:0] n22_O_4_0; // @[Top.scala 151:21]
  wire [7:0] n22_O_4_1; // @[Top.scala 151:21]
  wire [7:0] n22_O_5_0; // @[Top.scala 151:21]
  wire [7:0] n22_O_5_1; // @[Top.scala 151:21]
  wire [7:0] n22_O_6_0; // @[Top.scala 151:21]
  wire [7:0] n22_O_6_1; // @[Top.scala 151:21]
  wire [7:0] n22_O_7_0; // @[Top.scala 151:21]
  wire [7:0] n22_O_7_1; // @[Top.scala 151:21]
  wire [7:0] n22_O_8_0; // @[Top.scala 151:21]
  wire [7:0] n22_O_8_1; // @[Top.scala 151:21]
  wire [7:0] n22_O_9_0; // @[Top.scala 151:21]
  wire [7:0] n22_O_9_1; // @[Top.scala 151:21]
  wire [7:0] n22_O_10_0; // @[Top.scala 151:21]
  wire [7:0] n22_O_10_1; // @[Top.scala 151:21]
  wire [7:0] n22_O_11_0; // @[Top.scala 151:21]
  wire [7:0] n22_O_11_1; // @[Top.scala 151:21]
  wire [7:0] n22_O_12_0; // @[Top.scala 151:21]
  wire [7:0] n22_O_12_1; // @[Top.scala 151:21]
  wire [7:0] n22_O_13_0; // @[Top.scala 151:21]
  wire [7:0] n22_O_13_1; // @[Top.scala 151:21]
  wire [7:0] n22_O_14_0; // @[Top.scala 151:21]
  wire [7:0] n22_O_14_1; // @[Top.scala 151:21]
  wire [7:0] n22_O_15_0; // @[Top.scala 151:21]
  wire [7:0] n22_O_15_1; // @[Top.scala 151:21]
  wire  n26_valid_up; // @[Top.scala 155:21]
  wire  n26_valid_down; // @[Top.scala 155:21]
  wire [7:0] n26_I0_0_0; // @[Top.scala 155:21]
  wire [7:0] n26_I0_0_1; // @[Top.scala 155:21]
  wire [7:0] n26_I0_1_0; // @[Top.scala 155:21]
  wire [7:0] n26_I0_1_1; // @[Top.scala 155:21]
  wire [7:0] n26_I0_2_0; // @[Top.scala 155:21]
  wire [7:0] n26_I0_2_1; // @[Top.scala 155:21]
  wire [7:0] n26_I0_3_0; // @[Top.scala 155:21]
  wire [7:0] n26_I0_3_1; // @[Top.scala 155:21]
  wire [7:0] n26_I0_4_0; // @[Top.scala 155:21]
  wire [7:0] n26_I0_4_1; // @[Top.scala 155:21]
  wire [7:0] n26_I0_5_0; // @[Top.scala 155:21]
  wire [7:0] n26_I0_5_1; // @[Top.scala 155:21]
  wire [7:0] n26_I0_6_0; // @[Top.scala 155:21]
  wire [7:0] n26_I0_6_1; // @[Top.scala 155:21]
  wire [7:0] n26_I0_7_0; // @[Top.scala 155:21]
  wire [7:0] n26_I0_7_1; // @[Top.scala 155:21]
  wire [7:0] n26_I0_8_0; // @[Top.scala 155:21]
  wire [7:0] n26_I0_8_1; // @[Top.scala 155:21]
  wire [7:0] n26_I0_9_0; // @[Top.scala 155:21]
  wire [7:0] n26_I0_9_1; // @[Top.scala 155:21]
  wire [7:0] n26_I0_10_0; // @[Top.scala 155:21]
  wire [7:0] n26_I0_10_1; // @[Top.scala 155:21]
  wire [7:0] n26_I0_11_0; // @[Top.scala 155:21]
  wire [7:0] n26_I0_11_1; // @[Top.scala 155:21]
  wire [7:0] n26_I0_12_0; // @[Top.scala 155:21]
  wire [7:0] n26_I0_12_1; // @[Top.scala 155:21]
  wire [7:0] n26_I0_13_0; // @[Top.scala 155:21]
  wire [7:0] n26_I0_13_1; // @[Top.scala 155:21]
  wire [7:0] n26_I0_14_0; // @[Top.scala 155:21]
  wire [7:0] n26_I0_14_1; // @[Top.scala 155:21]
  wire [7:0] n26_I0_15_0; // @[Top.scala 155:21]
  wire [7:0] n26_I0_15_1; // @[Top.scala 155:21]
  wire [7:0] n26_I1_0; // @[Top.scala 155:21]
  wire [7:0] n26_I1_1; // @[Top.scala 155:21]
  wire [7:0] n26_I1_2; // @[Top.scala 155:21]
  wire [7:0] n26_I1_3; // @[Top.scala 155:21]
  wire [7:0] n26_I1_4; // @[Top.scala 155:21]
  wire [7:0] n26_I1_5; // @[Top.scala 155:21]
  wire [7:0] n26_I1_6; // @[Top.scala 155:21]
  wire [7:0] n26_I1_7; // @[Top.scala 155:21]
  wire [7:0] n26_I1_8; // @[Top.scala 155:21]
  wire [7:0] n26_I1_9; // @[Top.scala 155:21]
  wire [7:0] n26_I1_10; // @[Top.scala 155:21]
  wire [7:0] n26_I1_11; // @[Top.scala 155:21]
  wire [7:0] n26_I1_12; // @[Top.scala 155:21]
  wire [7:0] n26_I1_13; // @[Top.scala 155:21]
  wire [7:0] n26_I1_14; // @[Top.scala 155:21]
  wire [7:0] n26_I1_15; // @[Top.scala 155:21]
  wire [7:0] n26_O_0_0; // @[Top.scala 155:21]
  wire [7:0] n26_O_0_1; // @[Top.scala 155:21]
  wire [7:0] n26_O_0_2; // @[Top.scala 155:21]
  wire [7:0] n26_O_1_0; // @[Top.scala 155:21]
  wire [7:0] n26_O_1_1; // @[Top.scala 155:21]
  wire [7:0] n26_O_1_2; // @[Top.scala 155:21]
  wire [7:0] n26_O_2_0; // @[Top.scala 155:21]
  wire [7:0] n26_O_2_1; // @[Top.scala 155:21]
  wire [7:0] n26_O_2_2; // @[Top.scala 155:21]
  wire [7:0] n26_O_3_0; // @[Top.scala 155:21]
  wire [7:0] n26_O_3_1; // @[Top.scala 155:21]
  wire [7:0] n26_O_3_2; // @[Top.scala 155:21]
  wire [7:0] n26_O_4_0; // @[Top.scala 155:21]
  wire [7:0] n26_O_4_1; // @[Top.scala 155:21]
  wire [7:0] n26_O_4_2; // @[Top.scala 155:21]
  wire [7:0] n26_O_5_0; // @[Top.scala 155:21]
  wire [7:0] n26_O_5_1; // @[Top.scala 155:21]
  wire [7:0] n26_O_5_2; // @[Top.scala 155:21]
  wire [7:0] n26_O_6_0; // @[Top.scala 155:21]
  wire [7:0] n26_O_6_1; // @[Top.scala 155:21]
  wire [7:0] n26_O_6_2; // @[Top.scala 155:21]
  wire [7:0] n26_O_7_0; // @[Top.scala 155:21]
  wire [7:0] n26_O_7_1; // @[Top.scala 155:21]
  wire [7:0] n26_O_7_2; // @[Top.scala 155:21]
  wire [7:0] n26_O_8_0; // @[Top.scala 155:21]
  wire [7:0] n26_O_8_1; // @[Top.scala 155:21]
  wire [7:0] n26_O_8_2; // @[Top.scala 155:21]
  wire [7:0] n26_O_9_0; // @[Top.scala 155:21]
  wire [7:0] n26_O_9_1; // @[Top.scala 155:21]
  wire [7:0] n26_O_9_2; // @[Top.scala 155:21]
  wire [7:0] n26_O_10_0; // @[Top.scala 155:21]
  wire [7:0] n26_O_10_1; // @[Top.scala 155:21]
  wire [7:0] n26_O_10_2; // @[Top.scala 155:21]
  wire [7:0] n26_O_11_0; // @[Top.scala 155:21]
  wire [7:0] n26_O_11_1; // @[Top.scala 155:21]
  wire [7:0] n26_O_11_2; // @[Top.scala 155:21]
  wire [7:0] n26_O_12_0; // @[Top.scala 155:21]
  wire [7:0] n26_O_12_1; // @[Top.scala 155:21]
  wire [7:0] n26_O_12_2; // @[Top.scala 155:21]
  wire [7:0] n26_O_13_0; // @[Top.scala 155:21]
  wire [7:0] n26_O_13_1; // @[Top.scala 155:21]
  wire [7:0] n26_O_13_2; // @[Top.scala 155:21]
  wire [7:0] n26_O_14_0; // @[Top.scala 155:21]
  wire [7:0] n26_O_14_1; // @[Top.scala 155:21]
  wire [7:0] n26_O_14_2; // @[Top.scala 155:21]
  wire [7:0] n26_O_15_0; // @[Top.scala 155:21]
  wire [7:0] n26_O_15_1; // @[Top.scala 155:21]
  wire [7:0] n26_O_15_2; // @[Top.scala 155:21]
  wire  n30_valid_up; // @[Top.scala 159:21]
  wire  n30_valid_down; // @[Top.scala 159:21]
  wire [7:0] n30_I_0_0; // @[Top.scala 159:21]
  wire [7:0] n30_I_0_1; // @[Top.scala 159:21]
  wire [7:0] n30_I_0_2; // @[Top.scala 159:21]
  wire [7:0] n30_I_1_0; // @[Top.scala 159:21]
  wire [7:0] n30_I_1_1; // @[Top.scala 159:21]
  wire [7:0] n30_I_1_2; // @[Top.scala 159:21]
  wire [7:0] n30_I_2_0; // @[Top.scala 159:21]
  wire [7:0] n30_I_2_1; // @[Top.scala 159:21]
  wire [7:0] n30_I_2_2; // @[Top.scala 159:21]
  wire [7:0] n30_I_3_0; // @[Top.scala 159:21]
  wire [7:0] n30_I_3_1; // @[Top.scala 159:21]
  wire [7:0] n30_I_3_2; // @[Top.scala 159:21]
  wire [7:0] n30_I_4_0; // @[Top.scala 159:21]
  wire [7:0] n30_I_4_1; // @[Top.scala 159:21]
  wire [7:0] n30_I_4_2; // @[Top.scala 159:21]
  wire [7:0] n30_I_5_0; // @[Top.scala 159:21]
  wire [7:0] n30_I_5_1; // @[Top.scala 159:21]
  wire [7:0] n30_I_5_2; // @[Top.scala 159:21]
  wire [7:0] n30_I_6_0; // @[Top.scala 159:21]
  wire [7:0] n30_I_6_1; // @[Top.scala 159:21]
  wire [7:0] n30_I_6_2; // @[Top.scala 159:21]
  wire [7:0] n30_I_7_0; // @[Top.scala 159:21]
  wire [7:0] n30_I_7_1; // @[Top.scala 159:21]
  wire [7:0] n30_I_7_2; // @[Top.scala 159:21]
  wire [7:0] n30_I_8_0; // @[Top.scala 159:21]
  wire [7:0] n30_I_8_1; // @[Top.scala 159:21]
  wire [7:0] n30_I_8_2; // @[Top.scala 159:21]
  wire [7:0] n30_I_9_0; // @[Top.scala 159:21]
  wire [7:0] n30_I_9_1; // @[Top.scala 159:21]
  wire [7:0] n30_I_9_2; // @[Top.scala 159:21]
  wire [7:0] n30_I_10_0; // @[Top.scala 159:21]
  wire [7:0] n30_I_10_1; // @[Top.scala 159:21]
  wire [7:0] n30_I_10_2; // @[Top.scala 159:21]
  wire [7:0] n30_I_11_0; // @[Top.scala 159:21]
  wire [7:0] n30_I_11_1; // @[Top.scala 159:21]
  wire [7:0] n30_I_11_2; // @[Top.scala 159:21]
  wire [7:0] n30_I_12_0; // @[Top.scala 159:21]
  wire [7:0] n30_I_12_1; // @[Top.scala 159:21]
  wire [7:0] n30_I_12_2; // @[Top.scala 159:21]
  wire [7:0] n30_I_13_0; // @[Top.scala 159:21]
  wire [7:0] n30_I_13_1; // @[Top.scala 159:21]
  wire [7:0] n30_I_13_2; // @[Top.scala 159:21]
  wire [7:0] n30_I_14_0; // @[Top.scala 159:21]
  wire [7:0] n30_I_14_1; // @[Top.scala 159:21]
  wire [7:0] n30_I_14_2; // @[Top.scala 159:21]
  wire [7:0] n30_I_15_0; // @[Top.scala 159:21]
  wire [7:0] n30_I_15_1; // @[Top.scala 159:21]
  wire [7:0] n30_I_15_2; // @[Top.scala 159:21]
  wire [7:0] n30_O_0_0_0; // @[Top.scala 159:21]
  wire [7:0] n30_O_0_0_1; // @[Top.scala 159:21]
  wire [7:0] n30_O_0_0_2; // @[Top.scala 159:21]
  wire [7:0] n30_O_1_0_0; // @[Top.scala 159:21]
  wire [7:0] n30_O_1_0_1; // @[Top.scala 159:21]
  wire [7:0] n30_O_1_0_2; // @[Top.scala 159:21]
  wire [7:0] n30_O_2_0_0; // @[Top.scala 159:21]
  wire [7:0] n30_O_2_0_1; // @[Top.scala 159:21]
  wire [7:0] n30_O_2_0_2; // @[Top.scala 159:21]
  wire [7:0] n30_O_3_0_0; // @[Top.scala 159:21]
  wire [7:0] n30_O_3_0_1; // @[Top.scala 159:21]
  wire [7:0] n30_O_3_0_2; // @[Top.scala 159:21]
  wire [7:0] n30_O_4_0_0; // @[Top.scala 159:21]
  wire [7:0] n30_O_4_0_1; // @[Top.scala 159:21]
  wire [7:0] n30_O_4_0_2; // @[Top.scala 159:21]
  wire [7:0] n30_O_5_0_0; // @[Top.scala 159:21]
  wire [7:0] n30_O_5_0_1; // @[Top.scala 159:21]
  wire [7:0] n30_O_5_0_2; // @[Top.scala 159:21]
  wire [7:0] n30_O_6_0_0; // @[Top.scala 159:21]
  wire [7:0] n30_O_6_0_1; // @[Top.scala 159:21]
  wire [7:0] n30_O_6_0_2; // @[Top.scala 159:21]
  wire [7:0] n30_O_7_0_0; // @[Top.scala 159:21]
  wire [7:0] n30_O_7_0_1; // @[Top.scala 159:21]
  wire [7:0] n30_O_7_0_2; // @[Top.scala 159:21]
  wire [7:0] n30_O_8_0_0; // @[Top.scala 159:21]
  wire [7:0] n30_O_8_0_1; // @[Top.scala 159:21]
  wire [7:0] n30_O_8_0_2; // @[Top.scala 159:21]
  wire [7:0] n30_O_9_0_0; // @[Top.scala 159:21]
  wire [7:0] n30_O_9_0_1; // @[Top.scala 159:21]
  wire [7:0] n30_O_9_0_2; // @[Top.scala 159:21]
  wire [7:0] n30_O_10_0_0; // @[Top.scala 159:21]
  wire [7:0] n30_O_10_0_1; // @[Top.scala 159:21]
  wire [7:0] n30_O_10_0_2; // @[Top.scala 159:21]
  wire [7:0] n30_O_11_0_0; // @[Top.scala 159:21]
  wire [7:0] n30_O_11_0_1; // @[Top.scala 159:21]
  wire [7:0] n30_O_11_0_2; // @[Top.scala 159:21]
  wire [7:0] n30_O_12_0_0; // @[Top.scala 159:21]
  wire [7:0] n30_O_12_0_1; // @[Top.scala 159:21]
  wire [7:0] n30_O_12_0_2; // @[Top.scala 159:21]
  wire [7:0] n30_O_13_0_0; // @[Top.scala 159:21]
  wire [7:0] n30_O_13_0_1; // @[Top.scala 159:21]
  wire [7:0] n30_O_13_0_2; // @[Top.scala 159:21]
  wire [7:0] n30_O_14_0_0; // @[Top.scala 159:21]
  wire [7:0] n30_O_14_0_1; // @[Top.scala 159:21]
  wire [7:0] n30_O_14_0_2; // @[Top.scala 159:21]
  wire [7:0] n30_O_15_0_0; // @[Top.scala 159:21]
  wire [7:0] n30_O_15_0_1; // @[Top.scala 159:21]
  wire [7:0] n30_O_15_0_2; // @[Top.scala 159:21]
  wire  n35_valid_up; // @[Top.scala 162:21]
  wire  n35_valid_down; // @[Top.scala 162:21]
  wire [7:0] n35_I_0_0_0; // @[Top.scala 162:21]
  wire [7:0] n35_I_0_0_1; // @[Top.scala 162:21]
  wire [7:0] n35_I_0_0_2; // @[Top.scala 162:21]
  wire [7:0] n35_I_1_0_0; // @[Top.scala 162:21]
  wire [7:0] n35_I_1_0_1; // @[Top.scala 162:21]
  wire [7:0] n35_I_1_0_2; // @[Top.scala 162:21]
  wire [7:0] n35_I_2_0_0; // @[Top.scala 162:21]
  wire [7:0] n35_I_2_0_1; // @[Top.scala 162:21]
  wire [7:0] n35_I_2_0_2; // @[Top.scala 162:21]
  wire [7:0] n35_I_3_0_0; // @[Top.scala 162:21]
  wire [7:0] n35_I_3_0_1; // @[Top.scala 162:21]
  wire [7:0] n35_I_3_0_2; // @[Top.scala 162:21]
  wire [7:0] n35_I_4_0_0; // @[Top.scala 162:21]
  wire [7:0] n35_I_4_0_1; // @[Top.scala 162:21]
  wire [7:0] n35_I_4_0_2; // @[Top.scala 162:21]
  wire [7:0] n35_I_5_0_0; // @[Top.scala 162:21]
  wire [7:0] n35_I_5_0_1; // @[Top.scala 162:21]
  wire [7:0] n35_I_5_0_2; // @[Top.scala 162:21]
  wire [7:0] n35_I_6_0_0; // @[Top.scala 162:21]
  wire [7:0] n35_I_6_0_1; // @[Top.scala 162:21]
  wire [7:0] n35_I_6_0_2; // @[Top.scala 162:21]
  wire [7:0] n35_I_7_0_0; // @[Top.scala 162:21]
  wire [7:0] n35_I_7_0_1; // @[Top.scala 162:21]
  wire [7:0] n35_I_7_0_2; // @[Top.scala 162:21]
  wire [7:0] n35_I_8_0_0; // @[Top.scala 162:21]
  wire [7:0] n35_I_8_0_1; // @[Top.scala 162:21]
  wire [7:0] n35_I_8_0_2; // @[Top.scala 162:21]
  wire [7:0] n35_I_9_0_0; // @[Top.scala 162:21]
  wire [7:0] n35_I_9_0_1; // @[Top.scala 162:21]
  wire [7:0] n35_I_9_0_2; // @[Top.scala 162:21]
  wire [7:0] n35_I_10_0_0; // @[Top.scala 162:21]
  wire [7:0] n35_I_10_0_1; // @[Top.scala 162:21]
  wire [7:0] n35_I_10_0_2; // @[Top.scala 162:21]
  wire [7:0] n35_I_11_0_0; // @[Top.scala 162:21]
  wire [7:0] n35_I_11_0_1; // @[Top.scala 162:21]
  wire [7:0] n35_I_11_0_2; // @[Top.scala 162:21]
  wire [7:0] n35_I_12_0_0; // @[Top.scala 162:21]
  wire [7:0] n35_I_12_0_1; // @[Top.scala 162:21]
  wire [7:0] n35_I_12_0_2; // @[Top.scala 162:21]
  wire [7:0] n35_I_13_0_0; // @[Top.scala 162:21]
  wire [7:0] n35_I_13_0_1; // @[Top.scala 162:21]
  wire [7:0] n35_I_13_0_2; // @[Top.scala 162:21]
  wire [7:0] n35_I_14_0_0; // @[Top.scala 162:21]
  wire [7:0] n35_I_14_0_1; // @[Top.scala 162:21]
  wire [7:0] n35_I_14_0_2; // @[Top.scala 162:21]
  wire [7:0] n35_I_15_0_0; // @[Top.scala 162:21]
  wire [7:0] n35_I_15_0_1; // @[Top.scala 162:21]
  wire [7:0] n35_I_15_0_2; // @[Top.scala 162:21]
  wire [7:0] n35_O_0_0; // @[Top.scala 162:21]
  wire [7:0] n35_O_0_1; // @[Top.scala 162:21]
  wire [7:0] n35_O_0_2; // @[Top.scala 162:21]
  wire [7:0] n35_O_1_0; // @[Top.scala 162:21]
  wire [7:0] n35_O_1_1; // @[Top.scala 162:21]
  wire [7:0] n35_O_1_2; // @[Top.scala 162:21]
  wire [7:0] n35_O_2_0; // @[Top.scala 162:21]
  wire [7:0] n35_O_2_1; // @[Top.scala 162:21]
  wire [7:0] n35_O_2_2; // @[Top.scala 162:21]
  wire [7:0] n35_O_3_0; // @[Top.scala 162:21]
  wire [7:0] n35_O_3_1; // @[Top.scala 162:21]
  wire [7:0] n35_O_3_2; // @[Top.scala 162:21]
  wire [7:0] n35_O_4_0; // @[Top.scala 162:21]
  wire [7:0] n35_O_4_1; // @[Top.scala 162:21]
  wire [7:0] n35_O_4_2; // @[Top.scala 162:21]
  wire [7:0] n35_O_5_0; // @[Top.scala 162:21]
  wire [7:0] n35_O_5_1; // @[Top.scala 162:21]
  wire [7:0] n35_O_5_2; // @[Top.scala 162:21]
  wire [7:0] n35_O_6_0; // @[Top.scala 162:21]
  wire [7:0] n35_O_6_1; // @[Top.scala 162:21]
  wire [7:0] n35_O_6_2; // @[Top.scala 162:21]
  wire [7:0] n35_O_7_0; // @[Top.scala 162:21]
  wire [7:0] n35_O_7_1; // @[Top.scala 162:21]
  wire [7:0] n35_O_7_2; // @[Top.scala 162:21]
  wire [7:0] n35_O_8_0; // @[Top.scala 162:21]
  wire [7:0] n35_O_8_1; // @[Top.scala 162:21]
  wire [7:0] n35_O_8_2; // @[Top.scala 162:21]
  wire [7:0] n35_O_9_0; // @[Top.scala 162:21]
  wire [7:0] n35_O_9_1; // @[Top.scala 162:21]
  wire [7:0] n35_O_9_2; // @[Top.scala 162:21]
  wire [7:0] n35_O_10_0; // @[Top.scala 162:21]
  wire [7:0] n35_O_10_1; // @[Top.scala 162:21]
  wire [7:0] n35_O_10_2; // @[Top.scala 162:21]
  wire [7:0] n35_O_11_0; // @[Top.scala 162:21]
  wire [7:0] n35_O_11_1; // @[Top.scala 162:21]
  wire [7:0] n35_O_11_2; // @[Top.scala 162:21]
  wire [7:0] n35_O_12_0; // @[Top.scala 162:21]
  wire [7:0] n35_O_12_1; // @[Top.scala 162:21]
  wire [7:0] n35_O_12_2; // @[Top.scala 162:21]
  wire [7:0] n35_O_13_0; // @[Top.scala 162:21]
  wire [7:0] n35_O_13_1; // @[Top.scala 162:21]
  wire [7:0] n35_O_13_2; // @[Top.scala 162:21]
  wire [7:0] n35_O_14_0; // @[Top.scala 162:21]
  wire [7:0] n35_O_14_1; // @[Top.scala 162:21]
  wire [7:0] n35_O_14_2; // @[Top.scala 162:21]
  wire [7:0] n35_O_15_0; // @[Top.scala 162:21]
  wire [7:0] n35_O_15_1; // @[Top.scala 162:21]
  wire [7:0] n35_O_15_2; // @[Top.scala 162:21]
  wire  n36_valid_up; // @[Top.scala 165:21]
  wire  n36_valid_down; // @[Top.scala 165:21]
  wire [7:0] n36_I0_0_0; // @[Top.scala 165:21]
  wire [7:0] n36_I0_0_1; // @[Top.scala 165:21]
  wire [7:0] n36_I0_0_2; // @[Top.scala 165:21]
  wire [7:0] n36_I0_1_0; // @[Top.scala 165:21]
  wire [7:0] n36_I0_1_1; // @[Top.scala 165:21]
  wire [7:0] n36_I0_1_2; // @[Top.scala 165:21]
  wire [7:0] n36_I0_2_0; // @[Top.scala 165:21]
  wire [7:0] n36_I0_2_1; // @[Top.scala 165:21]
  wire [7:0] n36_I0_2_2; // @[Top.scala 165:21]
  wire [7:0] n36_I0_3_0; // @[Top.scala 165:21]
  wire [7:0] n36_I0_3_1; // @[Top.scala 165:21]
  wire [7:0] n36_I0_3_2; // @[Top.scala 165:21]
  wire [7:0] n36_I0_4_0; // @[Top.scala 165:21]
  wire [7:0] n36_I0_4_1; // @[Top.scala 165:21]
  wire [7:0] n36_I0_4_2; // @[Top.scala 165:21]
  wire [7:0] n36_I0_5_0; // @[Top.scala 165:21]
  wire [7:0] n36_I0_5_1; // @[Top.scala 165:21]
  wire [7:0] n36_I0_5_2; // @[Top.scala 165:21]
  wire [7:0] n36_I0_6_0; // @[Top.scala 165:21]
  wire [7:0] n36_I0_6_1; // @[Top.scala 165:21]
  wire [7:0] n36_I0_6_2; // @[Top.scala 165:21]
  wire [7:0] n36_I0_7_0; // @[Top.scala 165:21]
  wire [7:0] n36_I0_7_1; // @[Top.scala 165:21]
  wire [7:0] n36_I0_7_2; // @[Top.scala 165:21]
  wire [7:0] n36_I0_8_0; // @[Top.scala 165:21]
  wire [7:0] n36_I0_8_1; // @[Top.scala 165:21]
  wire [7:0] n36_I0_8_2; // @[Top.scala 165:21]
  wire [7:0] n36_I0_9_0; // @[Top.scala 165:21]
  wire [7:0] n36_I0_9_1; // @[Top.scala 165:21]
  wire [7:0] n36_I0_9_2; // @[Top.scala 165:21]
  wire [7:0] n36_I0_10_0; // @[Top.scala 165:21]
  wire [7:0] n36_I0_10_1; // @[Top.scala 165:21]
  wire [7:0] n36_I0_10_2; // @[Top.scala 165:21]
  wire [7:0] n36_I0_11_0; // @[Top.scala 165:21]
  wire [7:0] n36_I0_11_1; // @[Top.scala 165:21]
  wire [7:0] n36_I0_11_2; // @[Top.scala 165:21]
  wire [7:0] n36_I0_12_0; // @[Top.scala 165:21]
  wire [7:0] n36_I0_12_1; // @[Top.scala 165:21]
  wire [7:0] n36_I0_12_2; // @[Top.scala 165:21]
  wire [7:0] n36_I0_13_0; // @[Top.scala 165:21]
  wire [7:0] n36_I0_13_1; // @[Top.scala 165:21]
  wire [7:0] n36_I0_13_2; // @[Top.scala 165:21]
  wire [7:0] n36_I0_14_0; // @[Top.scala 165:21]
  wire [7:0] n36_I0_14_1; // @[Top.scala 165:21]
  wire [7:0] n36_I0_14_2; // @[Top.scala 165:21]
  wire [7:0] n36_I0_15_0; // @[Top.scala 165:21]
  wire [7:0] n36_I0_15_1; // @[Top.scala 165:21]
  wire [7:0] n36_I0_15_2; // @[Top.scala 165:21]
  wire [7:0] n36_I1_0_0; // @[Top.scala 165:21]
  wire [7:0] n36_I1_0_1; // @[Top.scala 165:21]
  wire [7:0] n36_I1_0_2; // @[Top.scala 165:21]
  wire [7:0] n36_I1_1_0; // @[Top.scala 165:21]
  wire [7:0] n36_I1_1_1; // @[Top.scala 165:21]
  wire [7:0] n36_I1_1_2; // @[Top.scala 165:21]
  wire [7:0] n36_I1_2_0; // @[Top.scala 165:21]
  wire [7:0] n36_I1_2_1; // @[Top.scala 165:21]
  wire [7:0] n36_I1_2_2; // @[Top.scala 165:21]
  wire [7:0] n36_I1_3_0; // @[Top.scala 165:21]
  wire [7:0] n36_I1_3_1; // @[Top.scala 165:21]
  wire [7:0] n36_I1_3_2; // @[Top.scala 165:21]
  wire [7:0] n36_I1_4_0; // @[Top.scala 165:21]
  wire [7:0] n36_I1_4_1; // @[Top.scala 165:21]
  wire [7:0] n36_I1_4_2; // @[Top.scala 165:21]
  wire [7:0] n36_I1_5_0; // @[Top.scala 165:21]
  wire [7:0] n36_I1_5_1; // @[Top.scala 165:21]
  wire [7:0] n36_I1_5_2; // @[Top.scala 165:21]
  wire [7:0] n36_I1_6_0; // @[Top.scala 165:21]
  wire [7:0] n36_I1_6_1; // @[Top.scala 165:21]
  wire [7:0] n36_I1_6_2; // @[Top.scala 165:21]
  wire [7:0] n36_I1_7_0; // @[Top.scala 165:21]
  wire [7:0] n36_I1_7_1; // @[Top.scala 165:21]
  wire [7:0] n36_I1_7_2; // @[Top.scala 165:21]
  wire [7:0] n36_I1_8_0; // @[Top.scala 165:21]
  wire [7:0] n36_I1_8_1; // @[Top.scala 165:21]
  wire [7:0] n36_I1_8_2; // @[Top.scala 165:21]
  wire [7:0] n36_I1_9_0; // @[Top.scala 165:21]
  wire [7:0] n36_I1_9_1; // @[Top.scala 165:21]
  wire [7:0] n36_I1_9_2; // @[Top.scala 165:21]
  wire [7:0] n36_I1_10_0; // @[Top.scala 165:21]
  wire [7:0] n36_I1_10_1; // @[Top.scala 165:21]
  wire [7:0] n36_I1_10_2; // @[Top.scala 165:21]
  wire [7:0] n36_I1_11_0; // @[Top.scala 165:21]
  wire [7:0] n36_I1_11_1; // @[Top.scala 165:21]
  wire [7:0] n36_I1_11_2; // @[Top.scala 165:21]
  wire [7:0] n36_I1_12_0; // @[Top.scala 165:21]
  wire [7:0] n36_I1_12_1; // @[Top.scala 165:21]
  wire [7:0] n36_I1_12_2; // @[Top.scala 165:21]
  wire [7:0] n36_I1_13_0; // @[Top.scala 165:21]
  wire [7:0] n36_I1_13_1; // @[Top.scala 165:21]
  wire [7:0] n36_I1_13_2; // @[Top.scala 165:21]
  wire [7:0] n36_I1_14_0; // @[Top.scala 165:21]
  wire [7:0] n36_I1_14_1; // @[Top.scala 165:21]
  wire [7:0] n36_I1_14_2; // @[Top.scala 165:21]
  wire [7:0] n36_I1_15_0; // @[Top.scala 165:21]
  wire [7:0] n36_I1_15_1; // @[Top.scala 165:21]
  wire [7:0] n36_I1_15_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_0_0_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_0_0_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_0_0_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_0_1_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_0_1_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_0_1_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_1_0_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_1_0_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_1_0_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_1_1_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_1_1_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_1_1_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_2_0_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_2_0_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_2_0_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_2_1_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_2_1_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_2_1_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_3_0_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_3_0_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_3_0_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_3_1_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_3_1_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_3_1_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_4_0_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_4_0_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_4_0_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_4_1_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_4_1_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_4_1_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_5_0_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_5_0_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_5_0_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_5_1_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_5_1_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_5_1_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_6_0_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_6_0_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_6_0_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_6_1_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_6_1_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_6_1_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_7_0_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_7_0_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_7_0_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_7_1_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_7_1_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_7_1_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_8_0_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_8_0_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_8_0_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_8_1_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_8_1_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_8_1_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_9_0_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_9_0_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_9_0_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_9_1_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_9_1_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_9_1_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_10_0_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_10_0_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_10_0_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_10_1_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_10_1_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_10_1_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_11_0_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_11_0_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_11_0_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_11_1_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_11_1_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_11_1_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_12_0_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_12_0_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_12_0_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_12_1_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_12_1_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_12_1_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_13_0_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_13_0_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_13_0_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_13_1_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_13_1_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_13_1_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_14_0_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_14_0_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_14_0_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_14_1_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_14_1_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_14_1_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_15_0_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_15_0_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_15_0_2; // @[Top.scala 165:21]
  wire [7:0] n36_O_15_1_0; // @[Top.scala 165:21]
  wire [7:0] n36_O_15_1_1; // @[Top.scala 165:21]
  wire [7:0] n36_O_15_1_2; // @[Top.scala 165:21]
  wire  n40_valid_up; // @[Top.scala 169:21]
  wire  n40_valid_down; // @[Top.scala 169:21]
  wire [7:0] n40_I_0; // @[Top.scala 169:21]
  wire [7:0] n40_I_1; // @[Top.scala 169:21]
  wire [7:0] n40_I_2; // @[Top.scala 169:21]
  wire [7:0] n40_I_3; // @[Top.scala 169:21]
  wire [7:0] n40_I_4; // @[Top.scala 169:21]
  wire [7:0] n40_I_5; // @[Top.scala 169:21]
  wire [7:0] n40_I_6; // @[Top.scala 169:21]
  wire [7:0] n40_I_7; // @[Top.scala 169:21]
  wire [7:0] n40_I_8; // @[Top.scala 169:21]
  wire [7:0] n40_I_9; // @[Top.scala 169:21]
  wire [7:0] n40_I_10; // @[Top.scala 169:21]
  wire [7:0] n40_I_11; // @[Top.scala 169:21]
  wire [7:0] n40_I_12; // @[Top.scala 169:21]
  wire [7:0] n40_I_13; // @[Top.scala 169:21]
  wire [7:0] n40_I_14; // @[Top.scala 169:21]
  wire [7:0] n40_I_15; // @[Top.scala 169:21]
  wire [7:0] n40_O_0; // @[Top.scala 169:21]
  wire [7:0] n40_O_1; // @[Top.scala 169:21]
  wire [7:0] n40_O_2; // @[Top.scala 169:21]
  wire [7:0] n40_O_3; // @[Top.scala 169:21]
  wire [7:0] n40_O_4; // @[Top.scala 169:21]
  wire [7:0] n40_O_5; // @[Top.scala 169:21]
  wire [7:0] n40_O_6; // @[Top.scala 169:21]
  wire [7:0] n40_O_7; // @[Top.scala 169:21]
  wire [7:0] n40_O_8; // @[Top.scala 169:21]
  wire [7:0] n40_O_9; // @[Top.scala 169:21]
  wire [7:0] n40_O_10; // @[Top.scala 169:21]
  wire [7:0] n40_O_11; // @[Top.scala 169:21]
  wire [7:0] n40_O_12; // @[Top.scala 169:21]
  wire [7:0] n40_O_13; // @[Top.scala 169:21]
  wire [7:0] n40_O_14; // @[Top.scala 169:21]
  wire [7:0] n40_O_15; // @[Top.scala 169:21]
  wire  n41_valid_up; // @[Top.scala 172:21]
  wire  n41_valid_down; // @[Top.scala 172:21]
  wire [7:0] n41_I_0; // @[Top.scala 172:21]
  wire [7:0] n41_I_1; // @[Top.scala 172:21]
  wire [7:0] n41_I_2; // @[Top.scala 172:21]
  wire [7:0] n41_I_3; // @[Top.scala 172:21]
  wire [7:0] n41_I_4; // @[Top.scala 172:21]
  wire [7:0] n41_I_5; // @[Top.scala 172:21]
  wire [7:0] n41_I_6; // @[Top.scala 172:21]
  wire [7:0] n41_I_7; // @[Top.scala 172:21]
  wire [7:0] n41_I_8; // @[Top.scala 172:21]
  wire [7:0] n41_I_9; // @[Top.scala 172:21]
  wire [7:0] n41_I_10; // @[Top.scala 172:21]
  wire [7:0] n41_I_11; // @[Top.scala 172:21]
  wire [7:0] n41_I_12; // @[Top.scala 172:21]
  wire [7:0] n41_I_13; // @[Top.scala 172:21]
  wire [7:0] n41_I_14; // @[Top.scala 172:21]
  wire [7:0] n41_I_15; // @[Top.scala 172:21]
  wire [7:0] n41_O_0; // @[Top.scala 172:21]
  wire [7:0] n41_O_1; // @[Top.scala 172:21]
  wire [7:0] n41_O_2; // @[Top.scala 172:21]
  wire [7:0] n41_O_3; // @[Top.scala 172:21]
  wire [7:0] n41_O_4; // @[Top.scala 172:21]
  wire [7:0] n41_O_5; // @[Top.scala 172:21]
  wire [7:0] n41_O_6; // @[Top.scala 172:21]
  wire [7:0] n41_O_7; // @[Top.scala 172:21]
  wire [7:0] n41_O_8; // @[Top.scala 172:21]
  wire [7:0] n41_O_9; // @[Top.scala 172:21]
  wire [7:0] n41_O_10; // @[Top.scala 172:21]
  wire [7:0] n41_O_11; // @[Top.scala 172:21]
  wire [7:0] n41_O_12; // @[Top.scala 172:21]
  wire [7:0] n41_O_13; // @[Top.scala 172:21]
  wire [7:0] n41_O_14; // @[Top.scala 172:21]
  wire [7:0] n41_O_15; // @[Top.scala 172:21]
  wire  n42_valid_up; // @[Top.scala 175:21]
  wire  n42_valid_down; // @[Top.scala 175:21]
  wire [7:0] n42_I0_0; // @[Top.scala 175:21]
  wire [7:0] n42_I0_1; // @[Top.scala 175:21]
  wire [7:0] n42_I0_2; // @[Top.scala 175:21]
  wire [7:0] n42_I0_3; // @[Top.scala 175:21]
  wire [7:0] n42_I0_4; // @[Top.scala 175:21]
  wire [7:0] n42_I0_5; // @[Top.scala 175:21]
  wire [7:0] n42_I0_6; // @[Top.scala 175:21]
  wire [7:0] n42_I0_7; // @[Top.scala 175:21]
  wire [7:0] n42_I0_8; // @[Top.scala 175:21]
  wire [7:0] n42_I0_9; // @[Top.scala 175:21]
  wire [7:0] n42_I0_10; // @[Top.scala 175:21]
  wire [7:0] n42_I0_11; // @[Top.scala 175:21]
  wire [7:0] n42_I0_12; // @[Top.scala 175:21]
  wire [7:0] n42_I0_13; // @[Top.scala 175:21]
  wire [7:0] n42_I0_14; // @[Top.scala 175:21]
  wire [7:0] n42_I0_15; // @[Top.scala 175:21]
  wire [7:0] n42_I1_0; // @[Top.scala 175:21]
  wire [7:0] n42_I1_1; // @[Top.scala 175:21]
  wire [7:0] n42_I1_2; // @[Top.scala 175:21]
  wire [7:0] n42_I1_3; // @[Top.scala 175:21]
  wire [7:0] n42_I1_4; // @[Top.scala 175:21]
  wire [7:0] n42_I1_5; // @[Top.scala 175:21]
  wire [7:0] n42_I1_6; // @[Top.scala 175:21]
  wire [7:0] n42_I1_7; // @[Top.scala 175:21]
  wire [7:0] n42_I1_8; // @[Top.scala 175:21]
  wire [7:0] n42_I1_9; // @[Top.scala 175:21]
  wire [7:0] n42_I1_10; // @[Top.scala 175:21]
  wire [7:0] n42_I1_11; // @[Top.scala 175:21]
  wire [7:0] n42_I1_12; // @[Top.scala 175:21]
  wire [7:0] n42_I1_13; // @[Top.scala 175:21]
  wire [7:0] n42_I1_14; // @[Top.scala 175:21]
  wire [7:0] n42_I1_15; // @[Top.scala 175:21]
  wire [7:0] n42_O_0_0; // @[Top.scala 175:21]
  wire [7:0] n42_O_0_1; // @[Top.scala 175:21]
  wire [7:0] n42_O_1_0; // @[Top.scala 175:21]
  wire [7:0] n42_O_1_1; // @[Top.scala 175:21]
  wire [7:0] n42_O_2_0; // @[Top.scala 175:21]
  wire [7:0] n42_O_2_1; // @[Top.scala 175:21]
  wire [7:0] n42_O_3_0; // @[Top.scala 175:21]
  wire [7:0] n42_O_3_1; // @[Top.scala 175:21]
  wire [7:0] n42_O_4_0; // @[Top.scala 175:21]
  wire [7:0] n42_O_4_1; // @[Top.scala 175:21]
  wire [7:0] n42_O_5_0; // @[Top.scala 175:21]
  wire [7:0] n42_O_5_1; // @[Top.scala 175:21]
  wire [7:0] n42_O_6_0; // @[Top.scala 175:21]
  wire [7:0] n42_O_6_1; // @[Top.scala 175:21]
  wire [7:0] n42_O_7_0; // @[Top.scala 175:21]
  wire [7:0] n42_O_7_1; // @[Top.scala 175:21]
  wire [7:0] n42_O_8_0; // @[Top.scala 175:21]
  wire [7:0] n42_O_8_1; // @[Top.scala 175:21]
  wire [7:0] n42_O_9_0; // @[Top.scala 175:21]
  wire [7:0] n42_O_9_1; // @[Top.scala 175:21]
  wire [7:0] n42_O_10_0; // @[Top.scala 175:21]
  wire [7:0] n42_O_10_1; // @[Top.scala 175:21]
  wire [7:0] n42_O_11_0; // @[Top.scala 175:21]
  wire [7:0] n42_O_11_1; // @[Top.scala 175:21]
  wire [7:0] n42_O_12_0; // @[Top.scala 175:21]
  wire [7:0] n42_O_12_1; // @[Top.scala 175:21]
  wire [7:0] n42_O_13_0; // @[Top.scala 175:21]
  wire [7:0] n42_O_13_1; // @[Top.scala 175:21]
  wire [7:0] n42_O_14_0; // @[Top.scala 175:21]
  wire [7:0] n42_O_14_1; // @[Top.scala 175:21]
  wire [7:0] n42_O_15_0; // @[Top.scala 175:21]
  wire [7:0] n42_O_15_1; // @[Top.scala 175:21]
  wire  n46_valid_up; // @[Top.scala 179:21]
  wire  n46_valid_down; // @[Top.scala 179:21]
  wire [7:0] n46_I0_0_0; // @[Top.scala 179:21]
  wire [7:0] n46_I0_0_1; // @[Top.scala 179:21]
  wire [7:0] n46_I0_1_0; // @[Top.scala 179:21]
  wire [7:0] n46_I0_1_1; // @[Top.scala 179:21]
  wire [7:0] n46_I0_2_0; // @[Top.scala 179:21]
  wire [7:0] n46_I0_2_1; // @[Top.scala 179:21]
  wire [7:0] n46_I0_3_0; // @[Top.scala 179:21]
  wire [7:0] n46_I0_3_1; // @[Top.scala 179:21]
  wire [7:0] n46_I0_4_0; // @[Top.scala 179:21]
  wire [7:0] n46_I0_4_1; // @[Top.scala 179:21]
  wire [7:0] n46_I0_5_0; // @[Top.scala 179:21]
  wire [7:0] n46_I0_5_1; // @[Top.scala 179:21]
  wire [7:0] n46_I0_6_0; // @[Top.scala 179:21]
  wire [7:0] n46_I0_6_1; // @[Top.scala 179:21]
  wire [7:0] n46_I0_7_0; // @[Top.scala 179:21]
  wire [7:0] n46_I0_7_1; // @[Top.scala 179:21]
  wire [7:0] n46_I0_8_0; // @[Top.scala 179:21]
  wire [7:0] n46_I0_8_1; // @[Top.scala 179:21]
  wire [7:0] n46_I0_9_0; // @[Top.scala 179:21]
  wire [7:0] n46_I0_9_1; // @[Top.scala 179:21]
  wire [7:0] n46_I0_10_0; // @[Top.scala 179:21]
  wire [7:0] n46_I0_10_1; // @[Top.scala 179:21]
  wire [7:0] n46_I0_11_0; // @[Top.scala 179:21]
  wire [7:0] n46_I0_11_1; // @[Top.scala 179:21]
  wire [7:0] n46_I0_12_0; // @[Top.scala 179:21]
  wire [7:0] n46_I0_12_1; // @[Top.scala 179:21]
  wire [7:0] n46_I0_13_0; // @[Top.scala 179:21]
  wire [7:0] n46_I0_13_1; // @[Top.scala 179:21]
  wire [7:0] n46_I0_14_0; // @[Top.scala 179:21]
  wire [7:0] n46_I0_14_1; // @[Top.scala 179:21]
  wire [7:0] n46_I0_15_0; // @[Top.scala 179:21]
  wire [7:0] n46_I0_15_1; // @[Top.scala 179:21]
  wire [7:0] n46_I1_0; // @[Top.scala 179:21]
  wire [7:0] n46_I1_1; // @[Top.scala 179:21]
  wire [7:0] n46_I1_2; // @[Top.scala 179:21]
  wire [7:0] n46_I1_3; // @[Top.scala 179:21]
  wire [7:0] n46_I1_4; // @[Top.scala 179:21]
  wire [7:0] n46_I1_5; // @[Top.scala 179:21]
  wire [7:0] n46_I1_6; // @[Top.scala 179:21]
  wire [7:0] n46_I1_7; // @[Top.scala 179:21]
  wire [7:0] n46_I1_8; // @[Top.scala 179:21]
  wire [7:0] n46_I1_9; // @[Top.scala 179:21]
  wire [7:0] n46_I1_10; // @[Top.scala 179:21]
  wire [7:0] n46_I1_11; // @[Top.scala 179:21]
  wire [7:0] n46_I1_12; // @[Top.scala 179:21]
  wire [7:0] n46_I1_13; // @[Top.scala 179:21]
  wire [7:0] n46_I1_14; // @[Top.scala 179:21]
  wire [7:0] n46_I1_15; // @[Top.scala 179:21]
  wire [7:0] n46_O_0_0; // @[Top.scala 179:21]
  wire [7:0] n46_O_0_1; // @[Top.scala 179:21]
  wire [7:0] n46_O_0_2; // @[Top.scala 179:21]
  wire [7:0] n46_O_1_0; // @[Top.scala 179:21]
  wire [7:0] n46_O_1_1; // @[Top.scala 179:21]
  wire [7:0] n46_O_1_2; // @[Top.scala 179:21]
  wire [7:0] n46_O_2_0; // @[Top.scala 179:21]
  wire [7:0] n46_O_2_1; // @[Top.scala 179:21]
  wire [7:0] n46_O_2_2; // @[Top.scala 179:21]
  wire [7:0] n46_O_3_0; // @[Top.scala 179:21]
  wire [7:0] n46_O_3_1; // @[Top.scala 179:21]
  wire [7:0] n46_O_3_2; // @[Top.scala 179:21]
  wire [7:0] n46_O_4_0; // @[Top.scala 179:21]
  wire [7:0] n46_O_4_1; // @[Top.scala 179:21]
  wire [7:0] n46_O_4_2; // @[Top.scala 179:21]
  wire [7:0] n46_O_5_0; // @[Top.scala 179:21]
  wire [7:0] n46_O_5_1; // @[Top.scala 179:21]
  wire [7:0] n46_O_5_2; // @[Top.scala 179:21]
  wire [7:0] n46_O_6_0; // @[Top.scala 179:21]
  wire [7:0] n46_O_6_1; // @[Top.scala 179:21]
  wire [7:0] n46_O_6_2; // @[Top.scala 179:21]
  wire [7:0] n46_O_7_0; // @[Top.scala 179:21]
  wire [7:0] n46_O_7_1; // @[Top.scala 179:21]
  wire [7:0] n46_O_7_2; // @[Top.scala 179:21]
  wire [7:0] n46_O_8_0; // @[Top.scala 179:21]
  wire [7:0] n46_O_8_1; // @[Top.scala 179:21]
  wire [7:0] n46_O_8_2; // @[Top.scala 179:21]
  wire [7:0] n46_O_9_0; // @[Top.scala 179:21]
  wire [7:0] n46_O_9_1; // @[Top.scala 179:21]
  wire [7:0] n46_O_9_2; // @[Top.scala 179:21]
  wire [7:0] n46_O_10_0; // @[Top.scala 179:21]
  wire [7:0] n46_O_10_1; // @[Top.scala 179:21]
  wire [7:0] n46_O_10_2; // @[Top.scala 179:21]
  wire [7:0] n46_O_11_0; // @[Top.scala 179:21]
  wire [7:0] n46_O_11_1; // @[Top.scala 179:21]
  wire [7:0] n46_O_11_2; // @[Top.scala 179:21]
  wire [7:0] n46_O_12_0; // @[Top.scala 179:21]
  wire [7:0] n46_O_12_1; // @[Top.scala 179:21]
  wire [7:0] n46_O_12_2; // @[Top.scala 179:21]
  wire [7:0] n46_O_13_0; // @[Top.scala 179:21]
  wire [7:0] n46_O_13_1; // @[Top.scala 179:21]
  wire [7:0] n46_O_13_2; // @[Top.scala 179:21]
  wire [7:0] n46_O_14_0; // @[Top.scala 179:21]
  wire [7:0] n46_O_14_1; // @[Top.scala 179:21]
  wire [7:0] n46_O_14_2; // @[Top.scala 179:21]
  wire [7:0] n46_O_15_0; // @[Top.scala 179:21]
  wire [7:0] n46_O_15_1; // @[Top.scala 179:21]
  wire [7:0] n46_O_15_2; // @[Top.scala 179:21]
  wire  n50_valid_up; // @[Top.scala 183:21]
  wire  n50_valid_down; // @[Top.scala 183:21]
  wire [7:0] n50_I_0_0; // @[Top.scala 183:21]
  wire [7:0] n50_I_0_1; // @[Top.scala 183:21]
  wire [7:0] n50_I_0_2; // @[Top.scala 183:21]
  wire [7:0] n50_I_1_0; // @[Top.scala 183:21]
  wire [7:0] n50_I_1_1; // @[Top.scala 183:21]
  wire [7:0] n50_I_1_2; // @[Top.scala 183:21]
  wire [7:0] n50_I_2_0; // @[Top.scala 183:21]
  wire [7:0] n50_I_2_1; // @[Top.scala 183:21]
  wire [7:0] n50_I_2_2; // @[Top.scala 183:21]
  wire [7:0] n50_I_3_0; // @[Top.scala 183:21]
  wire [7:0] n50_I_3_1; // @[Top.scala 183:21]
  wire [7:0] n50_I_3_2; // @[Top.scala 183:21]
  wire [7:0] n50_I_4_0; // @[Top.scala 183:21]
  wire [7:0] n50_I_4_1; // @[Top.scala 183:21]
  wire [7:0] n50_I_4_2; // @[Top.scala 183:21]
  wire [7:0] n50_I_5_0; // @[Top.scala 183:21]
  wire [7:0] n50_I_5_1; // @[Top.scala 183:21]
  wire [7:0] n50_I_5_2; // @[Top.scala 183:21]
  wire [7:0] n50_I_6_0; // @[Top.scala 183:21]
  wire [7:0] n50_I_6_1; // @[Top.scala 183:21]
  wire [7:0] n50_I_6_2; // @[Top.scala 183:21]
  wire [7:0] n50_I_7_0; // @[Top.scala 183:21]
  wire [7:0] n50_I_7_1; // @[Top.scala 183:21]
  wire [7:0] n50_I_7_2; // @[Top.scala 183:21]
  wire [7:0] n50_I_8_0; // @[Top.scala 183:21]
  wire [7:0] n50_I_8_1; // @[Top.scala 183:21]
  wire [7:0] n50_I_8_2; // @[Top.scala 183:21]
  wire [7:0] n50_I_9_0; // @[Top.scala 183:21]
  wire [7:0] n50_I_9_1; // @[Top.scala 183:21]
  wire [7:0] n50_I_9_2; // @[Top.scala 183:21]
  wire [7:0] n50_I_10_0; // @[Top.scala 183:21]
  wire [7:0] n50_I_10_1; // @[Top.scala 183:21]
  wire [7:0] n50_I_10_2; // @[Top.scala 183:21]
  wire [7:0] n50_I_11_0; // @[Top.scala 183:21]
  wire [7:0] n50_I_11_1; // @[Top.scala 183:21]
  wire [7:0] n50_I_11_2; // @[Top.scala 183:21]
  wire [7:0] n50_I_12_0; // @[Top.scala 183:21]
  wire [7:0] n50_I_12_1; // @[Top.scala 183:21]
  wire [7:0] n50_I_12_2; // @[Top.scala 183:21]
  wire [7:0] n50_I_13_0; // @[Top.scala 183:21]
  wire [7:0] n50_I_13_1; // @[Top.scala 183:21]
  wire [7:0] n50_I_13_2; // @[Top.scala 183:21]
  wire [7:0] n50_I_14_0; // @[Top.scala 183:21]
  wire [7:0] n50_I_14_1; // @[Top.scala 183:21]
  wire [7:0] n50_I_14_2; // @[Top.scala 183:21]
  wire [7:0] n50_I_15_0; // @[Top.scala 183:21]
  wire [7:0] n50_I_15_1; // @[Top.scala 183:21]
  wire [7:0] n50_I_15_2; // @[Top.scala 183:21]
  wire [7:0] n50_O_0_0_0; // @[Top.scala 183:21]
  wire [7:0] n50_O_0_0_1; // @[Top.scala 183:21]
  wire [7:0] n50_O_0_0_2; // @[Top.scala 183:21]
  wire [7:0] n50_O_1_0_0; // @[Top.scala 183:21]
  wire [7:0] n50_O_1_0_1; // @[Top.scala 183:21]
  wire [7:0] n50_O_1_0_2; // @[Top.scala 183:21]
  wire [7:0] n50_O_2_0_0; // @[Top.scala 183:21]
  wire [7:0] n50_O_2_0_1; // @[Top.scala 183:21]
  wire [7:0] n50_O_2_0_2; // @[Top.scala 183:21]
  wire [7:0] n50_O_3_0_0; // @[Top.scala 183:21]
  wire [7:0] n50_O_3_0_1; // @[Top.scala 183:21]
  wire [7:0] n50_O_3_0_2; // @[Top.scala 183:21]
  wire [7:0] n50_O_4_0_0; // @[Top.scala 183:21]
  wire [7:0] n50_O_4_0_1; // @[Top.scala 183:21]
  wire [7:0] n50_O_4_0_2; // @[Top.scala 183:21]
  wire [7:0] n50_O_5_0_0; // @[Top.scala 183:21]
  wire [7:0] n50_O_5_0_1; // @[Top.scala 183:21]
  wire [7:0] n50_O_5_0_2; // @[Top.scala 183:21]
  wire [7:0] n50_O_6_0_0; // @[Top.scala 183:21]
  wire [7:0] n50_O_6_0_1; // @[Top.scala 183:21]
  wire [7:0] n50_O_6_0_2; // @[Top.scala 183:21]
  wire [7:0] n50_O_7_0_0; // @[Top.scala 183:21]
  wire [7:0] n50_O_7_0_1; // @[Top.scala 183:21]
  wire [7:0] n50_O_7_0_2; // @[Top.scala 183:21]
  wire [7:0] n50_O_8_0_0; // @[Top.scala 183:21]
  wire [7:0] n50_O_8_0_1; // @[Top.scala 183:21]
  wire [7:0] n50_O_8_0_2; // @[Top.scala 183:21]
  wire [7:0] n50_O_9_0_0; // @[Top.scala 183:21]
  wire [7:0] n50_O_9_0_1; // @[Top.scala 183:21]
  wire [7:0] n50_O_9_0_2; // @[Top.scala 183:21]
  wire [7:0] n50_O_10_0_0; // @[Top.scala 183:21]
  wire [7:0] n50_O_10_0_1; // @[Top.scala 183:21]
  wire [7:0] n50_O_10_0_2; // @[Top.scala 183:21]
  wire [7:0] n50_O_11_0_0; // @[Top.scala 183:21]
  wire [7:0] n50_O_11_0_1; // @[Top.scala 183:21]
  wire [7:0] n50_O_11_0_2; // @[Top.scala 183:21]
  wire [7:0] n50_O_12_0_0; // @[Top.scala 183:21]
  wire [7:0] n50_O_12_0_1; // @[Top.scala 183:21]
  wire [7:0] n50_O_12_0_2; // @[Top.scala 183:21]
  wire [7:0] n50_O_13_0_0; // @[Top.scala 183:21]
  wire [7:0] n50_O_13_0_1; // @[Top.scala 183:21]
  wire [7:0] n50_O_13_0_2; // @[Top.scala 183:21]
  wire [7:0] n50_O_14_0_0; // @[Top.scala 183:21]
  wire [7:0] n50_O_14_0_1; // @[Top.scala 183:21]
  wire [7:0] n50_O_14_0_2; // @[Top.scala 183:21]
  wire [7:0] n50_O_15_0_0; // @[Top.scala 183:21]
  wire [7:0] n50_O_15_0_1; // @[Top.scala 183:21]
  wire [7:0] n50_O_15_0_2; // @[Top.scala 183:21]
  wire  n55_valid_up; // @[Top.scala 186:21]
  wire  n55_valid_down; // @[Top.scala 186:21]
  wire [7:0] n55_I_0_0_0; // @[Top.scala 186:21]
  wire [7:0] n55_I_0_0_1; // @[Top.scala 186:21]
  wire [7:0] n55_I_0_0_2; // @[Top.scala 186:21]
  wire [7:0] n55_I_1_0_0; // @[Top.scala 186:21]
  wire [7:0] n55_I_1_0_1; // @[Top.scala 186:21]
  wire [7:0] n55_I_1_0_2; // @[Top.scala 186:21]
  wire [7:0] n55_I_2_0_0; // @[Top.scala 186:21]
  wire [7:0] n55_I_2_0_1; // @[Top.scala 186:21]
  wire [7:0] n55_I_2_0_2; // @[Top.scala 186:21]
  wire [7:0] n55_I_3_0_0; // @[Top.scala 186:21]
  wire [7:0] n55_I_3_0_1; // @[Top.scala 186:21]
  wire [7:0] n55_I_3_0_2; // @[Top.scala 186:21]
  wire [7:0] n55_I_4_0_0; // @[Top.scala 186:21]
  wire [7:0] n55_I_4_0_1; // @[Top.scala 186:21]
  wire [7:0] n55_I_4_0_2; // @[Top.scala 186:21]
  wire [7:0] n55_I_5_0_0; // @[Top.scala 186:21]
  wire [7:0] n55_I_5_0_1; // @[Top.scala 186:21]
  wire [7:0] n55_I_5_0_2; // @[Top.scala 186:21]
  wire [7:0] n55_I_6_0_0; // @[Top.scala 186:21]
  wire [7:0] n55_I_6_0_1; // @[Top.scala 186:21]
  wire [7:0] n55_I_6_0_2; // @[Top.scala 186:21]
  wire [7:0] n55_I_7_0_0; // @[Top.scala 186:21]
  wire [7:0] n55_I_7_0_1; // @[Top.scala 186:21]
  wire [7:0] n55_I_7_0_2; // @[Top.scala 186:21]
  wire [7:0] n55_I_8_0_0; // @[Top.scala 186:21]
  wire [7:0] n55_I_8_0_1; // @[Top.scala 186:21]
  wire [7:0] n55_I_8_0_2; // @[Top.scala 186:21]
  wire [7:0] n55_I_9_0_0; // @[Top.scala 186:21]
  wire [7:0] n55_I_9_0_1; // @[Top.scala 186:21]
  wire [7:0] n55_I_9_0_2; // @[Top.scala 186:21]
  wire [7:0] n55_I_10_0_0; // @[Top.scala 186:21]
  wire [7:0] n55_I_10_0_1; // @[Top.scala 186:21]
  wire [7:0] n55_I_10_0_2; // @[Top.scala 186:21]
  wire [7:0] n55_I_11_0_0; // @[Top.scala 186:21]
  wire [7:0] n55_I_11_0_1; // @[Top.scala 186:21]
  wire [7:0] n55_I_11_0_2; // @[Top.scala 186:21]
  wire [7:0] n55_I_12_0_0; // @[Top.scala 186:21]
  wire [7:0] n55_I_12_0_1; // @[Top.scala 186:21]
  wire [7:0] n55_I_12_0_2; // @[Top.scala 186:21]
  wire [7:0] n55_I_13_0_0; // @[Top.scala 186:21]
  wire [7:0] n55_I_13_0_1; // @[Top.scala 186:21]
  wire [7:0] n55_I_13_0_2; // @[Top.scala 186:21]
  wire [7:0] n55_I_14_0_0; // @[Top.scala 186:21]
  wire [7:0] n55_I_14_0_1; // @[Top.scala 186:21]
  wire [7:0] n55_I_14_0_2; // @[Top.scala 186:21]
  wire [7:0] n55_I_15_0_0; // @[Top.scala 186:21]
  wire [7:0] n55_I_15_0_1; // @[Top.scala 186:21]
  wire [7:0] n55_I_15_0_2; // @[Top.scala 186:21]
  wire [7:0] n55_O_0_0; // @[Top.scala 186:21]
  wire [7:0] n55_O_0_1; // @[Top.scala 186:21]
  wire [7:0] n55_O_0_2; // @[Top.scala 186:21]
  wire [7:0] n55_O_1_0; // @[Top.scala 186:21]
  wire [7:0] n55_O_1_1; // @[Top.scala 186:21]
  wire [7:0] n55_O_1_2; // @[Top.scala 186:21]
  wire [7:0] n55_O_2_0; // @[Top.scala 186:21]
  wire [7:0] n55_O_2_1; // @[Top.scala 186:21]
  wire [7:0] n55_O_2_2; // @[Top.scala 186:21]
  wire [7:0] n55_O_3_0; // @[Top.scala 186:21]
  wire [7:0] n55_O_3_1; // @[Top.scala 186:21]
  wire [7:0] n55_O_3_2; // @[Top.scala 186:21]
  wire [7:0] n55_O_4_0; // @[Top.scala 186:21]
  wire [7:0] n55_O_4_1; // @[Top.scala 186:21]
  wire [7:0] n55_O_4_2; // @[Top.scala 186:21]
  wire [7:0] n55_O_5_0; // @[Top.scala 186:21]
  wire [7:0] n55_O_5_1; // @[Top.scala 186:21]
  wire [7:0] n55_O_5_2; // @[Top.scala 186:21]
  wire [7:0] n55_O_6_0; // @[Top.scala 186:21]
  wire [7:0] n55_O_6_1; // @[Top.scala 186:21]
  wire [7:0] n55_O_6_2; // @[Top.scala 186:21]
  wire [7:0] n55_O_7_0; // @[Top.scala 186:21]
  wire [7:0] n55_O_7_1; // @[Top.scala 186:21]
  wire [7:0] n55_O_7_2; // @[Top.scala 186:21]
  wire [7:0] n55_O_8_0; // @[Top.scala 186:21]
  wire [7:0] n55_O_8_1; // @[Top.scala 186:21]
  wire [7:0] n55_O_8_2; // @[Top.scala 186:21]
  wire [7:0] n55_O_9_0; // @[Top.scala 186:21]
  wire [7:0] n55_O_9_1; // @[Top.scala 186:21]
  wire [7:0] n55_O_9_2; // @[Top.scala 186:21]
  wire [7:0] n55_O_10_0; // @[Top.scala 186:21]
  wire [7:0] n55_O_10_1; // @[Top.scala 186:21]
  wire [7:0] n55_O_10_2; // @[Top.scala 186:21]
  wire [7:0] n55_O_11_0; // @[Top.scala 186:21]
  wire [7:0] n55_O_11_1; // @[Top.scala 186:21]
  wire [7:0] n55_O_11_2; // @[Top.scala 186:21]
  wire [7:0] n55_O_12_0; // @[Top.scala 186:21]
  wire [7:0] n55_O_12_1; // @[Top.scala 186:21]
  wire [7:0] n55_O_12_2; // @[Top.scala 186:21]
  wire [7:0] n55_O_13_0; // @[Top.scala 186:21]
  wire [7:0] n55_O_13_1; // @[Top.scala 186:21]
  wire [7:0] n55_O_13_2; // @[Top.scala 186:21]
  wire [7:0] n55_O_14_0; // @[Top.scala 186:21]
  wire [7:0] n55_O_14_1; // @[Top.scala 186:21]
  wire [7:0] n55_O_14_2; // @[Top.scala 186:21]
  wire [7:0] n55_O_15_0; // @[Top.scala 186:21]
  wire [7:0] n55_O_15_1; // @[Top.scala 186:21]
  wire [7:0] n55_O_15_2; // @[Top.scala 186:21]
  wire  n56_valid_up; // @[Top.scala 189:21]
  wire  n56_valid_down; // @[Top.scala 189:21]
  wire [7:0] n56_I0_0_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_0_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_0_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_0_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_0_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_0_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_1_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_1_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_1_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_1_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_1_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_1_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_2_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_2_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_2_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_2_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_2_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_2_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_3_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_3_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_3_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_3_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_3_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_3_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_4_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_4_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_4_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_4_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_4_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_4_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_5_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_5_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_5_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_5_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_5_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_5_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_6_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_6_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_6_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_6_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_6_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_6_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_7_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_7_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_7_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_7_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_7_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_7_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_8_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_8_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_8_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_8_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_8_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_8_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_9_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_9_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_9_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_9_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_9_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_9_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_10_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_10_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_10_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_10_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_10_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_10_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_11_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_11_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_11_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_11_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_11_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_11_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_12_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_12_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_12_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_12_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_12_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_12_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_13_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_13_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_13_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_13_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_13_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_13_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_14_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_14_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_14_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_14_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_14_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_14_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_15_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_15_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_15_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_I0_15_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_I0_15_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_I0_15_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_I1_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_I1_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_I1_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_I1_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_I1_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_I1_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_I1_2_0; // @[Top.scala 189:21]
  wire [7:0] n56_I1_2_1; // @[Top.scala 189:21]
  wire [7:0] n56_I1_2_2; // @[Top.scala 189:21]
  wire [7:0] n56_I1_3_0; // @[Top.scala 189:21]
  wire [7:0] n56_I1_3_1; // @[Top.scala 189:21]
  wire [7:0] n56_I1_3_2; // @[Top.scala 189:21]
  wire [7:0] n56_I1_4_0; // @[Top.scala 189:21]
  wire [7:0] n56_I1_4_1; // @[Top.scala 189:21]
  wire [7:0] n56_I1_4_2; // @[Top.scala 189:21]
  wire [7:0] n56_I1_5_0; // @[Top.scala 189:21]
  wire [7:0] n56_I1_5_1; // @[Top.scala 189:21]
  wire [7:0] n56_I1_5_2; // @[Top.scala 189:21]
  wire [7:0] n56_I1_6_0; // @[Top.scala 189:21]
  wire [7:0] n56_I1_6_1; // @[Top.scala 189:21]
  wire [7:0] n56_I1_6_2; // @[Top.scala 189:21]
  wire [7:0] n56_I1_7_0; // @[Top.scala 189:21]
  wire [7:0] n56_I1_7_1; // @[Top.scala 189:21]
  wire [7:0] n56_I1_7_2; // @[Top.scala 189:21]
  wire [7:0] n56_I1_8_0; // @[Top.scala 189:21]
  wire [7:0] n56_I1_8_1; // @[Top.scala 189:21]
  wire [7:0] n56_I1_8_2; // @[Top.scala 189:21]
  wire [7:0] n56_I1_9_0; // @[Top.scala 189:21]
  wire [7:0] n56_I1_9_1; // @[Top.scala 189:21]
  wire [7:0] n56_I1_9_2; // @[Top.scala 189:21]
  wire [7:0] n56_I1_10_0; // @[Top.scala 189:21]
  wire [7:0] n56_I1_10_1; // @[Top.scala 189:21]
  wire [7:0] n56_I1_10_2; // @[Top.scala 189:21]
  wire [7:0] n56_I1_11_0; // @[Top.scala 189:21]
  wire [7:0] n56_I1_11_1; // @[Top.scala 189:21]
  wire [7:0] n56_I1_11_2; // @[Top.scala 189:21]
  wire [7:0] n56_I1_12_0; // @[Top.scala 189:21]
  wire [7:0] n56_I1_12_1; // @[Top.scala 189:21]
  wire [7:0] n56_I1_12_2; // @[Top.scala 189:21]
  wire [7:0] n56_I1_13_0; // @[Top.scala 189:21]
  wire [7:0] n56_I1_13_1; // @[Top.scala 189:21]
  wire [7:0] n56_I1_13_2; // @[Top.scala 189:21]
  wire [7:0] n56_I1_14_0; // @[Top.scala 189:21]
  wire [7:0] n56_I1_14_1; // @[Top.scala 189:21]
  wire [7:0] n56_I1_14_2; // @[Top.scala 189:21]
  wire [7:0] n56_I1_15_0; // @[Top.scala 189:21]
  wire [7:0] n56_I1_15_1; // @[Top.scala 189:21]
  wire [7:0] n56_I1_15_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_0_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_0_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_0_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_0_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_0_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_0_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_0_2_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_0_2_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_0_2_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_1_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_1_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_1_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_1_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_1_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_1_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_1_2_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_1_2_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_1_2_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_2_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_2_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_2_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_2_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_2_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_2_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_2_2_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_2_2_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_2_2_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_3_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_3_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_3_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_3_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_3_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_3_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_3_2_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_3_2_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_3_2_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_4_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_4_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_4_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_4_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_4_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_4_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_4_2_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_4_2_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_4_2_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_5_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_5_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_5_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_5_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_5_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_5_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_5_2_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_5_2_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_5_2_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_6_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_6_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_6_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_6_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_6_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_6_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_6_2_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_6_2_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_6_2_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_7_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_7_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_7_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_7_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_7_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_7_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_7_2_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_7_2_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_7_2_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_8_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_8_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_8_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_8_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_8_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_8_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_8_2_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_8_2_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_8_2_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_9_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_9_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_9_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_9_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_9_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_9_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_9_2_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_9_2_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_9_2_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_10_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_10_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_10_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_10_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_10_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_10_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_10_2_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_10_2_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_10_2_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_11_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_11_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_11_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_11_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_11_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_11_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_11_2_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_11_2_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_11_2_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_12_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_12_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_12_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_12_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_12_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_12_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_12_2_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_12_2_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_12_2_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_13_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_13_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_13_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_13_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_13_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_13_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_13_2_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_13_2_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_13_2_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_14_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_14_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_14_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_14_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_14_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_14_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_14_2_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_14_2_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_14_2_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_15_0_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_15_0_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_15_0_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_15_1_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_15_1_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_15_1_2; // @[Top.scala 189:21]
  wire [7:0] n56_O_15_2_0; // @[Top.scala 189:21]
  wire [7:0] n56_O_15_2_1; // @[Top.scala 189:21]
  wire [7:0] n56_O_15_2_2; // @[Top.scala 189:21]
  wire  n60_valid_up; // @[Top.scala 193:21]
  wire  n60_valid_down; // @[Top.scala 193:21]
  wire [7:0] n60_I_0_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_0_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_0_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_0_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_0_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_0_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_0_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_0_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_0_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_1_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_1_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_1_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_1_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_1_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_1_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_1_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_1_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_1_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_2_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_2_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_2_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_2_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_2_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_2_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_2_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_2_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_2_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_3_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_3_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_3_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_3_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_3_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_3_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_3_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_3_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_3_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_4_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_4_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_4_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_4_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_4_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_4_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_4_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_4_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_4_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_5_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_5_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_5_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_5_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_5_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_5_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_5_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_5_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_5_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_6_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_6_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_6_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_6_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_6_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_6_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_6_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_6_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_6_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_7_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_7_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_7_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_7_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_7_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_7_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_7_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_7_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_7_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_8_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_8_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_8_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_8_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_8_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_8_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_8_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_8_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_8_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_9_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_9_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_9_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_9_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_9_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_9_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_9_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_9_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_9_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_10_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_10_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_10_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_10_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_10_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_10_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_10_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_10_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_10_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_11_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_11_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_11_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_11_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_11_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_11_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_11_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_11_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_11_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_12_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_12_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_12_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_12_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_12_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_12_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_12_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_12_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_12_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_13_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_13_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_13_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_13_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_13_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_13_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_13_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_13_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_13_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_14_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_14_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_14_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_14_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_14_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_14_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_14_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_14_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_14_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_15_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_15_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_15_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_15_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_15_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_15_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_I_15_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_I_15_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_I_15_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_0_0_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_0_0_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_0_0_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_0_0_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_0_0_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_0_0_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_0_0_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_0_0_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_0_0_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_1_0_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_1_0_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_1_0_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_1_0_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_1_0_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_1_0_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_1_0_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_1_0_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_1_0_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_2_0_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_2_0_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_2_0_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_2_0_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_2_0_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_2_0_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_2_0_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_2_0_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_2_0_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_3_0_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_3_0_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_3_0_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_3_0_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_3_0_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_3_0_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_3_0_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_3_0_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_3_0_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_4_0_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_4_0_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_4_0_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_4_0_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_4_0_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_4_0_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_4_0_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_4_0_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_4_0_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_5_0_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_5_0_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_5_0_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_5_0_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_5_0_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_5_0_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_5_0_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_5_0_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_5_0_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_6_0_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_6_0_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_6_0_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_6_0_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_6_0_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_6_0_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_6_0_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_6_0_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_6_0_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_7_0_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_7_0_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_7_0_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_7_0_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_7_0_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_7_0_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_7_0_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_7_0_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_7_0_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_8_0_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_8_0_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_8_0_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_8_0_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_8_0_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_8_0_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_8_0_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_8_0_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_8_0_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_9_0_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_9_0_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_9_0_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_9_0_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_9_0_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_9_0_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_9_0_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_9_0_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_9_0_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_10_0_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_10_0_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_10_0_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_10_0_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_10_0_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_10_0_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_10_0_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_10_0_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_10_0_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_11_0_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_11_0_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_11_0_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_11_0_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_11_0_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_11_0_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_11_0_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_11_0_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_11_0_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_12_0_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_12_0_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_12_0_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_12_0_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_12_0_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_12_0_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_12_0_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_12_0_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_12_0_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_13_0_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_13_0_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_13_0_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_13_0_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_13_0_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_13_0_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_13_0_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_13_0_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_13_0_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_14_0_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_14_0_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_14_0_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_14_0_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_14_0_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_14_0_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_14_0_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_14_0_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_14_0_2_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_15_0_0_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_15_0_0_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_15_0_0_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_15_0_1_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_15_0_1_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_15_0_1_2; // @[Top.scala 193:21]
  wire [7:0] n60_O_15_0_2_0; // @[Top.scala 193:21]
  wire [7:0] n60_O_15_0_2_1; // @[Top.scala 193:21]
  wire [7:0] n60_O_15_0_2_2; // @[Top.scala 193:21]
  wire  n65_valid_up; // @[Top.scala 196:21]
  wire  n65_valid_down; // @[Top.scala 196:21]
  wire [7:0] n65_I_0_0_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_0_0_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_0_0_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_0_0_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_0_0_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_0_0_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_0_0_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_0_0_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_0_0_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_1_0_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_1_0_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_1_0_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_1_0_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_1_0_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_1_0_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_1_0_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_1_0_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_1_0_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_2_0_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_2_0_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_2_0_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_2_0_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_2_0_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_2_0_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_2_0_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_2_0_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_2_0_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_3_0_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_3_0_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_3_0_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_3_0_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_3_0_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_3_0_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_3_0_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_3_0_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_3_0_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_4_0_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_4_0_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_4_0_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_4_0_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_4_0_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_4_0_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_4_0_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_4_0_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_4_0_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_5_0_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_5_0_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_5_0_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_5_0_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_5_0_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_5_0_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_5_0_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_5_0_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_5_0_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_6_0_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_6_0_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_6_0_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_6_0_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_6_0_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_6_0_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_6_0_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_6_0_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_6_0_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_7_0_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_7_0_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_7_0_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_7_0_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_7_0_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_7_0_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_7_0_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_7_0_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_7_0_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_8_0_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_8_0_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_8_0_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_8_0_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_8_0_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_8_0_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_8_0_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_8_0_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_8_0_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_9_0_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_9_0_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_9_0_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_9_0_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_9_0_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_9_0_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_9_0_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_9_0_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_9_0_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_10_0_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_10_0_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_10_0_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_10_0_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_10_0_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_10_0_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_10_0_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_10_0_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_10_0_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_11_0_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_11_0_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_11_0_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_11_0_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_11_0_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_11_0_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_11_0_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_11_0_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_11_0_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_12_0_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_12_0_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_12_0_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_12_0_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_12_0_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_12_0_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_12_0_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_12_0_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_12_0_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_13_0_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_13_0_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_13_0_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_13_0_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_13_0_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_13_0_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_13_0_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_13_0_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_13_0_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_14_0_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_14_0_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_14_0_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_14_0_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_14_0_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_14_0_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_14_0_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_14_0_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_14_0_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_15_0_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_15_0_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_15_0_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_15_0_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_15_0_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_15_0_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_I_15_0_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_I_15_0_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_I_15_0_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_0_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_0_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_0_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_0_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_0_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_0_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_0_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_0_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_0_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_1_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_1_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_1_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_1_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_1_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_1_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_1_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_1_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_1_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_2_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_2_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_2_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_2_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_2_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_2_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_2_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_2_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_2_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_3_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_3_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_3_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_3_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_3_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_3_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_3_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_3_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_3_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_4_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_4_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_4_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_4_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_4_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_4_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_4_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_4_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_4_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_5_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_5_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_5_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_5_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_5_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_5_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_5_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_5_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_5_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_6_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_6_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_6_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_6_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_6_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_6_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_6_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_6_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_6_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_7_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_7_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_7_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_7_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_7_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_7_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_7_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_7_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_7_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_8_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_8_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_8_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_8_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_8_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_8_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_8_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_8_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_8_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_9_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_9_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_9_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_9_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_9_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_9_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_9_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_9_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_9_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_10_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_10_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_10_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_10_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_10_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_10_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_10_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_10_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_10_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_11_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_11_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_11_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_11_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_11_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_11_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_11_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_11_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_11_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_12_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_12_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_12_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_12_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_12_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_12_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_12_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_12_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_12_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_13_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_13_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_13_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_13_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_13_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_13_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_13_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_13_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_13_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_14_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_14_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_14_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_14_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_14_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_14_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_14_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_14_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_14_2_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_15_0_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_15_0_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_15_0_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_15_1_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_15_1_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_15_1_2; // @[Top.scala 196:21]
  wire [7:0] n65_O_15_2_0; // @[Top.scala 196:21]
  wire [7:0] n65_O_15_2_1; // @[Top.scala 196:21]
  wire [7:0] n65_O_15_2_2; // @[Top.scala 196:21]
  wire  n105_clock; // @[Top.scala 199:22]
  wire  n105_reset; // @[Top.scala 199:22]
  wire  n105_valid_up; // @[Top.scala 199:22]
  wire  n105_valid_down; // @[Top.scala 199:22]
  wire [7:0] n105_I_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_0_0_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_0_0_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_0_1_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_0_1_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_0_1_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_0_2_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_0_2_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_0_2_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_1_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_1_0_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_1_0_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_1_1_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_1_1_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_1_1_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_1_2_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_1_2_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_1_2_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_2_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_2_0_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_2_0_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_2_1_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_2_1_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_2_1_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_2_2_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_2_2_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_2_2_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_3_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_3_0_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_3_0_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_3_1_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_3_1_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_3_1_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_3_2_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_3_2_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_3_2_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_4_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_4_0_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_4_0_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_4_1_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_4_1_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_4_1_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_4_2_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_4_2_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_4_2_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_5_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_5_0_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_5_0_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_5_1_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_5_1_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_5_1_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_5_2_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_5_2_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_5_2_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_6_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_6_0_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_6_0_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_6_1_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_6_1_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_6_1_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_6_2_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_6_2_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_6_2_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_7_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_7_0_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_7_0_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_7_1_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_7_1_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_7_1_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_7_2_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_7_2_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_7_2_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_8_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_8_0_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_8_0_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_8_1_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_8_1_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_8_1_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_8_2_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_8_2_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_8_2_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_9_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_9_0_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_9_0_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_9_1_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_9_1_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_9_1_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_9_2_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_9_2_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_9_2_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_10_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_10_0_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_10_0_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_10_1_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_10_1_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_10_1_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_10_2_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_10_2_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_10_2_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_11_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_11_0_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_11_0_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_11_1_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_11_1_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_11_1_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_11_2_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_11_2_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_11_2_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_12_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_12_0_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_12_0_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_12_1_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_12_1_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_12_1_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_12_2_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_12_2_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_12_2_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_13_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_13_0_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_13_0_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_13_1_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_13_1_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_13_1_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_13_2_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_13_2_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_13_2_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_14_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_14_0_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_14_0_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_14_1_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_14_1_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_14_1_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_14_2_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_14_2_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_14_2_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_15_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_15_0_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_15_0_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_15_1_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_15_1_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_15_1_2; // @[Top.scala 199:22]
  wire [7:0] n105_I_15_2_0; // @[Top.scala 199:22]
  wire [7:0] n105_I_15_2_1; // @[Top.scala 199:22]
  wire [7:0] n105_I_15_2_2; // @[Top.scala 199:22]
  wire [7:0] n105_O_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_O_1_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_O_2_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_O_3_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_O_4_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_O_5_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_O_6_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_O_7_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_O_8_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_O_9_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_O_10_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_O_11_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_O_12_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_O_13_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_O_14_0_0; // @[Top.scala 199:22]
  wire [7:0] n105_O_15_0_0; // @[Top.scala 199:22]
  wire  n106_valid_up; // @[Top.scala 202:22]
  wire  n106_valid_down; // @[Top.scala 202:22]
  wire [7:0] n106_I_0_0_0; // @[Top.scala 202:22]
  wire [7:0] n106_I_1_0_0; // @[Top.scala 202:22]
  wire [7:0] n106_I_2_0_0; // @[Top.scala 202:22]
  wire [7:0] n106_I_3_0_0; // @[Top.scala 202:22]
  wire [7:0] n106_I_4_0_0; // @[Top.scala 202:22]
  wire [7:0] n106_I_5_0_0; // @[Top.scala 202:22]
  wire [7:0] n106_I_6_0_0; // @[Top.scala 202:22]
  wire [7:0] n106_I_7_0_0; // @[Top.scala 202:22]
  wire [7:0] n106_I_8_0_0; // @[Top.scala 202:22]
  wire [7:0] n106_I_9_0_0; // @[Top.scala 202:22]
  wire [7:0] n106_I_10_0_0; // @[Top.scala 202:22]
  wire [7:0] n106_I_11_0_0; // @[Top.scala 202:22]
  wire [7:0] n106_I_12_0_0; // @[Top.scala 202:22]
  wire [7:0] n106_I_13_0_0; // @[Top.scala 202:22]
  wire [7:0] n106_I_14_0_0; // @[Top.scala 202:22]
  wire [7:0] n106_I_15_0_0; // @[Top.scala 202:22]
  wire [7:0] n106_O_0_0; // @[Top.scala 202:22]
  wire [7:0] n106_O_1_0; // @[Top.scala 202:22]
  wire [7:0] n106_O_2_0; // @[Top.scala 202:22]
  wire [7:0] n106_O_3_0; // @[Top.scala 202:22]
  wire [7:0] n106_O_4_0; // @[Top.scala 202:22]
  wire [7:0] n106_O_5_0; // @[Top.scala 202:22]
  wire [7:0] n106_O_6_0; // @[Top.scala 202:22]
  wire [7:0] n106_O_7_0; // @[Top.scala 202:22]
  wire [7:0] n106_O_8_0; // @[Top.scala 202:22]
  wire [7:0] n106_O_9_0; // @[Top.scala 202:22]
  wire [7:0] n106_O_10_0; // @[Top.scala 202:22]
  wire [7:0] n106_O_11_0; // @[Top.scala 202:22]
  wire [7:0] n106_O_12_0; // @[Top.scala 202:22]
  wire [7:0] n106_O_13_0; // @[Top.scala 202:22]
  wire [7:0] n106_O_14_0; // @[Top.scala 202:22]
  wire [7:0] n106_O_15_0; // @[Top.scala 202:22]
  wire  n107_valid_up; // @[Top.scala 205:22]
  wire  n107_valid_down; // @[Top.scala 205:22]
  wire [7:0] n107_I_0_0; // @[Top.scala 205:22]
  wire [7:0] n107_I_1_0; // @[Top.scala 205:22]
  wire [7:0] n107_I_2_0; // @[Top.scala 205:22]
  wire [7:0] n107_I_3_0; // @[Top.scala 205:22]
  wire [7:0] n107_I_4_0; // @[Top.scala 205:22]
  wire [7:0] n107_I_5_0; // @[Top.scala 205:22]
  wire [7:0] n107_I_6_0; // @[Top.scala 205:22]
  wire [7:0] n107_I_7_0; // @[Top.scala 205:22]
  wire [7:0] n107_I_8_0; // @[Top.scala 205:22]
  wire [7:0] n107_I_9_0; // @[Top.scala 205:22]
  wire [7:0] n107_I_10_0; // @[Top.scala 205:22]
  wire [7:0] n107_I_11_0; // @[Top.scala 205:22]
  wire [7:0] n107_I_12_0; // @[Top.scala 205:22]
  wire [7:0] n107_I_13_0; // @[Top.scala 205:22]
  wire [7:0] n107_I_14_0; // @[Top.scala 205:22]
  wire [7:0] n107_I_15_0; // @[Top.scala 205:22]
  wire [7:0] n107_O_0; // @[Top.scala 205:22]
  wire [7:0] n107_O_1; // @[Top.scala 205:22]
  wire [7:0] n107_O_2; // @[Top.scala 205:22]
  wire [7:0] n107_O_3; // @[Top.scala 205:22]
  wire [7:0] n107_O_4; // @[Top.scala 205:22]
  wire [7:0] n107_O_5; // @[Top.scala 205:22]
  wire [7:0] n107_O_6; // @[Top.scala 205:22]
  wire [7:0] n107_O_7; // @[Top.scala 205:22]
  wire [7:0] n107_O_8; // @[Top.scala 205:22]
  wire [7:0] n107_O_9; // @[Top.scala 205:22]
  wire [7:0] n107_O_10; // @[Top.scala 205:22]
  wire [7:0] n107_O_11; // @[Top.scala 205:22]
  wire [7:0] n107_O_12; // @[Top.scala 205:22]
  wire [7:0] n107_O_13; // @[Top.scala 205:22]
  wire [7:0] n107_O_14; // @[Top.scala 205:22]
  wire [7:0] n107_O_15; // @[Top.scala 205:22]
  wire  n108_clock; // @[Top.scala 208:22]
  wire  n108_reset; // @[Top.scala 208:22]
  wire  n108_valid_up; // @[Top.scala 208:22]
  wire  n108_valid_down; // @[Top.scala 208:22]
  wire [7:0] n108_I_0; // @[Top.scala 208:22]
  wire [7:0] n108_I_1; // @[Top.scala 208:22]
  wire [7:0] n108_I_2; // @[Top.scala 208:22]
  wire [7:0] n108_I_3; // @[Top.scala 208:22]
  wire [7:0] n108_I_4; // @[Top.scala 208:22]
  wire [7:0] n108_I_5; // @[Top.scala 208:22]
  wire [7:0] n108_I_6; // @[Top.scala 208:22]
  wire [7:0] n108_I_7; // @[Top.scala 208:22]
  wire [7:0] n108_I_8; // @[Top.scala 208:22]
  wire [7:0] n108_I_9; // @[Top.scala 208:22]
  wire [7:0] n108_I_10; // @[Top.scala 208:22]
  wire [7:0] n108_I_11; // @[Top.scala 208:22]
  wire [7:0] n108_I_12; // @[Top.scala 208:22]
  wire [7:0] n108_I_13; // @[Top.scala 208:22]
  wire [7:0] n108_I_14; // @[Top.scala 208:22]
  wire [7:0] n108_I_15; // @[Top.scala 208:22]
  wire [7:0] n108_O_0; // @[Top.scala 208:22]
  wire [7:0] n108_O_1; // @[Top.scala 208:22]
  wire [7:0] n108_O_2; // @[Top.scala 208:22]
  wire [7:0] n108_O_3; // @[Top.scala 208:22]
  wire [7:0] n108_O_4; // @[Top.scala 208:22]
  wire [7:0] n108_O_5; // @[Top.scala 208:22]
  wire [7:0] n108_O_6; // @[Top.scala 208:22]
  wire [7:0] n108_O_7; // @[Top.scala 208:22]
  wire [7:0] n108_O_8; // @[Top.scala 208:22]
  wire [7:0] n108_O_9; // @[Top.scala 208:22]
  wire [7:0] n108_O_10; // @[Top.scala 208:22]
  wire [7:0] n108_O_11; // @[Top.scala 208:22]
  wire [7:0] n108_O_12; // @[Top.scala 208:22]
  wire [7:0] n108_O_13; // @[Top.scala 208:22]
  wire [7:0] n108_O_14; // @[Top.scala 208:22]
  wire [7:0] n108_O_15; // @[Top.scala 208:22]
  wire  n109_clock; // @[Top.scala 211:22]
  wire  n109_reset; // @[Top.scala 211:22]
  wire  n109_valid_up; // @[Top.scala 211:22]
  wire  n109_valid_down; // @[Top.scala 211:22]
  wire [7:0] n109_I0_0; // @[Top.scala 211:22]
  wire [7:0] n109_I0_1; // @[Top.scala 211:22]
  wire [7:0] n109_I0_2; // @[Top.scala 211:22]
  wire [7:0] n109_I0_3; // @[Top.scala 211:22]
  wire [7:0] n109_I0_4; // @[Top.scala 211:22]
  wire [7:0] n109_I0_5; // @[Top.scala 211:22]
  wire [7:0] n109_I0_6; // @[Top.scala 211:22]
  wire [7:0] n109_I0_7; // @[Top.scala 211:22]
  wire [7:0] n109_I0_8; // @[Top.scala 211:22]
  wire [7:0] n109_I0_9; // @[Top.scala 211:22]
  wire [7:0] n109_I0_10; // @[Top.scala 211:22]
  wire [7:0] n109_I0_11; // @[Top.scala 211:22]
  wire [7:0] n109_I0_12; // @[Top.scala 211:22]
  wire [7:0] n109_I0_13; // @[Top.scala 211:22]
  wire [7:0] n109_I0_14; // @[Top.scala 211:22]
  wire [7:0] n109_I0_15; // @[Top.scala 211:22]
  wire [7:0] n109_I1_0; // @[Top.scala 211:22]
  wire [7:0] n109_I1_1; // @[Top.scala 211:22]
  wire [7:0] n109_I1_2; // @[Top.scala 211:22]
  wire [7:0] n109_I1_3; // @[Top.scala 211:22]
  wire [7:0] n109_I1_4; // @[Top.scala 211:22]
  wire [7:0] n109_I1_5; // @[Top.scala 211:22]
  wire [7:0] n109_I1_6; // @[Top.scala 211:22]
  wire [7:0] n109_I1_7; // @[Top.scala 211:22]
  wire [7:0] n109_I1_8; // @[Top.scala 211:22]
  wire [7:0] n109_I1_9; // @[Top.scala 211:22]
  wire [7:0] n109_I1_10; // @[Top.scala 211:22]
  wire [7:0] n109_I1_11; // @[Top.scala 211:22]
  wire [7:0] n109_I1_12; // @[Top.scala 211:22]
  wire [7:0] n109_I1_13; // @[Top.scala 211:22]
  wire [7:0] n109_I1_14; // @[Top.scala 211:22]
  wire [7:0] n109_I1_15; // @[Top.scala 211:22]
  wire [7:0] n109_O_0; // @[Top.scala 211:22]
  wire [7:0] n109_O_1; // @[Top.scala 211:22]
  wire [7:0] n109_O_2; // @[Top.scala 211:22]
  wire [7:0] n109_O_3; // @[Top.scala 211:22]
  wire [7:0] n109_O_4; // @[Top.scala 211:22]
  wire [7:0] n109_O_5; // @[Top.scala 211:22]
  wire [7:0] n109_O_6; // @[Top.scala 211:22]
  wire [7:0] n109_O_7; // @[Top.scala 211:22]
  wire [7:0] n109_O_8; // @[Top.scala 211:22]
  wire [7:0] n109_O_9; // @[Top.scala 211:22]
  wire [7:0] n109_O_10; // @[Top.scala 211:22]
  wire [7:0] n109_O_11; // @[Top.scala 211:22]
  wire [7:0] n109_O_12; // @[Top.scala 211:22]
  wire [7:0] n109_O_13; // @[Top.scala 211:22]
  wire [7:0] n109_O_14; // @[Top.scala 211:22]
  wire [7:0] n109_O_15; // @[Top.scala 211:22]
  wire  n136_clock; // @[Top.scala 215:22]
  wire  n136_reset; // @[Top.scala 215:22]
  wire  n136_valid_up; // @[Top.scala 215:22]
  wire  n136_valid_down; // @[Top.scala 215:22]
  wire [7:0] n136_I_0; // @[Top.scala 215:22]
  wire [7:0] n136_I_1; // @[Top.scala 215:22]
  wire [7:0] n136_I_2; // @[Top.scala 215:22]
  wire [7:0] n136_I_3; // @[Top.scala 215:22]
  wire [7:0] n136_I_4; // @[Top.scala 215:22]
  wire [7:0] n136_I_5; // @[Top.scala 215:22]
  wire [7:0] n136_I_6; // @[Top.scala 215:22]
  wire [7:0] n136_I_7; // @[Top.scala 215:22]
  wire [7:0] n136_I_8; // @[Top.scala 215:22]
  wire [7:0] n136_I_9; // @[Top.scala 215:22]
  wire [7:0] n136_I_10; // @[Top.scala 215:22]
  wire [7:0] n136_I_11; // @[Top.scala 215:22]
  wire [7:0] n136_I_12; // @[Top.scala 215:22]
  wire [7:0] n136_I_13; // @[Top.scala 215:22]
  wire [7:0] n136_I_14; // @[Top.scala 215:22]
  wire [7:0] n136_I_15; // @[Top.scala 215:22]
  wire [7:0] n136_O_0; // @[Top.scala 215:22]
  wire [7:0] n136_O_1; // @[Top.scala 215:22]
  wire [7:0] n136_O_2; // @[Top.scala 215:22]
  wire [7:0] n136_O_3; // @[Top.scala 215:22]
  wire [7:0] n136_O_4; // @[Top.scala 215:22]
  wire [7:0] n136_O_5; // @[Top.scala 215:22]
  wire [7:0] n136_O_6; // @[Top.scala 215:22]
  wire [7:0] n136_O_7; // @[Top.scala 215:22]
  wire [7:0] n136_O_8; // @[Top.scala 215:22]
  wire [7:0] n136_O_9; // @[Top.scala 215:22]
  wire [7:0] n136_O_10; // @[Top.scala 215:22]
  wire [7:0] n136_O_11; // @[Top.scala 215:22]
  wire [7:0] n136_O_12; // @[Top.scala 215:22]
  wire [7:0] n136_O_13; // @[Top.scala 215:22]
  wire [7:0] n136_O_14; // @[Top.scala 215:22]
  wire [7:0] n136_O_15; // @[Top.scala 215:22]
  wire  n137_clock; // @[Top.scala 218:22]
  wire  n137_reset; // @[Top.scala 218:22]
  wire  n137_valid_up; // @[Top.scala 218:22]
  wire  n137_valid_down; // @[Top.scala 218:22]
  wire [7:0] n137_I_0; // @[Top.scala 218:22]
  wire [7:0] n137_I_1; // @[Top.scala 218:22]
  wire [7:0] n137_I_2; // @[Top.scala 218:22]
  wire [7:0] n137_I_3; // @[Top.scala 218:22]
  wire [7:0] n137_I_4; // @[Top.scala 218:22]
  wire [7:0] n137_I_5; // @[Top.scala 218:22]
  wire [7:0] n137_I_6; // @[Top.scala 218:22]
  wire [7:0] n137_I_7; // @[Top.scala 218:22]
  wire [7:0] n137_I_8; // @[Top.scala 218:22]
  wire [7:0] n137_I_9; // @[Top.scala 218:22]
  wire [7:0] n137_I_10; // @[Top.scala 218:22]
  wire [7:0] n137_I_11; // @[Top.scala 218:22]
  wire [7:0] n137_I_12; // @[Top.scala 218:22]
  wire [7:0] n137_I_13; // @[Top.scala 218:22]
  wire [7:0] n137_I_14; // @[Top.scala 218:22]
  wire [7:0] n137_I_15; // @[Top.scala 218:22]
  wire [7:0] n137_O_0; // @[Top.scala 218:22]
  wire [7:0] n137_O_1; // @[Top.scala 218:22]
  wire [7:0] n137_O_2; // @[Top.scala 218:22]
  wire [7:0] n137_O_3; // @[Top.scala 218:22]
  wire [7:0] n137_O_4; // @[Top.scala 218:22]
  wire [7:0] n137_O_5; // @[Top.scala 218:22]
  wire [7:0] n137_O_6; // @[Top.scala 218:22]
  wire [7:0] n137_O_7; // @[Top.scala 218:22]
  wire [7:0] n137_O_8; // @[Top.scala 218:22]
  wire [7:0] n137_O_9; // @[Top.scala 218:22]
  wire [7:0] n137_O_10; // @[Top.scala 218:22]
  wire [7:0] n137_O_11; // @[Top.scala 218:22]
  wire [7:0] n137_O_12; // @[Top.scala 218:22]
  wire [7:0] n137_O_13; // @[Top.scala 218:22]
  wire [7:0] n137_O_14; // @[Top.scala 218:22]
  wire [7:0] n137_O_15; // @[Top.scala 218:22]
  wire  n138_clock; // @[Top.scala 221:22]
  wire  n138_reset; // @[Top.scala 221:22]
  wire  n138_valid_up; // @[Top.scala 221:22]
  wire  n138_valid_down; // @[Top.scala 221:22]
  wire [7:0] n138_I_0; // @[Top.scala 221:22]
  wire [7:0] n138_I_1; // @[Top.scala 221:22]
  wire [7:0] n138_I_2; // @[Top.scala 221:22]
  wire [7:0] n138_I_3; // @[Top.scala 221:22]
  wire [7:0] n138_I_4; // @[Top.scala 221:22]
  wire [7:0] n138_I_5; // @[Top.scala 221:22]
  wire [7:0] n138_I_6; // @[Top.scala 221:22]
  wire [7:0] n138_I_7; // @[Top.scala 221:22]
  wire [7:0] n138_I_8; // @[Top.scala 221:22]
  wire [7:0] n138_I_9; // @[Top.scala 221:22]
  wire [7:0] n138_I_10; // @[Top.scala 221:22]
  wire [7:0] n138_I_11; // @[Top.scala 221:22]
  wire [7:0] n138_I_12; // @[Top.scala 221:22]
  wire [7:0] n138_I_13; // @[Top.scala 221:22]
  wire [7:0] n138_I_14; // @[Top.scala 221:22]
  wire [7:0] n138_I_15; // @[Top.scala 221:22]
  wire [7:0] n138_O_0; // @[Top.scala 221:22]
  wire [7:0] n138_O_1; // @[Top.scala 221:22]
  wire [7:0] n138_O_2; // @[Top.scala 221:22]
  wire [7:0] n138_O_3; // @[Top.scala 221:22]
  wire [7:0] n138_O_4; // @[Top.scala 221:22]
  wire [7:0] n138_O_5; // @[Top.scala 221:22]
  wire [7:0] n138_O_6; // @[Top.scala 221:22]
  wire [7:0] n138_O_7; // @[Top.scala 221:22]
  wire [7:0] n138_O_8; // @[Top.scala 221:22]
  wire [7:0] n138_O_9; // @[Top.scala 221:22]
  wire [7:0] n138_O_10; // @[Top.scala 221:22]
  wire [7:0] n138_O_11; // @[Top.scala 221:22]
  wire [7:0] n138_O_12; // @[Top.scala 221:22]
  wire [7:0] n138_O_13; // @[Top.scala 221:22]
  wire [7:0] n138_O_14; // @[Top.scala 221:22]
  wire [7:0] n138_O_15; // @[Top.scala 221:22]
  FIFO n1 ( // @[Top.scala 116:20]
    .clock(n1_clock),
    .reset(n1_reset),
    .valid_up(n1_valid_up),
    .valid_down(n1_valid_down),
    .I_0(n1_I_0),
    .I_1(n1_I_1),
    .I_2(n1_I_2),
    .I_3(n1_I_3),
    .I_4(n1_I_4),
    .I_5(n1_I_5),
    .I_6(n1_I_6),
    .I_7(n1_I_7),
    .I_8(n1_I_8),
    .I_9(n1_I_9),
    .I_10(n1_I_10),
    .I_11(n1_I_11),
    .I_12(n1_I_12),
    .I_13(n1_I_13),
    .I_14(n1_I_14),
    .I_15(n1_I_15),
    .O_0(n1_O_0),
    .O_1(n1_O_1),
    .O_2(n1_O_2),
    .O_3(n1_O_3),
    .O_4(n1_O_4),
    .O_5(n1_O_5),
    .O_6(n1_O_6),
    .O_7(n1_O_7),
    .O_8(n1_O_8),
    .O_9(n1_O_9),
    .O_10(n1_O_10),
    .O_11(n1_O_11),
    .O_12(n1_O_12),
    .O_13(n1_O_13),
    .O_14(n1_O_14),
    .O_15(n1_O_15)
  );
  ShiftS n2 ( // @[Top.scala 119:20]
    .valid_up(n2_valid_up),
    .valid_down(n2_valid_down),
    .I_0(n2_I_0),
    .I_1(n2_I_1),
    .I_2(n2_I_2),
    .I_3(n2_I_3),
    .I_4(n2_I_4),
    .I_5(n2_I_5),
    .I_6(n2_I_6),
    .I_7(n2_I_7),
    .I_8(n2_I_8),
    .I_9(n2_I_9),
    .I_10(n2_I_10),
    .I_11(n2_I_11),
    .I_12(n2_I_12),
    .I_13(n2_I_13),
    .I_14(n2_I_14),
    .I_15(n2_I_15),
    .O_0(n2_O_0),
    .O_1(n2_O_1),
    .O_2(n2_O_2),
    .O_3(n2_O_3),
    .O_4(n2_O_4),
    .O_5(n2_O_5),
    .O_6(n2_O_6),
    .O_7(n2_O_7),
    .O_8(n2_O_8),
    .O_9(n2_O_9),
    .O_10(n2_O_10),
    .O_11(n2_O_11),
    .O_12(n2_O_12),
    .O_13(n2_O_13),
    .O_14(n2_O_14),
    .O_15(n2_O_15)
  );
  ShiftS n3 ( // @[Top.scala 122:20]
    .valid_up(n3_valid_up),
    .valid_down(n3_valid_down),
    .I_0(n3_I_0),
    .I_1(n3_I_1),
    .I_2(n3_I_2),
    .I_3(n3_I_3),
    .I_4(n3_I_4),
    .I_5(n3_I_5),
    .I_6(n3_I_6),
    .I_7(n3_I_7),
    .I_8(n3_I_8),
    .I_9(n3_I_9),
    .I_10(n3_I_10),
    .I_11(n3_I_11),
    .I_12(n3_I_12),
    .I_13(n3_I_13),
    .I_14(n3_I_14),
    .I_15(n3_I_15),
    .O_0(n3_O_0),
    .O_1(n3_O_1),
    .O_2(n3_O_2),
    .O_3(n3_O_3),
    .O_4(n3_O_4),
    .O_5(n3_O_5),
    .O_6(n3_O_6),
    .O_7(n3_O_7),
    .O_8(n3_O_8),
    .O_9(n3_O_9),
    .O_10(n3_O_10),
    .O_11(n3_O_11),
    .O_12(n3_O_12),
    .O_13(n3_O_13),
    .O_14(n3_O_14),
    .O_15(n3_O_15)
  );
  ShiftS_2 n4 ( // @[Top.scala 125:20]
    .valid_up(n4_valid_up),
    .valid_down(n4_valid_down),
    .I_0(n4_I_0),
    .I_1(n4_I_1),
    .I_2(n4_I_2),
    .I_3(n4_I_3),
    .I_4(n4_I_4),
    .I_5(n4_I_5),
    .I_6(n4_I_6),
    .I_7(n4_I_7),
    .I_8(n4_I_8),
    .I_9(n4_I_9),
    .I_10(n4_I_10),
    .I_11(n4_I_11),
    .I_12(n4_I_12),
    .I_13(n4_I_13),
    .I_14(n4_I_14),
    .I_15(n4_I_15),
    .O_0(n4_O_0),
    .O_1(n4_O_1),
    .O_2(n4_O_2),
    .O_3(n4_O_3),
    .O_4(n4_O_4),
    .O_5(n4_O_5),
    .O_6(n4_O_6),
    .O_7(n4_O_7),
    .O_8(n4_O_8),
    .O_9(n4_O_9),
    .O_10(n4_O_10),
    .O_11(n4_O_11),
    .O_12(n4_O_12),
    .O_13(n4_O_13),
    .O_14(n4_O_14),
    .O_15(n4_O_15)
  );
  ShiftS_2 n5 ( // @[Top.scala 128:20]
    .valid_up(n5_valid_up),
    .valid_down(n5_valid_down),
    .I_0(n5_I_0),
    .I_1(n5_I_1),
    .I_2(n5_I_2),
    .I_3(n5_I_3),
    .I_4(n5_I_4),
    .I_5(n5_I_5),
    .I_6(n5_I_6),
    .I_7(n5_I_7),
    .I_8(n5_I_8),
    .I_9(n5_I_9),
    .I_10(n5_I_10),
    .I_11(n5_I_11),
    .I_12(n5_I_12),
    .I_13(n5_I_13),
    .I_14(n5_I_14),
    .I_15(n5_I_15),
    .O_0(n5_O_0),
    .O_1(n5_O_1),
    .O_2(n5_O_2),
    .O_3(n5_O_3),
    .O_4(n5_O_4),
    .O_5(n5_O_5),
    .O_6(n5_O_6),
    .O_7(n5_O_7),
    .O_8(n5_O_8),
    .O_9(n5_O_9),
    .O_10(n5_O_10),
    .O_11(n5_O_11),
    .O_12(n5_O_12),
    .O_13(n5_O_13),
    .O_14(n5_O_14),
    .O_15(n5_O_15)
  );
  Map2S n6 ( // @[Top.scala 131:20]
    .valid_up(n6_valid_up),
    .valid_down(n6_valid_down),
    .I0_0(n6_I0_0),
    .I0_1(n6_I0_1),
    .I0_2(n6_I0_2),
    .I0_3(n6_I0_3),
    .I0_4(n6_I0_4),
    .I0_5(n6_I0_5),
    .I0_6(n6_I0_6),
    .I0_7(n6_I0_7),
    .I0_8(n6_I0_8),
    .I0_9(n6_I0_9),
    .I0_10(n6_I0_10),
    .I0_11(n6_I0_11),
    .I0_12(n6_I0_12),
    .I0_13(n6_I0_13),
    .I0_14(n6_I0_14),
    .I0_15(n6_I0_15),
    .I1_0(n6_I1_0),
    .I1_1(n6_I1_1),
    .I1_2(n6_I1_2),
    .I1_3(n6_I1_3),
    .I1_4(n6_I1_4),
    .I1_5(n6_I1_5),
    .I1_6(n6_I1_6),
    .I1_7(n6_I1_7),
    .I1_8(n6_I1_8),
    .I1_9(n6_I1_9),
    .I1_10(n6_I1_10),
    .I1_11(n6_I1_11),
    .I1_12(n6_I1_12),
    .I1_13(n6_I1_13),
    .I1_14(n6_I1_14),
    .I1_15(n6_I1_15),
    .O_0_0(n6_O_0_0),
    .O_0_1(n6_O_0_1),
    .O_1_0(n6_O_1_0),
    .O_1_1(n6_O_1_1),
    .O_2_0(n6_O_2_0),
    .O_2_1(n6_O_2_1),
    .O_3_0(n6_O_3_0),
    .O_3_1(n6_O_3_1),
    .O_4_0(n6_O_4_0),
    .O_4_1(n6_O_4_1),
    .O_5_0(n6_O_5_0),
    .O_5_1(n6_O_5_1),
    .O_6_0(n6_O_6_0),
    .O_6_1(n6_O_6_1),
    .O_7_0(n6_O_7_0),
    .O_7_1(n6_O_7_1),
    .O_8_0(n6_O_8_0),
    .O_8_1(n6_O_8_1),
    .O_9_0(n6_O_9_0),
    .O_9_1(n6_O_9_1),
    .O_10_0(n6_O_10_0),
    .O_10_1(n6_O_10_1),
    .O_11_0(n6_O_11_0),
    .O_11_1(n6_O_11_1),
    .O_12_0(n6_O_12_0),
    .O_12_1(n6_O_12_1),
    .O_13_0(n6_O_13_0),
    .O_13_1(n6_O_13_1),
    .O_14_0(n6_O_14_0),
    .O_14_1(n6_O_14_1),
    .O_15_0(n6_O_15_0),
    .O_15_1(n6_O_15_1)
  );
  Map2S_1 n10 ( // @[Top.scala 135:21]
    .valid_up(n10_valid_up),
    .valid_down(n10_valid_down),
    .I0_0_0(n10_I0_0_0),
    .I0_0_1(n10_I0_0_1),
    .I0_1_0(n10_I0_1_0),
    .I0_1_1(n10_I0_1_1),
    .I0_2_0(n10_I0_2_0),
    .I0_2_1(n10_I0_2_1),
    .I0_3_0(n10_I0_3_0),
    .I0_3_1(n10_I0_3_1),
    .I0_4_0(n10_I0_4_0),
    .I0_4_1(n10_I0_4_1),
    .I0_5_0(n10_I0_5_0),
    .I0_5_1(n10_I0_5_1),
    .I0_6_0(n10_I0_6_0),
    .I0_6_1(n10_I0_6_1),
    .I0_7_0(n10_I0_7_0),
    .I0_7_1(n10_I0_7_1),
    .I0_8_0(n10_I0_8_0),
    .I0_8_1(n10_I0_8_1),
    .I0_9_0(n10_I0_9_0),
    .I0_9_1(n10_I0_9_1),
    .I0_10_0(n10_I0_10_0),
    .I0_10_1(n10_I0_10_1),
    .I0_11_0(n10_I0_11_0),
    .I0_11_1(n10_I0_11_1),
    .I0_12_0(n10_I0_12_0),
    .I0_12_1(n10_I0_12_1),
    .I0_13_0(n10_I0_13_0),
    .I0_13_1(n10_I0_13_1),
    .I0_14_0(n10_I0_14_0),
    .I0_14_1(n10_I0_14_1),
    .I0_15_0(n10_I0_15_0),
    .I0_15_1(n10_I0_15_1),
    .I1_0(n10_I1_0),
    .I1_1(n10_I1_1),
    .I1_2(n10_I1_2),
    .I1_3(n10_I1_3),
    .I1_4(n10_I1_4),
    .I1_5(n10_I1_5),
    .I1_6(n10_I1_6),
    .I1_7(n10_I1_7),
    .I1_8(n10_I1_8),
    .I1_9(n10_I1_9),
    .I1_10(n10_I1_10),
    .I1_11(n10_I1_11),
    .I1_12(n10_I1_12),
    .I1_13(n10_I1_13),
    .I1_14(n10_I1_14),
    .I1_15(n10_I1_15),
    .O_0_0(n10_O_0_0),
    .O_0_1(n10_O_0_1),
    .O_0_2(n10_O_0_2),
    .O_1_0(n10_O_1_0),
    .O_1_1(n10_O_1_1),
    .O_1_2(n10_O_1_2),
    .O_2_0(n10_O_2_0),
    .O_2_1(n10_O_2_1),
    .O_2_2(n10_O_2_2),
    .O_3_0(n10_O_3_0),
    .O_3_1(n10_O_3_1),
    .O_3_2(n10_O_3_2),
    .O_4_0(n10_O_4_0),
    .O_4_1(n10_O_4_1),
    .O_4_2(n10_O_4_2),
    .O_5_0(n10_O_5_0),
    .O_5_1(n10_O_5_1),
    .O_5_2(n10_O_5_2),
    .O_6_0(n10_O_6_0),
    .O_6_1(n10_O_6_1),
    .O_6_2(n10_O_6_2),
    .O_7_0(n10_O_7_0),
    .O_7_1(n10_O_7_1),
    .O_7_2(n10_O_7_2),
    .O_8_0(n10_O_8_0),
    .O_8_1(n10_O_8_1),
    .O_8_2(n10_O_8_2),
    .O_9_0(n10_O_9_0),
    .O_9_1(n10_O_9_1),
    .O_9_2(n10_O_9_2),
    .O_10_0(n10_O_10_0),
    .O_10_1(n10_O_10_1),
    .O_10_2(n10_O_10_2),
    .O_11_0(n10_O_11_0),
    .O_11_1(n10_O_11_1),
    .O_11_2(n10_O_11_2),
    .O_12_0(n10_O_12_0),
    .O_12_1(n10_O_12_1),
    .O_12_2(n10_O_12_2),
    .O_13_0(n10_O_13_0),
    .O_13_1(n10_O_13_1),
    .O_13_2(n10_O_13_2),
    .O_14_0(n10_O_14_0),
    .O_14_1(n10_O_14_1),
    .O_14_2(n10_O_14_2),
    .O_15_0(n10_O_15_0),
    .O_15_1(n10_O_15_1),
    .O_15_2(n10_O_15_2)
  );
  PartitionS n14 ( // @[Top.scala 139:21]
    .valid_up(n14_valid_up),
    .valid_down(n14_valid_down),
    .I_0_0(n14_I_0_0),
    .I_0_1(n14_I_0_1),
    .I_0_2(n14_I_0_2),
    .I_1_0(n14_I_1_0),
    .I_1_1(n14_I_1_1),
    .I_1_2(n14_I_1_2),
    .I_2_0(n14_I_2_0),
    .I_2_1(n14_I_2_1),
    .I_2_2(n14_I_2_2),
    .I_3_0(n14_I_3_0),
    .I_3_1(n14_I_3_1),
    .I_3_2(n14_I_3_2),
    .I_4_0(n14_I_4_0),
    .I_4_1(n14_I_4_1),
    .I_4_2(n14_I_4_2),
    .I_5_0(n14_I_5_0),
    .I_5_1(n14_I_5_1),
    .I_5_2(n14_I_5_2),
    .I_6_0(n14_I_6_0),
    .I_6_1(n14_I_6_1),
    .I_6_2(n14_I_6_2),
    .I_7_0(n14_I_7_0),
    .I_7_1(n14_I_7_1),
    .I_7_2(n14_I_7_2),
    .I_8_0(n14_I_8_0),
    .I_8_1(n14_I_8_1),
    .I_8_2(n14_I_8_2),
    .I_9_0(n14_I_9_0),
    .I_9_1(n14_I_9_1),
    .I_9_2(n14_I_9_2),
    .I_10_0(n14_I_10_0),
    .I_10_1(n14_I_10_1),
    .I_10_2(n14_I_10_2),
    .I_11_0(n14_I_11_0),
    .I_11_1(n14_I_11_1),
    .I_11_2(n14_I_11_2),
    .I_12_0(n14_I_12_0),
    .I_12_1(n14_I_12_1),
    .I_12_2(n14_I_12_2),
    .I_13_0(n14_I_13_0),
    .I_13_1(n14_I_13_1),
    .I_13_2(n14_I_13_2),
    .I_14_0(n14_I_14_0),
    .I_14_1(n14_I_14_1),
    .I_14_2(n14_I_14_2),
    .I_15_0(n14_I_15_0),
    .I_15_1(n14_I_15_1),
    .I_15_2(n14_I_15_2),
    .O_0_0_0(n14_O_0_0_0),
    .O_0_0_1(n14_O_0_0_1),
    .O_0_0_2(n14_O_0_0_2),
    .O_1_0_0(n14_O_1_0_0),
    .O_1_0_1(n14_O_1_0_1),
    .O_1_0_2(n14_O_1_0_2),
    .O_2_0_0(n14_O_2_0_0),
    .O_2_0_1(n14_O_2_0_1),
    .O_2_0_2(n14_O_2_0_2),
    .O_3_0_0(n14_O_3_0_0),
    .O_3_0_1(n14_O_3_0_1),
    .O_3_0_2(n14_O_3_0_2),
    .O_4_0_0(n14_O_4_0_0),
    .O_4_0_1(n14_O_4_0_1),
    .O_4_0_2(n14_O_4_0_2),
    .O_5_0_0(n14_O_5_0_0),
    .O_5_0_1(n14_O_5_0_1),
    .O_5_0_2(n14_O_5_0_2),
    .O_6_0_0(n14_O_6_0_0),
    .O_6_0_1(n14_O_6_0_1),
    .O_6_0_2(n14_O_6_0_2),
    .O_7_0_0(n14_O_7_0_0),
    .O_7_0_1(n14_O_7_0_1),
    .O_7_0_2(n14_O_7_0_2),
    .O_8_0_0(n14_O_8_0_0),
    .O_8_0_1(n14_O_8_0_1),
    .O_8_0_2(n14_O_8_0_2),
    .O_9_0_0(n14_O_9_0_0),
    .O_9_0_1(n14_O_9_0_1),
    .O_9_0_2(n14_O_9_0_2),
    .O_10_0_0(n14_O_10_0_0),
    .O_10_0_1(n14_O_10_0_1),
    .O_10_0_2(n14_O_10_0_2),
    .O_11_0_0(n14_O_11_0_0),
    .O_11_0_1(n14_O_11_0_1),
    .O_11_0_2(n14_O_11_0_2),
    .O_12_0_0(n14_O_12_0_0),
    .O_12_0_1(n14_O_12_0_1),
    .O_12_0_2(n14_O_12_0_2),
    .O_13_0_0(n14_O_13_0_0),
    .O_13_0_1(n14_O_13_0_1),
    .O_13_0_2(n14_O_13_0_2),
    .O_14_0_0(n14_O_14_0_0),
    .O_14_0_1(n14_O_14_0_1),
    .O_14_0_2(n14_O_14_0_2),
    .O_15_0_0(n14_O_15_0_0),
    .O_15_0_1(n14_O_15_0_1),
    .O_15_0_2(n14_O_15_0_2)
  );
  MapS n19 ( // @[Top.scala 142:21]
    .valid_up(n19_valid_up),
    .valid_down(n19_valid_down),
    .I_0_0_0(n19_I_0_0_0),
    .I_0_0_1(n19_I_0_0_1),
    .I_0_0_2(n19_I_0_0_2),
    .I_1_0_0(n19_I_1_0_0),
    .I_1_0_1(n19_I_1_0_1),
    .I_1_0_2(n19_I_1_0_2),
    .I_2_0_0(n19_I_2_0_0),
    .I_2_0_1(n19_I_2_0_1),
    .I_2_0_2(n19_I_2_0_2),
    .I_3_0_0(n19_I_3_0_0),
    .I_3_0_1(n19_I_3_0_1),
    .I_3_0_2(n19_I_3_0_2),
    .I_4_0_0(n19_I_4_0_0),
    .I_4_0_1(n19_I_4_0_1),
    .I_4_0_2(n19_I_4_0_2),
    .I_5_0_0(n19_I_5_0_0),
    .I_5_0_1(n19_I_5_0_1),
    .I_5_0_2(n19_I_5_0_2),
    .I_6_0_0(n19_I_6_0_0),
    .I_6_0_1(n19_I_6_0_1),
    .I_6_0_2(n19_I_6_0_2),
    .I_7_0_0(n19_I_7_0_0),
    .I_7_0_1(n19_I_7_0_1),
    .I_7_0_2(n19_I_7_0_2),
    .I_8_0_0(n19_I_8_0_0),
    .I_8_0_1(n19_I_8_0_1),
    .I_8_0_2(n19_I_8_0_2),
    .I_9_0_0(n19_I_9_0_0),
    .I_9_0_1(n19_I_9_0_1),
    .I_9_0_2(n19_I_9_0_2),
    .I_10_0_0(n19_I_10_0_0),
    .I_10_0_1(n19_I_10_0_1),
    .I_10_0_2(n19_I_10_0_2),
    .I_11_0_0(n19_I_11_0_0),
    .I_11_0_1(n19_I_11_0_1),
    .I_11_0_2(n19_I_11_0_2),
    .I_12_0_0(n19_I_12_0_0),
    .I_12_0_1(n19_I_12_0_1),
    .I_12_0_2(n19_I_12_0_2),
    .I_13_0_0(n19_I_13_0_0),
    .I_13_0_1(n19_I_13_0_1),
    .I_13_0_2(n19_I_13_0_2),
    .I_14_0_0(n19_I_14_0_0),
    .I_14_0_1(n19_I_14_0_1),
    .I_14_0_2(n19_I_14_0_2),
    .I_15_0_0(n19_I_15_0_0),
    .I_15_0_1(n19_I_15_0_1),
    .I_15_0_2(n19_I_15_0_2),
    .O_0_0(n19_O_0_0),
    .O_0_1(n19_O_0_1),
    .O_0_2(n19_O_0_2),
    .O_1_0(n19_O_1_0),
    .O_1_1(n19_O_1_1),
    .O_1_2(n19_O_1_2),
    .O_2_0(n19_O_2_0),
    .O_2_1(n19_O_2_1),
    .O_2_2(n19_O_2_2),
    .O_3_0(n19_O_3_0),
    .O_3_1(n19_O_3_1),
    .O_3_2(n19_O_3_2),
    .O_4_0(n19_O_4_0),
    .O_4_1(n19_O_4_1),
    .O_4_2(n19_O_4_2),
    .O_5_0(n19_O_5_0),
    .O_5_1(n19_O_5_1),
    .O_5_2(n19_O_5_2),
    .O_6_0(n19_O_6_0),
    .O_6_1(n19_O_6_1),
    .O_6_2(n19_O_6_2),
    .O_7_0(n19_O_7_0),
    .O_7_1(n19_O_7_1),
    .O_7_2(n19_O_7_2),
    .O_8_0(n19_O_8_0),
    .O_8_1(n19_O_8_1),
    .O_8_2(n19_O_8_2),
    .O_9_0(n19_O_9_0),
    .O_9_1(n19_O_9_1),
    .O_9_2(n19_O_9_2),
    .O_10_0(n19_O_10_0),
    .O_10_1(n19_O_10_1),
    .O_10_2(n19_O_10_2),
    .O_11_0(n19_O_11_0),
    .O_11_1(n19_O_11_1),
    .O_11_2(n19_O_11_2),
    .O_12_0(n19_O_12_0),
    .O_12_1(n19_O_12_1),
    .O_12_2(n19_O_12_2),
    .O_13_0(n19_O_13_0),
    .O_13_1(n19_O_13_1),
    .O_13_2(n19_O_13_2),
    .O_14_0(n19_O_14_0),
    .O_14_1(n19_O_14_1),
    .O_14_2(n19_O_14_2),
    .O_15_0(n19_O_15_0),
    .O_15_1(n19_O_15_1),
    .O_15_2(n19_O_15_2)
  );
  ShiftS_2 n20 ( // @[Top.scala 145:21]
    .valid_up(n20_valid_up),
    .valid_down(n20_valid_down),
    .I_0(n20_I_0),
    .I_1(n20_I_1),
    .I_2(n20_I_2),
    .I_3(n20_I_3),
    .I_4(n20_I_4),
    .I_5(n20_I_5),
    .I_6(n20_I_6),
    .I_7(n20_I_7),
    .I_8(n20_I_8),
    .I_9(n20_I_9),
    .I_10(n20_I_10),
    .I_11(n20_I_11),
    .I_12(n20_I_12),
    .I_13(n20_I_13),
    .I_14(n20_I_14),
    .I_15(n20_I_15),
    .O_0(n20_O_0),
    .O_1(n20_O_1),
    .O_2(n20_O_2),
    .O_3(n20_O_3),
    .O_4(n20_O_4),
    .O_5(n20_O_5),
    .O_6(n20_O_6),
    .O_7(n20_O_7),
    .O_8(n20_O_8),
    .O_9(n20_O_9),
    .O_10(n20_O_10),
    .O_11(n20_O_11),
    .O_12(n20_O_12),
    .O_13(n20_O_13),
    .O_14(n20_O_14),
    .O_15(n20_O_15)
  );
  ShiftS_2 n21 ( // @[Top.scala 148:21]
    .valid_up(n21_valid_up),
    .valid_down(n21_valid_down),
    .I_0(n21_I_0),
    .I_1(n21_I_1),
    .I_2(n21_I_2),
    .I_3(n21_I_3),
    .I_4(n21_I_4),
    .I_5(n21_I_5),
    .I_6(n21_I_6),
    .I_7(n21_I_7),
    .I_8(n21_I_8),
    .I_9(n21_I_9),
    .I_10(n21_I_10),
    .I_11(n21_I_11),
    .I_12(n21_I_12),
    .I_13(n21_I_13),
    .I_14(n21_I_14),
    .I_15(n21_I_15),
    .O_0(n21_O_0),
    .O_1(n21_O_1),
    .O_2(n21_O_2),
    .O_3(n21_O_3),
    .O_4(n21_O_4),
    .O_5(n21_O_5),
    .O_6(n21_O_6),
    .O_7(n21_O_7),
    .O_8(n21_O_8),
    .O_9(n21_O_9),
    .O_10(n21_O_10),
    .O_11(n21_O_11),
    .O_12(n21_O_12),
    .O_13(n21_O_13),
    .O_14(n21_O_14),
    .O_15(n21_O_15)
  );
  Map2S n22 ( // @[Top.scala 151:21]
    .valid_up(n22_valid_up),
    .valid_down(n22_valid_down),
    .I0_0(n22_I0_0),
    .I0_1(n22_I0_1),
    .I0_2(n22_I0_2),
    .I0_3(n22_I0_3),
    .I0_4(n22_I0_4),
    .I0_5(n22_I0_5),
    .I0_6(n22_I0_6),
    .I0_7(n22_I0_7),
    .I0_8(n22_I0_8),
    .I0_9(n22_I0_9),
    .I0_10(n22_I0_10),
    .I0_11(n22_I0_11),
    .I0_12(n22_I0_12),
    .I0_13(n22_I0_13),
    .I0_14(n22_I0_14),
    .I0_15(n22_I0_15),
    .I1_0(n22_I1_0),
    .I1_1(n22_I1_1),
    .I1_2(n22_I1_2),
    .I1_3(n22_I1_3),
    .I1_4(n22_I1_4),
    .I1_5(n22_I1_5),
    .I1_6(n22_I1_6),
    .I1_7(n22_I1_7),
    .I1_8(n22_I1_8),
    .I1_9(n22_I1_9),
    .I1_10(n22_I1_10),
    .I1_11(n22_I1_11),
    .I1_12(n22_I1_12),
    .I1_13(n22_I1_13),
    .I1_14(n22_I1_14),
    .I1_15(n22_I1_15),
    .O_0_0(n22_O_0_0),
    .O_0_1(n22_O_0_1),
    .O_1_0(n22_O_1_0),
    .O_1_1(n22_O_1_1),
    .O_2_0(n22_O_2_0),
    .O_2_1(n22_O_2_1),
    .O_3_0(n22_O_3_0),
    .O_3_1(n22_O_3_1),
    .O_4_0(n22_O_4_0),
    .O_4_1(n22_O_4_1),
    .O_5_0(n22_O_5_0),
    .O_5_1(n22_O_5_1),
    .O_6_0(n22_O_6_0),
    .O_6_1(n22_O_6_1),
    .O_7_0(n22_O_7_0),
    .O_7_1(n22_O_7_1),
    .O_8_0(n22_O_8_0),
    .O_8_1(n22_O_8_1),
    .O_9_0(n22_O_9_0),
    .O_9_1(n22_O_9_1),
    .O_10_0(n22_O_10_0),
    .O_10_1(n22_O_10_1),
    .O_11_0(n22_O_11_0),
    .O_11_1(n22_O_11_1),
    .O_12_0(n22_O_12_0),
    .O_12_1(n22_O_12_1),
    .O_13_0(n22_O_13_0),
    .O_13_1(n22_O_13_1),
    .O_14_0(n22_O_14_0),
    .O_14_1(n22_O_14_1),
    .O_15_0(n22_O_15_0),
    .O_15_1(n22_O_15_1)
  );
  Map2S_1 n26 ( // @[Top.scala 155:21]
    .valid_up(n26_valid_up),
    .valid_down(n26_valid_down),
    .I0_0_0(n26_I0_0_0),
    .I0_0_1(n26_I0_0_1),
    .I0_1_0(n26_I0_1_0),
    .I0_1_1(n26_I0_1_1),
    .I0_2_0(n26_I0_2_0),
    .I0_2_1(n26_I0_2_1),
    .I0_3_0(n26_I0_3_0),
    .I0_3_1(n26_I0_3_1),
    .I0_4_0(n26_I0_4_0),
    .I0_4_1(n26_I0_4_1),
    .I0_5_0(n26_I0_5_0),
    .I0_5_1(n26_I0_5_1),
    .I0_6_0(n26_I0_6_0),
    .I0_6_1(n26_I0_6_1),
    .I0_7_0(n26_I0_7_0),
    .I0_7_1(n26_I0_7_1),
    .I0_8_0(n26_I0_8_0),
    .I0_8_1(n26_I0_8_1),
    .I0_9_0(n26_I0_9_0),
    .I0_9_1(n26_I0_9_1),
    .I0_10_0(n26_I0_10_0),
    .I0_10_1(n26_I0_10_1),
    .I0_11_0(n26_I0_11_0),
    .I0_11_1(n26_I0_11_1),
    .I0_12_0(n26_I0_12_0),
    .I0_12_1(n26_I0_12_1),
    .I0_13_0(n26_I0_13_0),
    .I0_13_1(n26_I0_13_1),
    .I0_14_0(n26_I0_14_0),
    .I0_14_1(n26_I0_14_1),
    .I0_15_0(n26_I0_15_0),
    .I0_15_1(n26_I0_15_1),
    .I1_0(n26_I1_0),
    .I1_1(n26_I1_1),
    .I1_2(n26_I1_2),
    .I1_3(n26_I1_3),
    .I1_4(n26_I1_4),
    .I1_5(n26_I1_5),
    .I1_6(n26_I1_6),
    .I1_7(n26_I1_7),
    .I1_8(n26_I1_8),
    .I1_9(n26_I1_9),
    .I1_10(n26_I1_10),
    .I1_11(n26_I1_11),
    .I1_12(n26_I1_12),
    .I1_13(n26_I1_13),
    .I1_14(n26_I1_14),
    .I1_15(n26_I1_15),
    .O_0_0(n26_O_0_0),
    .O_0_1(n26_O_0_1),
    .O_0_2(n26_O_0_2),
    .O_1_0(n26_O_1_0),
    .O_1_1(n26_O_1_1),
    .O_1_2(n26_O_1_2),
    .O_2_0(n26_O_2_0),
    .O_2_1(n26_O_2_1),
    .O_2_2(n26_O_2_2),
    .O_3_0(n26_O_3_0),
    .O_3_1(n26_O_3_1),
    .O_3_2(n26_O_3_2),
    .O_4_0(n26_O_4_0),
    .O_4_1(n26_O_4_1),
    .O_4_2(n26_O_4_2),
    .O_5_0(n26_O_5_0),
    .O_5_1(n26_O_5_1),
    .O_5_2(n26_O_5_2),
    .O_6_0(n26_O_6_0),
    .O_6_1(n26_O_6_1),
    .O_6_2(n26_O_6_2),
    .O_7_0(n26_O_7_0),
    .O_7_1(n26_O_7_1),
    .O_7_2(n26_O_7_2),
    .O_8_0(n26_O_8_0),
    .O_8_1(n26_O_8_1),
    .O_8_2(n26_O_8_2),
    .O_9_0(n26_O_9_0),
    .O_9_1(n26_O_9_1),
    .O_9_2(n26_O_9_2),
    .O_10_0(n26_O_10_0),
    .O_10_1(n26_O_10_1),
    .O_10_2(n26_O_10_2),
    .O_11_0(n26_O_11_0),
    .O_11_1(n26_O_11_1),
    .O_11_2(n26_O_11_2),
    .O_12_0(n26_O_12_0),
    .O_12_1(n26_O_12_1),
    .O_12_2(n26_O_12_2),
    .O_13_0(n26_O_13_0),
    .O_13_1(n26_O_13_1),
    .O_13_2(n26_O_13_2),
    .O_14_0(n26_O_14_0),
    .O_14_1(n26_O_14_1),
    .O_14_2(n26_O_14_2),
    .O_15_0(n26_O_15_0),
    .O_15_1(n26_O_15_1),
    .O_15_2(n26_O_15_2)
  );
  PartitionS n30 ( // @[Top.scala 159:21]
    .valid_up(n30_valid_up),
    .valid_down(n30_valid_down),
    .I_0_0(n30_I_0_0),
    .I_0_1(n30_I_0_1),
    .I_0_2(n30_I_0_2),
    .I_1_0(n30_I_1_0),
    .I_1_1(n30_I_1_1),
    .I_1_2(n30_I_1_2),
    .I_2_0(n30_I_2_0),
    .I_2_1(n30_I_2_1),
    .I_2_2(n30_I_2_2),
    .I_3_0(n30_I_3_0),
    .I_3_1(n30_I_3_1),
    .I_3_2(n30_I_3_2),
    .I_4_0(n30_I_4_0),
    .I_4_1(n30_I_4_1),
    .I_4_2(n30_I_4_2),
    .I_5_0(n30_I_5_0),
    .I_5_1(n30_I_5_1),
    .I_5_2(n30_I_5_2),
    .I_6_0(n30_I_6_0),
    .I_6_1(n30_I_6_1),
    .I_6_2(n30_I_6_2),
    .I_7_0(n30_I_7_0),
    .I_7_1(n30_I_7_1),
    .I_7_2(n30_I_7_2),
    .I_8_0(n30_I_8_0),
    .I_8_1(n30_I_8_1),
    .I_8_2(n30_I_8_2),
    .I_9_0(n30_I_9_0),
    .I_9_1(n30_I_9_1),
    .I_9_2(n30_I_9_2),
    .I_10_0(n30_I_10_0),
    .I_10_1(n30_I_10_1),
    .I_10_2(n30_I_10_2),
    .I_11_0(n30_I_11_0),
    .I_11_1(n30_I_11_1),
    .I_11_2(n30_I_11_2),
    .I_12_0(n30_I_12_0),
    .I_12_1(n30_I_12_1),
    .I_12_2(n30_I_12_2),
    .I_13_0(n30_I_13_0),
    .I_13_1(n30_I_13_1),
    .I_13_2(n30_I_13_2),
    .I_14_0(n30_I_14_0),
    .I_14_1(n30_I_14_1),
    .I_14_2(n30_I_14_2),
    .I_15_0(n30_I_15_0),
    .I_15_1(n30_I_15_1),
    .I_15_2(n30_I_15_2),
    .O_0_0_0(n30_O_0_0_0),
    .O_0_0_1(n30_O_0_0_1),
    .O_0_0_2(n30_O_0_0_2),
    .O_1_0_0(n30_O_1_0_0),
    .O_1_0_1(n30_O_1_0_1),
    .O_1_0_2(n30_O_1_0_2),
    .O_2_0_0(n30_O_2_0_0),
    .O_2_0_1(n30_O_2_0_1),
    .O_2_0_2(n30_O_2_0_2),
    .O_3_0_0(n30_O_3_0_0),
    .O_3_0_1(n30_O_3_0_1),
    .O_3_0_2(n30_O_3_0_2),
    .O_4_0_0(n30_O_4_0_0),
    .O_4_0_1(n30_O_4_0_1),
    .O_4_0_2(n30_O_4_0_2),
    .O_5_0_0(n30_O_5_0_0),
    .O_5_0_1(n30_O_5_0_1),
    .O_5_0_2(n30_O_5_0_2),
    .O_6_0_0(n30_O_6_0_0),
    .O_6_0_1(n30_O_6_0_1),
    .O_6_0_2(n30_O_6_0_2),
    .O_7_0_0(n30_O_7_0_0),
    .O_7_0_1(n30_O_7_0_1),
    .O_7_0_2(n30_O_7_0_2),
    .O_8_0_0(n30_O_8_0_0),
    .O_8_0_1(n30_O_8_0_1),
    .O_8_0_2(n30_O_8_0_2),
    .O_9_0_0(n30_O_9_0_0),
    .O_9_0_1(n30_O_9_0_1),
    .O_9_0_2(n30_O_9_0_2),
    .O_10_0_0(n30_O_10_0_0),
    .O_10_0_1(n30_O_10_0_1),
    .O_10_0_2(n30_O_10_0_2),
    .O_11_0_0(n30_O_11_0_0),
    .O_11_0_1(n30_O_11_0_1),
    .O_11_0_2(n30_O_11_0_2),
    .O_12_0_0(n30_O_12_0_0),
    .O_12_0_1(n30_O_12_0_1),
    .O_12_0_2(n30_O_12_0_2),
    .O_13_0_0(n30_O_13_0_0),
    .O_13_0_1(n30_O_13_0_1),
    .O_13_0_2(n30_O_13_0_2),
    .O_14_0_0(n30_O_14_0_0),
    .O_14_0_1(n30_O_14_0_1),
    .O_14_0_2(n30_O_14_0_2),
    .O_15_0_0(n30_O_15_0_0),
    .O_15_0_1(n30_O_15_0_1),
    .O_15_0_2(n30_O_15_0_2)
  );
  MapS n35 ( // @[Top.scala 162:21]
    .valid_up(n35_valid_up),
    .valid_down(n35_valid_down),
    .I_0_0_0(n35_I_0_0_0),
    .I_0_0_1(n35_I_0_0_1),
    .I_0_0_2(n35_I_0_0_2),
    .I_1_0_0(n35_I_1_0_0),
    .I_1_0_1(n35_I_1_0_1),
    .I_1_0_2(n35_I_1_0_2),
    .I_2_0_0(n35_I_2_0_0),
    .I_2_0_1(n35_I_2_0_1),
    .I_2_0_2(n35_I_2_0_2),
    .I_3_0_0(n35_I_3_0_0),
    .I_3_0_1(n35_I_3_0_1),
    .I_3_0_2(n35_I_3_0_2),
    .I_4_0_0(n35_I_4_0_0),
    .I_4_0_1(n35_I_4_0_1),
    .I_4_0_2(n35_I_4_0_2),
    .I_5_0_0(n35_I_5_0_0),
    .I_5_0_1(n35_I_5_0_1),
    .I_5_0_2(n35_I_5_0_2),
    .I_6_0_0(n35_I_6_0_0),
    .I_6_0_1(n35_I_6_0_1),
    .I_6_0_2(n35_I_6_0_2),
    .I_7_0_0(n35_I_7_0_0),
    .I_7_0_1(n35_I_7_0_1),
    .I_7_0_2(n35_I_7_0_2),
    .I_8_0_0(n35_I_8_0_0),
    .I_8_0_1(n35_I_8_0_1),
    .I_8_0_2(n35_I_8_0_2),
    .I_9_0_0(n35_I_9_0_0),
    .I_9_0_1(n35_I_9_0_1),
    .I_9_0_2(n35_I_9_0_2),
    .I_10_0_0(n35_I_10_0_0),
    .I_10_0_1(n35_I_10_0_1),
    .I_10_0_2(n35_I_10_0_2),
    .I_11_0_0(n35_I_11_0_0),
    .I_11_0_1(n35_I_11_0_1),
    .I_11_0_2(n35_I_11_0_2),
    .I_12_0_0(n35_I_12_0_0),
    .I_12_0_1(n35_I_12_0_1),
    .I_12_0_2(n35_I_12_0_2),
    .I_13_0_0(n35_I_13_0_0),
    .I_13_0_1(n35_I_13_0_1),
    .I_13_0_2(n35_I_13_0_2),
    .I_14_0_0(n35_I_14_0_0),
    .I_14_0_1(n35_I_14_0_1),
    .I_14_0_2(n35_I_14_0_2),
    .I_15_0_0(n35_I_15_0_0),
    .I_15_0_1(n35_I_15_0_1),
    .I_15_0_2(n35_I_15_0_2),
    .O_0_0(n35_O_0_0),
    .O_0_1(n35_O_0_1),
    .O_0_2(n35_O_0_2),
    .O_1_0(n35_O_1_0),
    .O_1_1(n35_O_1_1),
    .O_1_2(n35_O_1_2),
    .O_2_0(n35_O_2_0),
    .O_2_1(n35_O_2_1),
    .O_2_2(n35_O_2_2),
    .O_3_0(n35_O_3_0),
    .O_3_1(n35_O_3_1),
    .O_3_2(n35_O_3_2),
    .O_4_0(n35_O_4_0),
    .O_4_1(n35_O_4_1),
    .O_4_2(n35_O_4_2),
    .O_5_0(n35_O_5_0),
    .O_5_1(n35_O_5_1),
    .O_5_2(n35_O_5_2),
    .O_6_0(n35_O_6_0),
    .O_6_1(n35_O_6_1),
    .O_6_2(n35_O_6_2),
    .O_7_0(n35_O_7_0),
    .O_7_1(n35_O_7_1),
    .O_7_2(n35_O_7_2),
    .O_8_0(n35_O_8_0),
    .O_8_1(n35_O_8_1),
    .O_8_2(n35_O_8_2),
    .O_9_0(n35_O_9_0),
    .O_9_1(n35_O_9_1),
    .O_9_2(n35_O_9_2),
    .O_10_0(n35_O_10_0),
    .O_10_1(n35_O_10_1),
    .O_10_2(n35_O_10_2),
    .O_11_0(n35_O_11_0),
    .O_11_1(n35_O_11_1),
    .O_11_2(n35_O_11_2),
    .O_12_0(n35_O_12_0),
    .O_12_1(n35_O_12_1),
    .O_12_2(n35_O_12_2),
    .O_13_0(n35_O_13_0),
    .O_13_1(n35_O_13_1),
    .O_13_2(n35_O_13_2),
    .O_14_0(n35_O_14_0),
    .O_14_1(n35_O_14_1),
    .O_14_2(n35_O_14_2),
    .O_15_0(n35_O_15_0),
    .O_15_1(n35_O_15_1),
    .O_15_2(n35_O_15_2)
  );
  Map2S_4 n36 ( // @[Top.scala 165:21]
    .valid_up(n36_valid_up),
    .valid_down(n36_valid_down),
    .I0_0_0(n36_I0_0_0),
    .I0_0_1(n36_I0_0_1),
    .I0_0_2(n36_I0_0_2),
    .I0_1_0(n36_I0_1_0),
    .I0_1_1(n36_I0_1_1),
    .I0_1_2(n36_I0_1_2),
    .I0_2_0(n36_I0_2_0),
    .I0_2_1(n36_I0_2_1),
    .I0_2_2(n36_I0_2_2),
    .I0_3_0(n36_I0_3_0),
    .I0_3_1(n36_I0_3_1),
    .I0_3_2(n36_I0_3_2),
    .I0_4_0(n36_I0_4_0),
    .I0_4_1(n36_I0_4_1),
    .I0_4_2(n36_I0_4_2),
    .I0_5_0(n36_I0_5_0),
    .I0_5_1(n36_I0_5_1),
    .I0_5_2(n36_I0_5_2),
    .I0_6_0(n36_I0_6_0),
    .I0_6_1(n36_I0_6_1),
    .I0_6_2(n36_I0_6_2),
    .I0_7_0(n36_I0_7_0),
    .I0_7_1(n36_I0_7_1),
    .I0_7_2(n36_I0_7_2),
    .I0_8_0(n36_I0_8_0),
    .I0_8_1(n36_I0_8_1),
    .I0_8_2(n36_I0_8_2),
    .I0_9_0(n36_I0_9_0),
    .I0_9_1(n36_I0_9_1),
    .I0_9_2(n36_I0_9_2),
    .I0_10_0(n36_I0_10_0),
    .I0_10_1(n36_I0_10_1),
    .I0_10_2(n36_I0_10_2),
    .I0_11_0(n36_I0_11_0),
    .I0_11_1(n36_I0_11_1),
    .I0_11_2(n36_I0_11_2),
    .I0_12_0(n36_I0_12_0),
    .I0_12_1(n36_I0_12_1),
    .I0_12_2(n36_I0_12_2),
    .I0_13_0(n36_I0_13_0),
    .I0_13_1(n36_I0_13_1),
    .I0_13_2(n36_I0_13_2),
    .I0_14_0(n36_I0_14_0),
    .I0_14_1(n36_I0_14_1),
    .I0_14_2(n36_I0_14_2),
    .I0_15_0(n36_I0_15_0),
    .I0_15_1(n36_I0_15_1),
    .I0_15_2(n36_I0_15_2),
    .I1_0_0(n36_I1_0_0),
    .I1_0_1(n36_I1_0_1),
    .I1_0_2(n36_I1_0_2),
    .I1_1_0(n36_I1_1_0),
    .I1_1_1(n36_I1_1_1),
    .I1_1_2(n36_I1_1_2),
    .I1_2_0(n36_I1_2_0),
    .I1_2_1(n36_I1_2_1),
    .I1_2_2(n36_I1_2_2),
    .I1_3_0(n36_I1_3_0),
    .I1_3_1(n36_I1_3_1),
    .I1_3_2(n36_I1_3_2),
    .I1_4_0(n36_I1_4_0),
    .I1_4_1(n36_I1_4_1),
    .I1_4_2(n36_I1_4_2),
    .I1_5_0(n36_I1_5_0),
    .I1_5_1(n36_I1_5_1),
    .I1_5_2(n36_I1_5_2),
    .I1_6_0(n36_I1_6_0),
    .I1_6_1(n36_I1_6_1),
    .I1_6_2(n36_I1_6_2),
    .I1_7_0(n36_I1_7_0),
    .I1_7_1(n36_I1_7_1),
    .I1_7_2(n36_I1_7_2),
    .I1_8_0(n36_I1_8_0),
    .I1_8_1(n36_I1_8_1),
    .I1_8_2(n36_I1_8_2),
    .I1_9_0(n36_I1_9_0),
    .I1_9_1(n36_I1_9_1),
    .I1_9_2(n36_I1_9_2),
    .I1_10_0(n36_I1_10_0),
    .I1_10_1(n36_I1_10_1),
    .I1_10_2(n36_I1_10_2),
    .I1_11_0(n36_I1_11_0),
    .I1_11_1(n36_I1_11_1),
    .I1_11_2(n36_I1_11_2),
    .I1_12_0(n36_I1_12_0),
    .I1_12_1(n36_I1_12_1),
    .I1_12_2(n36_I1_12_2),
    .I1_13_0(n36_I1_13_0),
    .I1_13_1(n36_I1_13_1),
    .I1_13_2(n36_I1_13_2),
    .I1_14_0(n36_I1_14_0),
    .I1_14_1(n36_I1_14_1),
    .I1_14_2(n36_I1_14_2),
    .I1_15_0(n36_I1_15_0),
    .I1_15_1(n36_I1_15_1),
    .I1_15_2(n36_I1_15_2),
    .O_0_0_0(n36_O_0_0_0),
    .O_0_0_1(n36_O_0_0_1),
    .O_0_0_2(n36_O_0_0_2),
    .O_0_1_0(n36_O_0_1_0),
    .O_0_1_1(n36_O_0_1_1),
    .O_0_1_2(n36_O_0_1_2),
    .O_1_0_0(n36_O_1_0_0),
    .O_1_0_1(n36_O_1_0_1),
    .O_1_0_2(n36_O_1_0_2),
    .O_1_1_0(n36_O_1_1_0),
    .O_1_1_1(n36_O_1_1_1),
    .O_1_1_2(n36_O_1_1_2),
    .O_2_0_0(n36_O_2_0_0),
    .O_2_0_1(n36_O_2_0_1),
    .O_2_0_2(n36_O_2_0_2),
    .O_2_1_0(n36_O_2_1_0),
    .O_2_1_1(n36_O_2_1_1),
    .O_2_1_2(n36_O_2_1_2),
    .O_3_0_0(n36_O_3_0_0),
    .O_3_0_1(n36_O_3_0_1),
    .O_3_0_2(n36_O_3_0_2),
    .O_3_1_0(n36_O_3_1_0),
    .O_3_1_1(n36_O_3_1_1),
    .O_3_1_2(n36_O_3_1_2),
    .O_4_0_0(n36_O_4_0_0),
    .O_4_0_1(n36_O_4_0_1),
    .O_4_0_2(n36_O_4_0_2),
    .O_4_1_0(n36_O_4_1_0),
    .O_4_1_1(n36_O_4_1_1),
    .O_4_1_2(n36_O_4_1_2),
    .O_5_0_0(n36_O_5_0_0),
    .O_5_0_1(n36_O_5_0_1),
    .O_5_0_2(n36_O_5_0_2),
    .O_5_1_0(n36_O_5_1_0),
    .O_5_1_1(n36_O_5_1_1),
    .O_5_1_2(n36_O_5_1_2),
    .O_6_0_0(n36_O_6_0_0),
    .O_6_0_1(n36_O_6_0_1),
    .O_6_0_2(n36_O_6_0_2),
    .O_6_1_0(n36_O_6_1_0),
    .O_6_1_1(n36_O_6_1_1),
    .O_6_1_2(n36_O_6_1_2),
    .O_7_0_0(n36_O_7_0_0),
    .O_7_0_1(n36_O_7_0_1),
    .O_7_0_2(n36_O_7_0_2),
    .O_7_1_0(n36_O_7_1_0),
    .O_7_1_1(n36_O_7_1_1),
    .O_7_1_2(n36_O_7_1_2),
    .O_8_0_0(n36_O_8_0_0),
    .O_8_0_1(n36_O_8_0_1),
    .O_8_0_2(n36_O_8_0_2),
    .O_8_1_0(n36_O_8_1_0),
    .O_8_1_1(n36_O_8_1_1),
    .O_8_1_2(n36_O_8_1_2),
    .O_9_0_0(n36_O_9_0_0),
    .O_9_0_1(n36_O_9_0_1),
    .O_9_0_2(n36_O_9_0_2),
    .O_9_1_0(n36_O_9_1_0),
    .O_9_1_1(n36_O_9_1_1),
    .O_9_1_2(n36_O_9_1_2),
    .O_10_0_0(n36_O_10_0_0),
    .O_10_0_1(n36_O_10_0_1),
    .O_10_0_2(n36_O_10_0_2),
    .O_10_1_0(n36_O_10_1_0),
    .O_10_1_1(n36_O_10_1_1),
    .O_10_1_2(n36_O_10_1_2),
    .O_11_0_0(n36_O_11_0_0),
    .O_11_0_1(n36_O_11_0_1),
    .O_11_0_2(n36_O_11_0_2),
    .O_11_1_0(n36_O_11_1_0),
    .O_11_1_1(n36_O_11_1_1),
    .O_11_1_2(n36_O_11_1_2),
    .O_12_0_0(n36_O_12_0_0),
    .O_12_0_1(n36_O_12_0_1),
    .O_12_0_2(n36_O_12_0_2),
    .O_12_1_0(n36_O_12_1_0),
    .O_12_1_1(n36_O_12_1_1),
    .O_12_1_2(n36_O_12_1_2),
    .O_13_0_0(n36_O_13_0_0),
    .O_13_0_1(n36_O_13_0_1),
    .O_13_0_2(n36_O_13_0_2),
    .O_13_1_0(n36_O_13_1_0),
    .O_13_1_1(n36_O_13_1_1),
    .O_13_1_2(n36_O_13_1_2),
    .O_14_0_0(n36_O_14_0_0),
    .O_14_0_1(n36_O_14_0_1),
    .O_14_0_2(n36_O_14_0_2),
    .O_14_1_0(n36_O_14_1_0),
    .O_14_1_1(n36_O_14_1_1),
    .O_14_1_2(n36_O_14_1_2),
    .O_15_0_0(n36_O_15_0_0),
    .O_15_0_1(n36_O_15_0_1),
    .O_15_0_2(n36_O_15_0_2),
    .O_15_1_0(n36_O_15_1_0),
    .O_15_1_1(n36_O_15_1_1),
    .O_15_1_2(n36_O_15_1_2)
  );
  ShiftS_2 n40 ( // @[Top.scala 169:21]
    .valid_up(n40_valid_up),
    .valid_down(n40_valid_down),
    .I_0(n40_I_0),
    .I_1(n40_I_1),
    .I_2(n40_I_2),
    .I_3(n40_I_3),
    .I_4(n40_I_4),
    .I_5(n40_I_5),
    .I_6(n40_I_6),
    .I_7(n40_I_7),
    .I_8(n40_I_8),
    .I_9(n40_I_9),
    .I_10(n40_I_10),
    .I_11(n40_I_11),
    .I_12(n40_I_12),
    .I_13(n40_I_13),
    .I_14(n40_I_14),
    .I_15(n40_I_15),
    .O_0(n40_O_0),
    .O_1(n40_O_1),
    .O_2(n40_O_2),
    .O_3(n40_O_3),
    .O_4(n40_O_4),
    .O_5(n40_O_5),
    .O_6(n40_O_6),
    .O_7(n40_O_7),
    .O_8(n40_O_8),
    .O_9(n40_O_9),
    .O_10(n40_O_10),
    .O_11(n40_O_11),
    .O_12(n40_O_12),
    .O_13(n40_O_13),
    .O_14(n40_O_14),
    .O_15(n40_O_15)
  );
  ShiftS_2 n41 ( // @[Top.scala 172:21]
    .valid_up(n41_valid_up),
    .valid_down(n41_valid_down),
    .I_0(n41_I_0),
    .I_1(n41_I_1),
    .I_2(n41_I_2),
    .I_3(n41_I_3),
    .I_4(n41_I_4),
    .I_5(n41_I_5),
    .I_6(n41_I_6),
    .I_7(n41_I_7),
    .I_8(n41_I_8),
    .I_9(n41_I_9),
    .I_10(n41_I_10),
    .I_11(n41_I_11),
    .I_12(n41_I_12),
    .I_13(n41_I_13),
    .I_14(n41_I_14),
    .I_15(n41_I_15),
    .O_0(n41_O_0),
    .O_1(n41_O_1),
    .O_2(n41_O_2),
    .O_3(n41_O_3),
    .O_4(n41_O_4),
    .O_5(n41_O_5),
    .O_6(n41_O_6),
    .O_7(n41_O_7),
    .O_8(n41_O_8),
    .O_9(n41_O_9),
    .O_10(n41_O_10),
    .O_11(n41_O_11),
    .O_12(n41_O_12),
    .O_13(n41_O_13),
    .O_14(n41_O_14),
    .O_15(n41_O_15)
  );
  Map2S n42 ( // @[Top.scala 175:21]
    .valid_up(n42_valid_up),
    .valid_down(n42_valid_down),
    .I0_0(n42_I0_0),
    .I0_1(n42_I0_1),
    .I0_2(n42_I0_2),
    .I0_3(n42_I0_3),
    .I0_4(n42_I0_4),
    .I0_5(n42_I0_5),
    .I0_6(n42_I0_6),
    .I0_7(n42_I0_7),
    .I0_8(n42_I0_8),
    .I0_9(n42_I0_9),
    .I0_10(n42_I0_10),
    .I0_11(n42_I0_11),
    .I0_12(n42_I0_12),
    .I0_13(n42_I0_13),
    .I0_14(n42_I0_14),
    .I0_15(n42_I0_15),
    .I1_0(n42_I1_0),
    .I1_1(n42_I1_1),
    .I1_2(n42_I1_2),
    .I1_3(n42_I1_3),
    .I1_4(n42_I1_4),
    .I1_5(n42_I1_5),
    .I1_6(n42_I1_6),
    .I1_7(n42_I1_7),
    .I1_8(n42_I1_8),
    .I1_9(n42_I1_9),
    .I1_10(n42_I1_10),
    .I1_11(n42_I1_11),
    .I1_12(n42_I1_12),
    .I1_13(n42_I1_13),
    .I1_14(n42_I1_14),
    .I1_15(n42_I1_15),
    .O_0_0(n42_O_0_0),
    .O_0_1(n42_O_0_1),
    .O_1_0(n42_O_1_0),
    .O_1_1(n42_O_1_1),
    .O_2_0(n42_O_2_0),
    .O_2_1(n42_O_2_1),
    .O_3_0(n42_O_3_0),
    .O_3_1(n42_O_3_1),
    .O_4_0(n42_O_4_0),
    .O_4_1(n42_O_4_1),
    .O_5_0(n42_O_5_0),
    .O_5_1(n42_O_5_1),
    .O_6_0(n42_O_6_0),
    .O_6_1(n42_O_6_1),
    .O_7_0(n42_O_7_0),
    .O_7_1(n42_O_7_1),
    .O_8_0(n42_O_8_0),
    .O_8_1(n42_O_8_1),
    .O_9_0(n42_O_9_0),
    .O_9_1(n42_O_9_1),
    .O_10_0(n42_O_10_0),
    .O_10_1(n42_O_10_1),
    .O_11_0(n42_O_11_0),
    .O_11_1(n42_O_11_1),
    .O_12_0(n42_O_12_0),
    .O_12_1(n42_O_12_1),
    .O_13_0(n42_O_13_0),
    .O_13_1(n42_O_13_1),
    .O_14_0(n42_O_14_0),
    .O_14_1(n42_O_14_1),
    .O_15_0(n42_O_15_0),
    .O_15_1(n42_O_15_1)
  );
  Map2S_1 n46 ( // @[Top.scala 179:21]
    .valid_up(n46_valid_up),
    .valid_down(n46_valid_down),
    .I0_0_0(n46_I0_0_0),
    .I0_0_1(n46_I0_0_1),
    .I0_1_0(n46_I0_1_0),
    .I0_1_1(n46_I0_1_1),
    .I0_2_0(n46_I0_2_0),
    .I0_2_1(n46_I0_2_1),
    .I0_3_0(n46_I0_3_0),
    .I0_3_1(n46_I0_3_1),
    .I0_4_0(n46_I0_4_0),
    .I0_4_1(n46_I0_4_1),
    .I0_5_0(n46_I0_5_0),
    .I0_5_1(n46_I0_5_1),
    .I0_6_0(n46_I0_6_0),
    .I0_6_1(n46_I0_6_1),
    .I0_7_0(n46_I0_7_0),
    .I0_7_1(n46_I0_7_1),
    .I0_8_0(n46_I0_8_0),
    .I0_8_1(n46_I0_8_1),
    .I0_9_0(n46_I0_9_0),
    .I0_9_1(n46_I0_9_1),
    .I0_10_0(n46_I0_10_0),
    .I0_10_1(n46_I0_10_1),
    .I0_11_0(n46_I0_11_0),
    .I0_11_1(n46_I0_11_1),
    .I0_12_0(n46_I0_12_0),
    .I0_12_1(n46_I0_12_1),
    .I0_13_0(n46_I0_13_0),
    .I0_13_1(n46_I0_13_1),
    .I0_14_0(n46_I0_14_0),
    .I0_14_1(n46_I0_14_1),
    .I0_15_0(n46_I0_15_0),
    .I0_15_1(n46_I0_15_1),
    .I1_0(n46_I1_0),
    .I1_1(n46_I1_1),
    .I1_2(n46_I1_2),
    .I1_3(n46_I1_3),
    .I1_4(n46_I1_4),
    .I1_5(n46_I1_5),
    .I1_6(n46_I1_6),
    .I1_7(n46_I1_7),
    .I1_8(n46_I1_8),
    .I1_9(n46_I1_9),
    .I1_10(n46_I1_10),
    .I1_11(n46_I1_11),
    .I1_12(n46_I1_12),
    .I1_13(n46_I1_13),
    .I1_14(n46_I1_14),
    .I1_15(n46_I1_15),
    .O_0_0(n46_O_0_0),
    .O_0_1(n46_O_0_1),
    .O_0_2(n46_O_0_2),
    .O_1_0(n46_O_1_0),
    .O_1_1(n46_O_1_1),
    .O_1_2(n46_O_1_2),
    .O_2_0(n46_O_2_0),
    .O_2_1(n46_O_2_1),
    .O_2_2(n46_O_2_2),
    .O_3_0(n46_O_3_0),
    .O_3_1(n46_O_3_1),
    .O_3_2(n46_O_3_2),
    .O_4_0(n46_O_4_0),
    .O_4_1(n46_O_4_1),
    .O_4_2(n46_O_4_2),
    .O_5_0(n46_O_5_0),
    .O_5_1(n46_O_5_1),
    .O_5_2(n46_O_5_2),
    .O_6_0(n46_O_6_0),
    .O_6_1(n46_O_6_1),
    .O_6_2(n46_O_6_2),
    .O_7_0(n46_O_7_0),
    .O_7_1(n46_O_7_1),
    .O_7_2(n46_O_7_2),
    .O_8_0(n46_O_8_0),
    .O_8_1(n46_O_8_1),
    .O_8_2(n46_O_8_2),
    .O_9_0(n46_O_9_0),
    .O_9_1(n46_O_9_1),
    .O_9_2(n46_O_9_2),
    .O_10_0(n46_O_10_0),
    .O_10_1(n46_O_10_1),
    .O_10_2(n46_O_10_2),
    .O_11_0(n46_O_11_0),
    .O_11_1(n46_O_11_1),
    .O_11_2(n46_O_11_2),
    .O_12_0(n46_O_12_0),
    .O_12_1(n46_O_12_1),
    .O_12_2(n46_O_12_2),
    .O_13_0(n46_O_13_0),
    .O_13_1(n46_O_13_1),
    .O_13_2(n46_O_13_2),
    .O_14_0(n46_O_14_0),
    .O_14_1(n46_O_14_1),
    .O_14_2(n46_O_14_2),
    .O_15_0(n46_O_15_0),
    .O_15_1(n46_O_15_1),
    .O_15_2(n46_O_15_2)
  );
  PartitionS n50 ( // @[Top.scala 183:21]
    .valid_up(n50_valid_up),
    .valid_down(n50_valid_down),
    .I_0_0(n50_I_0_0),
    .I_0_1(n50_I_0_1),
    .I_0_2(n50_I_0_2),
    .I_1_0(n50_I_1_0),
    .I_1_1(n50_I_1_1),
    .I_1_2(n50_I_1_2),
    .I_2_0(n50_I_2_0),
    .I_2_1(n50_I_2_1),
    .I_2_2(n50_I_2_2),
    .I_3_0(n50_I_3_0),
    .I_3_1(n50_I_3_1),
    .I_3_2(n50_I_3_2),
    .I_4_0(n50_I_4_0),
    .I_4_1(n50_I_4_1),
    .I_4_2(n50_I_4_2),
    .I_5_0(n50_I_5_0),
    .I_5_1(n50_I_5_1),
    .I_5_2(n50_I_5_2),
    .I_6_0(n50_I_6_0),
    .I_6_1(n50_I_6_1),
    .I_6_2(n50_I_6_2),
    .I_7_0(n50_I_7_0),
    .I_7_1(n50_I_7_1),
    .I_7_2(n50_I_7_2),
    .I_8_0(n50_I_8_0),
    .I_8_1(n50_I_8_1),
    .I_8_2(n50_I_8_2),
    .I_9_0(n50_I_9_0),
    .I_9_1(n50_I_9_1),
    .I_9_2(n50_I_9_2),
    .I_10_0(n50_I_10_0),
    .I_10_1(n50_I_10_1),
    .I_10_2(n50_I_10_2),
    .I_11_0(n50_I_11_0),
    .I_11_1(n50_I_11_1),
    .I_11_2(n50_I_11_2),
    .I_12_0(n50_I_12_0),
    .I_12_1(n50_I_12_1),
    .I_12_2(n50_I_12_2),
    .I_13_0(n50_I_13_0),
    .I_13_1(n50_I_13_1),
    .I_13_2(n50_I_13_2),
    .I_14_0(n50_I_14_0),
    .I_14_1(n50_I_14_1),
    .I_14_2(n50_I_14_2),
    .I_15_0(n50_I_15_0),
    .I_15_1(n50_I_15_1),
    .I_15_2(n50_I_15_2),
    .O_0_0_0(n50_O_0_0_0),
    .O_0_0_1(n50_O_0_0_1),
    .O_0_0_2(n50_O_0_0_2),
    .O_1_0_0(n50_O_1_0_0),
    .O_1_0_1(n50_O_1_0_1),
    .O_1_0_2(n50_O_1_0_2),
    .O_2_0_0(n50_O_2_0_0),
    .O_2_0_1(n50_O_2_0_1),
    .O_2_0_2(n50_O_2_0_2),
    .O_3_0_0(n50_O_3_0_0),
    .O_3_0_1(n50_O_3_0_1),
    .O_3_0_2(n50_O_3_0_2),
    .O_4_0_0(n50_O_4_0_0),
    .O_4_0_1(n50_O_4_0_1),
    .O_4_0_2(n50_O_4_0_2),
    .O_5_0_0(n50_O_5_0_0),
    .O_5_0_1(n50_O_5_0_1),
    .O_5_0_2(n50_O_5_0_2),
    .O_6_0_0(n50_O_6_0_0),
    .O_6_0_1(n50_O_6_0_1),
    .O_6_0_2(n50_O_6_0_2),
    .O_7_0_0(n50_O_7_0_0),
    .O_7_0_1(n50_O_7_0_1),
    .O_7_0_2(n50_O_7_0_2),
    .O_8_0_0(n50_O_8_0_0),
    .O_8_0_1(n50_O_8_0_1),
    .O_8_0_2(n50_O_8_0_2),
    .O_9_0_0(n50_O_9_0_0),
    .O_9_0_1(n50_O_9_0_1),
    .O_9_0_2(n50_O_9_0_2),
    .O_10_0_0(n50_O_10_0_0),
    .O_10_0_1(n50_O_10_0_1),
    .O_10_0_2(n50_O_10_0_2),
    .O_11_0_0(n50_O_11_0_0),
    .O_11_0_1(n50_O_11_0_1),
    .O_11_0_2(n50_O_11_0_2),
    .O_12_0_0(n50_O_12_0_0),
    .O_12_0_1(n50_O_12_0_1),
    .O_12_0_2(n50_O_12_0_2),
    .O_13_0_0(n50_O_13_0_0),
    .O_13_0_1(n50_O_13_0_1),
    .O_13_0_2(n50_O_13_0_2),
    .O_14_0_0(n50_O_14_0_0),
    .O_14_0_1(n50_O_14_0_1),
    .O_14_0_2(n50_O_14_0_2),
    .O_15_0_0(n50_O_15_0_0),
    .O_15_0_1(n50_O_15_0_1),
    .O_15_0_2(n50_O_15_0_2)
  );
  MapS n55 ( // @[Top.scala 186:21]
    .valid_up(n55_valid_up),
    .valid_down(n55_valid_down),
    .I_0_0_0(n55_I_0_0_0),
    .I_0_0_1(n55_I_0_0_1),
    .I_0_0_2(n55_I_0_0_2),
    .I_1_0_0(n55_I_1_0_0),
    .I_1_0_1(n55_I_1_0_1),
    .I_1_0_2(n55_I_1_0_2),
    .I_2_0_0(n55_I_2_0_0),
    .I_2_0_1(n55_I_2_0_1),
    .I_2_0_2(n55_I_2_0_2),
    .I_3_0_0(n55_I_3_0_0),
    .I_3_0_1(n55_I_3_0_1),
    .I_3_0_2(n55_I_3_0_2),
    .I_4_0_0(n55_I_4_0_0),
    .I_4_0_1(n55_I_4_0_1),
    .I_4_0_2(n55_I_4_0_2),
    .I_5_0_0(n55_I_5_0_0),
    .I_5_0_1(n55_I_5_0_1),
    .I_5_0_2(n55_I_5_0_2),
    .I_6_0_0(n55_I_6_0_0),
    .I_6_0_1(n55_I_6_0_1),
    .I_6_0_2(n55_I_6_0_2),
    .I_7_0_0(n55_I_7_0_0),
    .I_7_0_1(n55_I_7_0_1),
    .I_7_0_2(n55_I_7_0_2),
    .I_8_0_0(n55_I_8_0_0),
    .I_8_0_1(n55_I_8_0_1),
    .I_8_0_2(n55_I_8_0_2),
    .I_9_0_0(n55_I_9_0_0),
    .I_9_0_1(n55_I_9_0_1),
    .I_9_0_2(n55_I_9_0_2),
    .I_10_0_0(n55_I_10_0_0),
    .I_10_0_1(n55_I_10_0_1),
    .I_10_0_2(n55_I_10_0_2),
    .I_11_0_0(n55_I_11_0_0),
    .I_11_0_1(n55_I_11_0_1),
    .I_11_0_2(n55_I_11_0_2),
    .I_12_0_0(n55_I_12_0_0),
    .I_12_0_1(n55_I_12_0_1),
    .I_12_0_2(n55_I_12_0_2),
    .I_13_0_0(n55_I_13_0_0),
    .I_13_0_1(n55_I_13_0_1),
    .I_13_0_2(n55_I_13_0_2),
    .I_14_0_0(n55_I_14_0_0),
    .I_14_0_1(n55_I_14_0_1),
    .I_14_0_2(n55_I_14_0_2),
    .I_15_0_0(n55_I_15_0_0),
    .I_15_0_1(n55_I_15_0_1),
    .I_15_0_2(n55_I_15_0_2),
    .O_0_0(n55_O_0_0),
    .O_0_1(n55_O_0_1),
    .O_0_2(n55_O_0_2),
    .O_1_0(n55_O_1_0),
    .O_1_1(n55_O_1_1),
    .O_1_2(n55_O_1_2),
    .O_2_0(n55_O_2_0),
    .O_2_1(n55_O_2_1),
    .O_2_2(n55_O_2_2),
    .O_3_0(n55_O_3_0),
    .O_3_1(n55_O_3_1),
    .O_3_2(n55_O_3_2),
    .O_4_0(n55_O_4_0),
    .O_4_1(n55_O_4_1),
    .O_4_2(n55_O_4_2),
    .O_5_0(n55_O_5_0),
    .O_5_1(n55_O_5_1),
    .O_5_2(n55_O_5_2),
    .O_6_0(n55_O_6_0),
    .O_6_1(n55_O_6_1),
    .O_6_2(n55_O_6_2),
    .O_7_0(n55_O_7_0),
    .O_7_1(n55_O_7_1),
    .O_7_2(n55_O_7_2),
    .O_8_0(n55_O_8_0),
    .O_8_1(n55_O_8_1),
    .O_8_2(n55_O_8_2),
    .O_9_0(n55_O_9_0),
    .O_9_1(n55_O_9_1),
    .O_9_2(n55_O_9_2),
    .O_10_0(n55_O_10_0),
    .O_10_1(n55_O_10_1),
    .O_10_2(n55_O_10_2),
    .O_11_0(n55_O_11_0),
    .O_11_1(n55_O_11_1),
    .O_11_2(n55_O_11_2),
    .O_12_0(n55_O_12_0),
    .O_12_1(n55_O_12_1),
    .O_12_2(n55_O_12_2),
    .O_13_0(n55_O_13_0),
    .O_13_1(n55_O_13_1),
    .O_13_2(n55_O_13_2),
    .O_14_0(n55_O_14_0),
    .O_14_1(n55_O_14_1),
    .O_14_2(n55_O_14_2),
    .O_15_0(n55_O_15_0),
    .O_15_1(n55_O_15_1),
    .O_15_2(n55_O_15_2)
  );
  Map2S_7 n56 ( // @[Top.scala 189:21]
    .valid_up(n56_valid_up),
    .valid_down(n56_valid_down),
    .I0_0_0_0(n56_I0_0_0_0),
    .I0_0_0_1(n56_I0_0_0_1),
    .I0_0_0_2(n56_I0_0_0_2),
    .I0_0_1_0(n56_I0_0_1_0),
    .I0_0_1_1(n56_I0_0_1_1),
    .I0_0_1_2(n56_I0_0_1_2),
    .I0_1_0_0(n56_I0_1_0_0),
    .I0_1_0_1(n56_I0_1_0_1),
    .I0_1_0_2(n56_I0_1_0_2),
    .I0_1_1_0(n56_I0_1_1_0),
    .I0_1_1_1(n56_I0_1_1_1),
    .I0_1_1_2(n56_I0_1_1_2),
    .I0_2_0_0(n56_I0_2_0_0),
    .I0_2_0_1(n56_I0_2_0_1),
    .I0_2_0_2(n56_I0_2_0_2),
    .I0_2_1_0(n56_I0_2_1_0),
    .I0_2_1_1(n56_I0_2_1_1),
    .I0_2_1_2(n56_I0_2_1_2),
    .I0_3_0_0(n56_I0_3_0_0),
    .I0_3_0_1(n56_I0_3_0_1),
    .I0_3_0_2(n56_I0_3_0_2),
    .I0_3_1_0(n56_I0_3_1_0),
    .I0_3_1_1(n56_I0_3_1_1),
    .I0_3_1_2(n56_I0_3_1_2),
    .I0_4_0_0(n56_I0_4_0_0),
    .I0_4_0_1(n56_I0_4_0_1),
    .I0_4_0_2(n56_I0_4_0_2),
    .I0_4_1_0(n56_I0_4_1_0),
    .I0_4_1_1(n56_I0_4_1_1),
    .I0_4_1_2(n56_I0_4_1_2),
    .I0_5_0_0(n56_I0_5_0_0),
    .I0_5_0_1(n56_I0_5_0_1),
    .I0_5_0_2(n56_I0_5_0_2),
    .I0_5_1_0(n56_I0_5_1_0),
    .I0_5_1_1(n56_I0_5_1_1),
    .I0_5_1_2(n56_I0_5_1_2),
    .I0_6_0_0(n56_I0_6_0_0),
    .I0_6_0_1(n56_I0_6_0_1),
    .I0_6_0_2(n56_I0_6_0_2),
    .I0_6_1_0(n56_I0_6_1_0),
    .I0_6_1_1(n56_I0_6_1_1),
    .I0_6_1_2(n56_I0_6_1_2),
    .I0_7_0_0(n56_I0_7_0_0),
    .I0_7_0_1(n56_I0_7_0_1),
    .I0_7_0_2(n56_I0_7_0_2),
    .I0_7_1_0(n56_I0_7_1_0),
    .I0_7_1_1(n56_I0_7_1_1),
    .I0_7_1_2(n56_I0_7_1_2),
    .I0_8_0_0(n56_I0_8_0_0),
    .I0_8_0_1(n56_I0_8_0_1),
    .I0_8_0_2(n56_I0_8_0_2),
    .I0_8_1_0(n56_I0_8_1_0),
    .I0_8_1_1(n56_I0_8_1_1),
    .I0_8_1_2(n56_I0_8_1_2),
    .I0_9_0_0(n56_I0_9_0_0),
    .I0_9_0_1(n56_I0_9_0_1),
    .I0_9_0_2(n56_I0_9_0_2),
    .I0_9_1_0(n56_I0_9_1_0),
    .I0_9_1_1(n56_I0_9_1_1),
    .I0_9_1_2(n56_I0_9_1_2),
    .I0_10_0_0(n56_I0_10_0_0),
    .I0_10_0_1(n56_I0_10_0_1),
    .I0_10_0_2(n56_I0_10_0_2),
    .I0_10_1_0(n56_I0_10_1_0),
    .I0_10_1_1(n56_I0_10_1_1),
    .I0_10_1_2(n56_I0_10_1_2),
    .I0_11_0_0(n56_I0_11_0_0),
    .I0_11_0_1(n56_I0_11_0_1),
    .I0_11_0_2(n56_I0_11_0_2),
    .I0_11_1_0(n56_I0_11_1_0),
    .I0_11_1_1(n56_I0_11_1_1),
    .I0_11_1_2(n56_I0_11_1_2),
    .I0_12_0_0(n56_I0_12_0_0),
    .I0_12_0_1(n56_I0_12_0_1),
    .I0_12_0_2(n56_I0_12_0_2),
    .I0_12_1_0(n56_I0_12_1_0),
    .I0_12_1_1(n56_I0_12_1_1),
    .I0_12_1_2(n56_I0_12_1_2),
    .I0_13_0_0(n56_I0_13_0_0),
    .I0_13_0_1(n56_I0_13_0_1),
    .I0_13_0_2(n56_I0_13_0_2),
    .I0_13_1_0(n56_I0_13_1_0),
    .I0_13_1_1(n56_I0_13_1_1),
    .I0_13_1_2(n56_I0_13_1_2),
    .I0_14_0_0(n56_I0_14_0_0),
    .I0_14_0_1(n56_I0_14_0_1),
    .I0_14_0_2(n56_I0_14_0_2),
    .I0_14_1_0(n56_I0_14_1_0),
    .I0_14_1_1(n56_I0_14_1_1),
    .I0_14_1_2(n56_I0_14_1_2),
    .I0_15_0_0(n56_I0_15_0_0),
    .I0_15_0_1(n56_I0_15_0_1),
    .I0_15_0_2(n56_I0_15_0_2),
    .I0_15_1_0(n56_I0_15_1_0),
    .I0_15_1_1(n56_I0_15_1_1),
    .I0_15_1_2(n56_I0_15_1_2),
    .I1_0_0(n56_I1_0_0),
    .I1_0_1(n56_I1_0_1),
    .I1_0_2(n56_I1_0_2),
    .I1_1_0(n56_I1_1_0),
    .I1_1_1(n56_I1_1_1),
    .I1_1_2(n56_I1_1_2),
    .I1_2_0(n56_I1_2_0),
    .I1_2_1(n56_I1_2_1),
    .I1_2_2(n56_I1_2_2),
    .I1_3_0(n56_I1_3_0),
    .I1_3_1(n56_I1_3_1),
    .I1_3_2(n56_I1_3_2),
    .I1_4_0(n56_I1_4_0),
    .I1_4_1(n56_I1_4_1),
    .I1_4_2(n56_I1_4_2),
    .I1_5_0(n56_I1_5_0),
    .I1_5_1(n56_I1_5_1),
    .I1_5_2(n56_I1_5_2),
    .I1_6_0(n56_I1_6_0),
    .I1_6_1(n56_I1_6_1),
    .I1_6_2(n56_I1_6_2),
    .I1_7_0(n56_I1_7_0),
    .I1_7_1(n56_I1_7_1),
    .I1_7_2(n56_I1_7_2),
    .I1_8_0(n56_I1_8_0),
    .I1_8_1(n56_I1_8_1),
    .I1_8_2(n56_I1_8_2),
    .I1_9_0(n56_I1_9_0),
    .I1_9_1(n56_I1_9_1),
    .I1_9_2(n56_I1_9_2),
    .I1_10_0(n56_I1_10_0),
    .I1_10_1(n56_I1_10_1),
    .I1_10_2(n56_I1_10_2),
    .I1_11_0(n56_I1_11_0),
    .I1_11_1(n56_I1_11_1),
    .I1_11_2(n56_I1_11_2),
    .I1_12_0(n56_I1_12_0),
    .I1_12_1(n56_I1_12_1),
    .I1_12_2(n56_I1_12_2),
    .I1_13_0(n56_I1_13_0),
    .I1_13_1(n56_I1_13_1),
    .I1_13_2(n56_I1_13_2),
    .I1_14_0(n56_I1_14_0),
    .I1_14_1(n56_I1_14_1),
    .I1_14_2(n56_I1_14_2),
    .I1_15_0(n56_I1_15_0),
    .I1_15_1(n56_I1_15_1),
    .I1_15_2(n56_I1_15_2),
    .O_0_0_0(n56_O_0_0_0),
    .O_0_0_1(n56_O_0_0_1),
    .O_0_0_2(n56_O_0_0_2),
    .O_0_1_0(n56_O_0_1_0),
    .O_0_1_1(n56_O_0_1_1),
    .O_0_1_2(n56_O_0_1_2),
    .O_0_2_0(n56_O_0_2_0),
    .O_0_2_1(n56_O_0_2_1),
    .O_0_2_2(n56_O_0_2_2),
    .O_1_0_0(n56_O_1_0_0),
    .O_1_0_1(n56_O_1_0_1),
    .O_1_0_2(n56_O_1_0_2),
    .O_1_1_0(n56_O_1_1_0),
    .O_1_1_1(n56_O_1_1_1),
    .O_1_1_2(n56_O_1_1_2),
    .O_1_2_0(n56_O_1_2_0),
    .O_1_2_1(n56_O_1_2_1),
    .O_1_2_2(n56_O_1_2_2),
    .O_2_0_0(n56_O_2_0_0),
    .O_2_0_1(n56_O_2_0_1),
    .O_2_0_2(n56_O_2_0_2),
    .O_2_1_0(n56_O_2_1_0),
    .O_2_1_1(n56_O_2_1_1),
    .O_2_1_2(n56_O_2_1_2),
    .O_2_2_0(n56_O_2_2_0),
    .O_2_2_1(n56_O_2_2_1),
    .O_2_2_2(n56_O_2_2_2),
    .O_3_0_0(n56_O_3_0_0),
    .O_3_0_1(n56_O_3_0_1),
    .O_3_0_2(n56_O_3_0_2),
    .O_3_1_0(n56_O_3_1_0),
    .O_3_1_1(n56_O_3_1_1),
    .O_3_1_2(n56_O_3_1_2),
    .O_3_2_0(n56_O_3_2_0),
    .O_3_2_1(n56_O_3_2_1),
    .O_3_2_2(n56_O_3_2_2),
    .O_4_0_0(n56_O_4_0_0),
    .O_4_0_1(n56_O_4_0_1),
    .O_4_0_2(n56_O_4_0_2),
    .O_4_1_0(n56_O_4_1_0),
    .O_4_1_1(n56_O_4_1_1),
    .O_4_1_2(n56_O_4_1_2),
    .O_4_2_0(n56_O_4_2_0),
    .O_4_2_1(n56_O_4_2_1),
    .O_4_2_2(n56_O_4_2_2),
    .O_5_0_0(n56_O_5_0_0),
    .O_5_0_1(n56_O_5_0_1),
    .O_5_0_2(n56_O_5_0_2),
    .O_5_1_0(n56_O_5_1_0),
    .O_5_1_1(n56_O_5_1_1),
    .O_5_1_2(n56_O_5_1_2),
    .O_5_2_0(n56_O_5_2_0),
    .O_5_2_1(n56_O_5_2_1),
    .O_5_2_2(n56_O_5_2_2),
    .O_6_0_0(n56_O_6_0_0),
    .O_6_0_1(n56_O_6_0_1),
    .O_6_0_2(n56_O_6_0_2),
    .O_6_1_0(n56_O_6_1_0),
    .O_6_1_1(n56_O_6_1_1),
    .O_6_1_2(n56_O_6_1_2),
    .O_6_2_0(n56_O_6_2_0),
    .O_6_2_1(n56_O_6_2_1),
    .O_6_2_2(n56_O_6_2_2),
    .O_7_0_0(n56_O_7_0_0),
    .O_7_0_1(n56_O_7_0_1),
    .O_7_0_2(n56_O_7_0_2),
    .O_7_1_0(n56_O_7_1_0),
    .O_7_1_1(n56_O_7_1_1),
    .O_7_1_2(n56_O_7_1_2),
    .O_7_2_0(n56_O_7_2_0),
    .O_7_2_1(n56_O_7_2_1),
    .O_7_2_2(n56_O_7_2_2),
    .O_8_0_0(n56_O_8_0_0),
    .O_8_0_1(n56_O_8_0_1),
    .O_8_0_2(n56_O_8_0_2),
    .O_8_1_0(n56_O_8_1_0),
    .O_8_1_1(n56_O_8_1_1),
    .O_8_1_2(n56_O_8_1_2),
    .O_8_2_0(n56_O_8_2_0),
    .O_8_2_1(n56_O_8_2_1),
    .O_8_2_2(n56_O_8_2_2),
    .O_9_0_0(n56_O_9_0_0),
    .O_9_0_1(n56_O_9_0_1),
    .O_9_0_2(n56_O_9_0_2),
    .O_9_1_0(n56_O_9_1_0),
    .O_9_1_1(n56_O_9_1_1),
    .O_9_1_2(n56_O_9_1_2),
    .O_9_2_0(n56_O_9_2_0),
    .O_9_2_1(n56_O_9_2_1),
    .O_9_2_2(n56_O_9_2_2),
    .O_10_0_0(n56_O_10_0_0),
    .O_10_0_1(n56_O_10_0_1),
    .O_10_0_2(n56_O_10_0_2),
    .O_10_1_0(n56_O_10_1_0),
    .O_10_1_1(n56_O_10_1_1),
    .O_10_1_2(n56_O_10_1_2),
    .O_10_2_0(n56_O_10_2_0),
    .O_10_2_1(n56_O_10_2_1),
    .O_10_2_2(n56_O_10_2_2),
    .O_11_0_0(n56_O_11_0_0),
    .O_11_0_1(n56_O_11_0_1),
    .O_11_0_2(n56_O_11_0_2),
    .O_11_1_0(n56_O_11_1_0),
    .O_11_1_1(n56_O_11_1_1),
    .O_11_1_2(n56_O_11_1_2),
    .O_11_2_0(n56_O_11_2_0),
    .O_11_2_1(n56_O_11_2_1),
    .O_11_2_2(n56_O_11_2_2),
    .O_12_0_0(n56_O_12_0_0),
    .O_12_0_1(n56_O_12_0_1),
    .O_12_0_2(n56_O_12_0_2),
    .O_12_1_0(n56_O_12_1_0),
    .O_12_1_1(n56_O_12_1_1),
    .O_12_1_2(n56_O_12_1_2),
    .O_12_2_0(n56_O_12_2_0),
    .O_12_2_1(n56_O_12_2_1),
    .O_12_2_2(n56_O_12_2_2),
    .O_13_0_0(n56_O_13_0_0),
    .O_13_0_1(n56_O_13_0_1),
    .O_13_0_2(n56_O_13_0_2),
    .O_13_1_0(n56_O_13_1_0),
    .O_13_1_1(n56_O_13_1_1),
    .O_13_1_2(n56_O_13_1_2),
    .O_13_2_0(n56_O_13_2_0),
    .O_13_2_1(n56_O_13_2_1),
    .O_13_2_2(n56_O_13_2_2),
    .O_14_0_0(n56_O_14_0_0),
    .O_14_0_1(n56_O_14_0_1),
    .O_14_0_2(n56_O_14_0_2),
    .O_14_1_0(n56_O_14_1_0),
    .O_14_1_1(n56_O_14_1_1),
    .O_14_1_2(n56_O_14_1_2),
    .O_14_2_0(n56_O_14_2_0),
    .O_14_2_1(n56_O_14_2_1),
    .O_14_2_2(n56_O_14_2_2),
    .O_15_0_0(n56_O_15_0_0),
    .O_15_0_1(n56_O_15_0_1),
    .O_15_0_2(n56_O_15_0_2),
    .O_15_1_0(n56_O_15_1_0),
    .O_15_1_1(n56_O_15_1_1),
    .O_15_1_2(n56_O_15_1_2),
    .O_15_2_0(n56_O_15_2_0),
    .O_15_2_1(n56_O_15_2_1),
    .O_15_2_2(n56_O_15_2_2)
  );
  PartitionS_3 n60 ( // @[Top.scala 193:21]
    .valid_up(n60_valid_up),
    .valid_down(n60_valid_down),
    .I_0_0_0(n60_I_0_0_0),
    .I_0_0_1(n60_I_0_0_1),
    .I_0_0_2(n60_I_0_0_2),
    .I_0_1_0(n60_I_0_1_0),
    .I_0_1_1(n60_I_0_1_1),
    .I_0_1_2(n60_I_0_1_2),
    .I_0_2_0(n60_I_0_2_0),
    .I_0_2_1(n60_I_0_2_1),
    .I_0_2_2(n60_I_0_2_2),
    .I_1_0_0(n60_I_1_0_0),
    .I_1_0_1(n60_I_1_0_1),
    .I_1_0_2(n60_I_1_0_2),
    .I_1_1_0(n60_I_1_1_0),
    .I_1_1_1(n60_I_1_1_1),
    .I_1_1_2(n60_I_1_1_2),
    .I_1_2_0(n60_I_1_2_0),
    .I_1_2_1(n60_I_1_2_1),
    .I_1_2_2(n60_I_1_2_2),
    .I_2_0_0(n60_I_2_0_0),
    .I_2_0_1(n60_I_2_0_1),
    .I_2_0_2(n60_I_2_0_2),
    .I_2_1_0(n60_I_2_1_0),
    .I_2_1_1(n60_I_2_1_1),
    .I_2_1_2(n60_I_2_1_2),
    .I_2_2_0(n60_I_2_2_0),
    .I_2_2_1(n60_I_2_2_1),
    .I_2_2_2(n60_I_2_2_2),
    .I_3_0_0(n60_I_3_0_0),
    .I_3_0_1(n60_I_3_0_1),
    .I_3_0_2(n60_I_3_0_2),
    .I_3_1_0(n60_I_3_1_0),
    .I_3_1_1(n60_I_3_1_1),
    .I_3_1_2(n60_I_3_1_2),
    .I_3_2_0(n60_I_3_2_0),
    .I_3_2_1(n60_I_3_2_1),
    .I_3_2_2(n60_I_3_2_2),
    .I_4_0_0(n60_I_4_0_0),
    .I_4_0_1(n60_I_4_0_1),
    .I_4_0_2(n60_I_4_0_2),
    .I_4_1_0(n60_I_4_1_0),
    .I_4_1_1(n60_I_4_1_1),
    .I_4_1_2(n60_I_4_1_2),
    .I_4_2_0(n60_I_4_2_0),
    .I_4_2_1(n60_I_4_2_1),
    .I_4_2_2(n60_I_4_2_2),
    .I_5_0_0(n60_I_5_0_0),
    .I_5_0_1(n60_I_5_0_1),
    .I_5_0_2(n60_I_5_0_2),
    .I_5_1_0(n60_I_5_1_0),
    .I_5_1_1(n60_I_5_1_1),
    .I_5_1_2(n60_I_5_1_2),
    .I_5_2_0(n60_I_5_2_0),
    .I_5_2_1(n60_I_5_2_1),
    .I_5_2_2(n60_I_5_2_2),
    .I_6_0_0(n60_I_6_0_0),
    .I_6_0_1(n60_I_6_0_1),
    .I_6_0_2(n60_I_6_0_2),
    .I_6_1_0(n60_I_6_1_0),
    .I_6_1_1(n60_I_6_1_1),
    .I_6_1_2(n60_I_6_1_2),
    .I_6_2_0(n60_I_6_2_0),
    .I_6_2_1(n60_I_6_2_1),
    .I_6_2_2(n60_I_6_2_2),
    .I_7_0_0(n60_I_7_0_0),
    .I_7_0_1(n60_I_7_0_1),
    .I_7_0_2(n60_I_7_0_2),
    .I_7_1_0(n60_I_7_1_0),
    .I_7_1_1(n60_I_7_1_1),
    .I_7_1_2(n60_I_7_1_2),
    .I_7_2_0(n60_I_7_2_0),
    .I_7_2_1(n60_I_7_2_1),
    .I_7_2_2(n60_I_7_2_2),
    .I_8_0_0(n60_I_8_0_0),
    .I_8_0_1(n60_I_8_0_1),
    .I_8_0_2(n60_I_8_0_2),
    .I_8_1_0(n60_I_8_1_0),
    .I_8_1_1(n60_I_8_1_1),
    .I_8_1_2(n60_I_8_1_2),
    .I_8_2_0(n60_I_8_2_0),
    .I_8_2_1(n60_I_8_2_1),
    .I_8_2_2(n60_I_8_2_2),
    .I_9_0_0(n60_I_9_0_0),
    .I_9_0_1(n60_I_9_0_1),
    .I_9_0_2(n60_I_9_0_2),
    .I_9_1_0(n60_I_9_1_0),
    .I_9_1_1(n60_I_9_1_1),
    .I_9_1_2(n60_I_9_1_2),
    .I_9_2_0(n60_I_9_2_0),
    .I_9_2_1(n60_I_9_2_1),
    .I_9_2_2(n60_I_9_2_2),
    .I_10_0_0(n60_I_10_0_0),
    .I_10_0_1(n60_I_10_0_1),
    .I_10_0_2(n60_I_10_0_2),
    .I_10_1_0(n60_I_10_1_0),
    .I_10_1_1(n60_I_10_1_1),
    .I_10_1_2(n60_I_10_1_2),
    .I_10_2_0(n60_I_10_2_0),
    .I_10_2_1(n60_I_10_2_1),
    .I_10_2_2(n60_I_10_2_2),
    .I_11_0_0(n60_I_11_0_0),
    .I_11_0_1(n60_I_11_0_1),
    .I_11_0_2(n60_I_11_0_2),
    .I_11_1_0(n60_I_11_1_0),
    .I_11_1_1(n60_I_11_1_1),
    .I_11_1_2(n60_I_11_1_2),
    .I_11_2_0(n60_I_11_2_0),
    .I_11_2_1(n60_I_11_2_1),
    .I_11_2_2(n60_I_11_2_2),
    .I_12_0_0(n60_I_12_0_0),
    .I_12_0_1(n60_I_12_0_1),
    .I_12_0_2(n60_I_12_0_2),
    .I_12_1_0(n60_I_12_1_0),
    .I_12_1_1(n60_I_12_1_1),
    .I_12_1_2(n60_I_12_1_2),
    .I_12_2_0(n60_I_12_2_0),
    .I_12_2_1(n60_I_12_2_1),
    .I_12_2_2(n60_I_12_2_2),
    .I_13_0_0(n60_I_13_0_0),
    .I_13_0_1(n60_I_13_0_1),
    .I_13_0_2(n60_I_13_0_2),
    .I_13_1_0(n60_I_13_1_0),
    .I_13_1_1(n60_I_13_1_1),
    .I_13_1_2(n60_I_13_1_2),
    .I_13_2_0(n60_I_13_2_0),
    .I_13_2_1(n60_I_13_2_1),
    .I_13_2_2(n60_I_13_2_2),
    .I_14_0_0(n60_I_14_0_0),
    .I_14_0_1(n60_I_14_0_1),
    .I_14_0_2(n60_I_14_0_2),
    .I_14_1_0(n60_I_14_1_0),
    .I_14_1_1(n60_I_14_1_1),
    .I_14_1_2(n60_I_14_1_2),
    .I_14_2_0(n60_I_14_2_0),
    .I_14_2_1(n60_I_14_2_1),
    .I_14_2_2(n60_I_14_2_2),
    .I_15_0_0(n60_I_15_0_0),
    .I_15_0_1(n60_I_15_0_1),
    .I_15_0_2(n60_I_15_0_2),
    .I_15_1_0(n60_I_15_1_0),
    .I_15_1_1(n60_I_15_1_1),
    .I_15_1_2(n60_I_15_1_2),
    .I_15_2_0(n60_I_15_2_0),
    .I_15_2_1(n60_I_15_2_1),
    .I_15_2_2(n60_I_15_2_2),
    .O_0_0_0_0(n60_O_0_0_0_0),
    .O_0_0_0_1(n60_O_0_0_0_1),
    .O_0_0_0_2(n60_O_0_0_0_2),
    .O_0_0_1_0(n60_O_0_0_1_0),
    .O_0_0_1_1(n60_O_0_0_1_1),
    .O_0_0_1_2(n60_O_0_0_1_2),
    .O_0_0_2_0(n60_O_0_0_2_0),
    .O_0_0_2_1(n60_O_0_0_2_1),
    .O_0_0_2_2(n60_O_0_0_2_2),
    .O_1_0_0_0(n60_O_1_0_0_0),
    .O_1_0_0_1(n60_O_1_0_0_1),
    .O_1_0_0_2(n60_O_1_0_0_2),
    .O_1_0_1_0(n60_O_1_0_1_0),
    .O_1_0_1_1(n60_O_1_0_1_1),
    .O_1_0_1_2(n60_O_1_0_1_2),
    .O_1_0_2_0(n60_O_1_0_2_0),
    .O_1_0_2_1(n60_O_1_0_2_1),
    .O_1_0_2_2(n60_O_1_0_2_2),
    .O_2_0_0_0(n60_O_2_0_0_0),
    .O_2_0_0_1(n60_O_2_0_0_1),
    .O_2_0_0_2(n60_O_2_0_0_2),
    .O_2_0_1_0(n60_O_2_0_1_0),
    .O_2_0_1_1(n60_O_2_0_1_1),
    .O_2_0_1_2(n60_O_2_0_1_2),
    .O_2_0_2_0(n60_O_2_0_2_0),
    .O_2_0_2_1(n60_O_2_0_2_1),
    .O_2_0_2_2(n60_O_2_0_2_2),
    .O_3_0_0_0(n60_O_3_0_0_0),
    .O_3_0_0_1(n60_O_3_0_0_1),
    .O_3_0_0_2(n60_O_3_0_0_2),
    .O_3_0_1_0(n60_O_3_0_1_0),
    .O_3_0_1_1(n60_O_3_0_1_1),
    .O_3_0_1_2(n60_O_3_0_1_2),
    .O_3_0_2_0(n60_O_3_0_2_0),
    .O_3_0_2_1(n60_O_3_0_2_1),
    .O_3_0_2_2(n60_O_3_0_2_2),
    .O_4_0_0_0(n60_O_4_0_0_0),
    .O_4_0_0_1(n60_O_4_0_0_1),
    .O_4_0_0_2(n60_O_4_0_0_2),
    .O_4_0_1_0(n60_O_4_0_1_0),
    .O_4_0_1_1(n60_O_4_0_1_1),
    .O_4_0_1_2(n60_O_4_0_1_2),
    .O_4_0_2_0(n60_O_4_0_2_0),
    .O_4_0_2_1(n60_O_4_0_2_1),
    .O_4_0_2_2(n60_O_4_0_2_2),
    .O_5_0_0_0(n60_O_5_0_0_0),
    .O_5_0_0_1(n60_O_5_0_0_1),
    .O_5_0_0_2(n60_O_5_0_0_2),
    .O_5_0_1_0(n60_O_5_0_1_0),
    .O_5_0_1_1(n60_O_5_0_1_1),
    .O_5_0_1_2(n60_O_5_0_1_2),
    .O_5_0_2_0(n60_O_5_0_2_0),
    .O_5_0_2_1(n60_O_5_0_2_1),
    .O_5_0_2_2(n60_O_5_0_2_2),
    .O_6_0_0_0(n60_O_6_0_0_0),
    .O_6_0_0_1(n60_O_6_0_0_1),
    .O_6_0_0_2(n60_O_6_0_0_2),
    .O_6_0_1_0(n60_O_6_0_1_0),
    .O_6_0_1_1(n60_O_6_0_1_1),
    .O_6_0_1_2(n60_O_6_0_1_2),
    .O_6_0_2_0(n60_O_6_0_2_0),
    .O_6_0_2_1(n60_O_6_0_2_1),
    .O_6_0_2_2(n60_O_6_0_2_2),
    .O_7_0_0_0(n60_O_7_0_0_0),
    .O_7_0_0_1(n60_O_7_0_0_1),
    .O_7_0_0_2(n60_O_7_0_0_2),
    .O_7_0_1_0(n60_O_7_0_1_0),
    .O_7_0_1_1(n60_O_7_0_1_1),
    .O_7_0_1_2(n60_O_7_0_1_2),
    .O_7_0_2_0(n60_O_7_0_2_0),
    .O_7_0_2_1(n60_O_7_0_2_1),
    .O_7_0_2_2(n60_O_7_0_2_2),
    .O_8_0_0_0(n60_O_8_0_0_0),
    .O_8_0_0_1(n60_O_8_0_0_1),
    .O_8_0_0_2(n60_O_8_0_0_2),
    .O_8_0_1_0(n60_O_8_0_1_0),
    .O_8_0_1_1(n60_O_8_0_1_1),
    .O_8_0_1_2(n60_O_8_0_1_2),
    .O_8_0_2_0(n60_O_8_0_2_0),
    .O_8_0_2_1(n60_O_8_0_2_1),
    .O_8_0_2_2(n60_O_8_0_2_2),
    .O_9_0_0_0(n60_O_9_0_0_0),
    .O_9_0_0_1(n60_O_9_0_0_1),
    .O_9_0_0_2(n60_O_9_0_0_2),
    .O_9_0_1_0(n60_O_9_0_1_0),
    .O_9_0_1_1(n60_O_9_0_1_1),
    .O_9_0_1_2(n60_O_9_0_1_2),
    .O_9_0_2_0(n60_O_9_0_2_0),
    .O_9_0_2_1(n60_O_9_0_2_1),
    .O_9_0_2_2(n60_O_9_0_2_2),
    .O_10_0_0_0(n60_O_10_0_0_0),
    .O_10_0_0_1(n60_O_10_0_0_1),
    .O_10_0_0_2(n60_O_10_0_0_2),
    .O_10_0_1_0(n60_O_10_0_1_0),
    .O_10_0_1_1(n60_O_10_0_1_1),
    .O_10_0_1_2(n60_O_10_0_1_2),
    .O_10_0_2_0(n60_O_10_0_2_0),
    .O_10_0_2_1(n60_O_10_0_2_1),
    .O_10_0_2_2(n60_O_10_0_2_2),
    .O_11_0_0_0(n60_O_11_0_0_0),
    .O_11_0_0_1(n60_O_11_0_0_1),
    .O_11_0_0_2(n60_O_11_0_0_2),
    .O_11_0_1_0(n60_O_11_0_1_0),
    .O_11_0_1_1(n60_O_11_0_1_1),
    .O_11_0_1_2(n60_O_11_0_1_2),
    .O_11_0_2_0(n60_O_11_0_2_0),
    .O_11_0_2_1(n60_O_11_0_2_1),
    .O_11_0_2_2(n60_O_11_0_2_2),
    .O_12_0_0_0(n60_O_12_0_0_0),
    .O_12_0_0_1(n60_O_12_0_0_1),
    .O_12_0_0_2(n60_O_12_0_0_2),
    .O_12_0_1_0(n60_O_12_0_1_0),
    .O_12_0_1_1(n60_O_12_0_1_1),
    .O_12_0_1_2(n60_O_12_0_1_2),
    .O_12_0_2_0(n60_O_12_0_2_0),
    .O_12_0_2_1(n60_O_12_0_2_1),
    .O_12_0_2_2(n60_O_12_0_2_2),
    .O_13_0_0_0(n60_O_13_0_0_0),
    .O_13_0_0_1(n60_O_13_0_0_1),
    .O_13_0_0_2(n60_O_13_0_0_2),
    .O_13_0_1_0(n60_O_13_0_1_0),
    .O_13_0_1_1(n60_O_13_0_1_1),
    .O_13_0_1_2(n60_O_13_0_1_2),
    .O_13_0_2_0(n60_O_13_0_2_0),
    .O_13_0_2_1(n60_O_13_0_2_1),
    .O_13_0_2_2(n60_O_13_0_2_2),
    .O_14_0_0_0(n60_O_14_0_0_0),
    .O_14_0_0_1(n60_O_14_0_0_1),
    .O_14_0_0_2(n60_O_14_0_0_2),
    .O_14_0_1_0(n60_O_14_0_1_0),
    .O_14_0_1_1(n60_O_14_0_1_1),
    .O_14_0_1_2(n60_O_14_0_1_2),
    .O_14_0_2_0(n60_O_14_0_2_0),
    .O_14_0_2_1(n60_O_14_0_2_1),
    .O_14_0_2_2(n60_O_14_0_2_2),
    .O_15_0_0_0(n60_O_15_0_0_0),
    .O_15_0_0_1(n60_O_15_0_0_1),
    .O_15_0_0_2(n60_O_15_0_0_2),
    .O_15_0_1_0(n60_O_15_0_1_0),
    .O_15_0_1_1(n60_O_15_0_1_1),
    .O_15_0_1_2(n60_O_15_0_1_2),
    .O_15_0_2_0(n60_O_15_0_2_0),
    .O_15_0_2_1(n60_O_15_0_2_1),
    .O_15_0_2_2(n60_O_15_0_2_2)
  );
  MapS_3 n65 ( // @[Top.scala 196:21]
    .valid_up(n65_valid_up),
    .valid_down(n65_valid_down),
    .I_0_0_0_0(n65_I_0_0_0_0),
    .I_0_0_0_1(n65_I_0_0_0_1),
    .I_0_0_0_2(n65_I_0_0_0_2),
    .I_0_0_1_0(n65_I_0_0_1_0),
    .I_0_0_1_1(n65_I_0_0_1_1),
    .I_0_0_1_2(n65_I_0_0_1_2),
    .I_0_0_2_0(n65_I_0_0_2_0),
    .I_0_0_2_1(n65_I_0_0_2_1),
    .I_0_0_2_2(n65_I_0_0_2_2),
    .I_1_0_0_0(n65_I_1_0_0_0),
    .I_1_0_0_1(n65_I_1_0_0_1),
    .I_1_0_0_2(n65_I_1_0_0_2),
    .I_1_0_1_0(n65_I_1_0_1_0),
    .I_1_0_1_1(n65_I_1_0_1_1),
    .I_1_0_1_2(n65_I_1_0_1_2),
    .I_1_0_2_0(n65_I_1_0_2_0),
    .I_1_0_2_1(n65_I_1_0_2_1),
    .I_1_0_2_2(n65_I_1_0_2_2),
    .I_2_0_0_0(n65_I_2_0_0_0),
    .I_2_0_0_1(n65_I_2_0_0_1),
    .I_2_0_0_2(n65_I_2_0_0_2),
    .I_2_0_1_0(n65_I_2_0_1_0),
    .I_2_0_1_1(n65_I_2_0_1_1),
    .I_2_0_1_2(n65_I_2_0_1_2),
    .I_2_0_2_0(n65_I_2_0_2_0),
    .I_2_0_2_1(n65_I_2_0_2_1),
    .I_2_0_2_2(n65_I_2_0_2_2),
    .I_3_0_0_0(n65_I_3_0_0_0),
    .I_3_0_0_1(n65_I_3_0_0_1),
    .I_3_0_0_2(n65_I_3_0_0_2),
    .I_3_0_1_0(n65_I_3_0_1_0),
    .I_3_0_1_1(n65_I_3_0_1_1),
    .I_3_0_1_2(n65_I_3_0_1_2),
    .I_3_0_2_0(n65_I_3_0_2_0),
    .I_3_0_2_1(n65_I_3_0_2_1),
    .I_3_0_2_2(n65_I_3_0_2_2),
    .I_4_0_0_0(n65_I_4_0_0_0),
    .I_4_0_0_1(n65_I_4_0_0_1),
    .I_4_0_0_2(n65_I_4_0_0_2),
    .I_4_0_1_0(n65_I_4_0_1_0),
    .I_4_0_1_1(n65_I_4_0_1_1),
    .I_4_0_1_2(n65_I_4_0_1_2),
    .I_4_0_2_0(n65_I_4_0_2_0),
    .I_4_0_2_1(n65_I_4_0_2_1),
    .I_4_0_2_2(n65_I_4_0_2_2),
    .I_5_0_0_0(n65_I_5_0_0_0),
    .I_5_0_0_1(n65_I_5_0_0_1),
    .I_5_0_0_2(n65_I_5_0_0_2),
    .I_5_0_1_0(n65_I_5_0_1_0),
    .I_5_0_1_1(n65_I_5_0_1_1),
    .I_5_0_1_2(n65_I_5_0_1_2),
    .I_5_0_2_0(n65_I_5_0_2_0),
    .I_5_0_2_1(n65_I_5_0_2_1),
    .I_5_0_2_2(n65_I_5_0_2_2),
    .I_6_0_0_0(n65_I_6_0_0_0),
    .I_6_0_0_1(n65_I_6_0_0_1),
    .I_6_0_0_2(n65_I_6_0_0_2),
    .I_6_0_1_0(n65_I_6_0_1_0),
    .I_6_0_1_1(n65_I_6_0_1_1),
    .I_6_0_1_2(n65_I_6_0_1_2),
    .I_6_0_2_0(n65_I_6_0_2_0),
    .I_6_0_2_1(n65_I_6_0_2_1),
    .I_6_0_2_2(n65_I_6_0_2_2),
    .I_7_0_0_0(n65_I_7_0_0_0),
    .I_7_0_0_1(n65_I_7_0_0_1),
    .I_7_0_0_2(n65_I_7_0_0_2),
    .I_7_0_1_0(n65_I_7_0_1_0),
    .I_7_0_1_1(n65_I_7_0_1_1),
    .I_7_0_1_2(n65_I_7_0_1_2),
    .I_7_0_2_0(n65_I_7_0_2_0),
    .I_7_0_2_1(n65_I_7_0_2_1),
    .I_7_0_2_2(n65_I_7_0_2_2),
    .I_8_0_0_0(n65_I_8_0_0_0),
    .I_8_0_0_1(n65_I_8_0_0_1),
    .I_8_0_0_2(n65_I_8_0_0_2),
    .I_8_0_1_0(n65_I_8_0_1_0),
    .I_8_0_1_1(n65_I_8_0_1_1),
    .I_8_0_1_2(n65_I_8_0_1_2),
    .I_8_0_2_0(n65_I_8_0_2_0),
    .I_8_0_2_1(n65_I_8_0_2_1),
    .I_8_0_2_2(n65_I_8_0_2_2),
    .I_9_0_0_0(n65_I_9_0_0_0),
    .I_9_0_0_1(n65_I_9_0_0_1),
    .I_9_0_0_2(n65_I_9_0_0_2),
    .I_9_0_1_0(n65_I_9_0_1_0),
    .I_9_0_1_1(n65_I_9_0_1_1),
    .I_9_0_1_2(n65_I_9_0_1_2),
    .I_9_0_2_0(n65_I_9_0_2_0),
    .I_9_0_2_1(n65_I_9_0_2_1),
    .I_9_0_2_2(n65_I_9_0_2_2),
    .I_10_0_0_0(n65_I_10_0_0_0),
    .I_10_0_0_1(n65_I_10_0_0_1),
    .I_10_0_0_2(n65_I_10_0_0_2),
    .I_10_0_1_0(n65_I_10_0_1_0),
    .I_10_0_1_1(n65_I_10_0_1_1),
    .I_10_0_1_2(n65_I_10_0_1_2),
    .I_10_0_2_0(n65_I_10_0_2_0),
    .I_10_0_2_1(n65_I_10_0_2_1),
    .I_10_0_2_2(n65_I_10_0_2_2),
    .I_11_0_0_0(n65_I_11_0_0_0),
    .I_11_0_0_1(n65_I_11_0_0_1),
    .I_11_0_0_2(n65_I_11_0_0_2),
    .I_11_0_1_0(n65_I_11_0_1_0),
    .I_11_0_1_1(n65_I_11_0_1_1),
    .I_11_0_1_2(n65_I_11_0_1_2),
    .I_11_0_2_0(n65_I_11_0_2_0),
    .I_11_0_2_1(n65_I_11_0_2_1),
    .I_11_0_2_2(n65_I_11_0_2_2),
    .I_12_0_0_0(n65_I_12_0_0_0),
    .I_12_0_0_1(n65_I_12_0_0_1),
    .I_12_0_0_2(n65_I_12_0_0_2),
    .I_12_0_1_0(n65_I_12_0_1_0),
    .I_12_0_1_1(n65_I_12_0_1_1),
    .I_12_0_1_2(n65_I_12_0_1_2),
    .I_12_0_2_0(n65_I_12_0_2_0),
    .I_12_0_2_1(n65_I_12_0_2_1),
    .I_12_0_2_2(n65_I_12_0_2_2),
    .I_13_0_0_0(n65_I_13_0_0_0),
    .I_13_0_0_1(n65_I_13_0_0_1),
    .I_13_0_0_2(n65_I_13_0_0_2),
    .I_13_0_1_0(n65_I_13_0_1_0),
    .I_13_0_1_1(n65_I_13_0_1_1),
    .I_13_0_1_2(n65_I_13_0_1_2),
    .I_13_0_2_0(n65_I_13_0_2_0),
    .I_13_0_2_1(n65_I_13_0_2_1),
    .I_13_0_2_2(n65_I_13_0_2_2),
    .I_14_0_0_0(n65_I_14_0_0_0),
    .I_14_0_0_1(n65_I_14_0_0_1),
    .I_14_0_0_2(n65_I_14_0_0_2),
    .I_14_0_1_0(n65_I_14_0_1_0),
    .I_14_0_1_1(n65_I_14_0_1_1),
    .I_14_0_1_2(n65_I_14_0_1_2),
    .I_14_0_2_0(n65_I_14_0_2_0),
    .I_14_0_2_1(n65_I_14_0_2_1),
    .I_14_0_2_2(n65_I_14_0_2_2),
    .I_15_0_0_0(n65_I_15_0_0_0),
    .I_15_0_0_1(n65_I_15_0_0_1),
    .I_15_0_0_2(n65_I_15_0_0_2),
    .I_15_0_1_0(n65_I_15_0_1_0),
    .I_15_0_1_1(n65_I_15_0_1_1),
    .I_15_0_1_2(n65_I_15_0_1_2),
    .I_15_0_2_0(n65_I_15_0_2_0),
    .I_15_0_2_1(n65_I_15_0_2_1),
    .I_15_0_2_2(n65_I_15_0_2_2),
    .O_0_0_0(n65_O_0_0_0),
    .O_0_0_1(n65_O_0_0_1),
    .O_0_0_2(n65_O_0_0_2),
    .O_0_1_0(n65_O_0_1_0),
    .O_0_1_1(n65_O_0_1_1),
    .O_0_1_2(n65_O_0_1_2),
    .O_0_2_0(n65_O_0_2_0),
    .O_0_2_1(n65_O_0_2_1),
    .O_0_2_2(n65_O_0_2_2),
    .O_1_0_0(n65_O_1_0_0),
    .O_1_0_1(n65_O_1_0_1),
    .O_1_0_2(n65_O_1_0_2),
    .O_1_1_0(n65_O_1_1_0),
    .O_1_1_1(n65_O_1_1_1),
    .O_1_1_2(n65_O_1_1_2),
    .O_1_2_0(n65_O_1_2_0),
    .O_1_2_1(n65_O_1_2_1),
    .O_1_2_2(n65_O_1_2_2),
    .O_2_0_0(n65_O_2_0_0),
    .O_2_0_1(n65_O_2_0_1),
    .O_2_0_2(n65_O_2_0_2),
    .O_2_1_0(n65_O_2_1_0),
    .O_2_1_1(n65_O_2_1_1),
    .O_2_1_2(n65_O_2_1_2),
    .O_2_2_0(n65_O_2_2_0),
    .O_2_2_1(n65_O_2_2_1),
    .O_2_2_2(n65_O_2_2_2),
    .O_3_0_0(n65_O_3_0_0),
    .O_3_0_1(n65_O_3_0_1),
    .O_3_0_2(n65_O_3_0_2),
    .O_3_1_0(n65_O_3_1_0),
    .O_3_1_1(n65_O_3_1_1),
    .O_3_1_2(n65_O_3_1_2),
    .O_3_2_0(n65_O_3_2_0),
    .O_3_2_1(n65_O_3_2_1),
    .O_3_2_2(n65_O_3_2_2),
    .O_4_0_0(n65_O_4_0_0),
    .O_4_0_1(n65_O_4_0_1),
    .O_4_0_2(n65_O_4_0_2),
    .O_4_1_0(n65_O_4_1_0),
    .O_4_1_1(n65_O_4_1_1),
    .O_4_1_2(n65_O_4_1_2),
    .O_4_2_0(n65_O_4_2_0),
    .O_4_2_1(n65_O_4_2_1),
    .O_4_2_2(n65_O_4_2_2),
    .O_5_0_0(n65_O_5_0_0),
    .O_5_0_1(n65_O_5_0_1),
    .O_5_0_2(n65_O_5_0_2),
    .O_5_1_0(n65_O_5_1_0),
    .O_5_1_1(n65_O_5_1_1),
    .O_5_1_2(n65_O_5_1_2),
    .O_5_2_0(n65_O_5_2_0),
    .O_5_2_1(n65_O_5_2_1),
    .O_5_2_2(n65_O_5_2_2),
    .O_6_0_0(n65_O_6_0_0),
    .O_6_0_1(n65_O_6_0_1),
    .O_6_0_2(n65_O_6_0_2),
    .O_6_1_0(n65_O_6_1_0),
    .O_6_1_1(n65_O_6_1_1),
    .O_6_1_2(n65_O_6_1_2),
    .O_6_2_0(n65_O_6_2_0),
    .O_6_2_1(n65_O_6_2_1),
    .O_6_2_2(n65_O_6_2_2),
    .O_7_0_0(n65_O_7_0_0),
    .O_7_0_1(n65_O_7_0_1),
    .O_7_0_2(n65_O_7_0_2),
    .O_7_1_0(n65_O_7_1_0),
    .O_7_1_1(n65_O_7_1_1),
    .O_7_1_2(n65_O_7_1_2),
    .O_7_2_0(n65_O_7_2_0),
    .O_7_2_1(n65_O_7_2_1),
    .O_7_2_2(n65_O_7_2_2),
    .O_8_0_0(n65_O_8_0_0),
    .O_8_0_1(n65_O_8_0_1),
    .O_8_0_2(n65_O_8_0_2),
    .O_8_1_0(n65_O_8_1_0),
    .O_8_1_1(n65_O_8_1_1),
    .O_8_1_2(n65_O_8_1_2),
    .O_8_2_0(n65_O_8_2_0),
    .O_8_2_1(n65_O_8_2_1),
    .O_8_2_2(n65_O_8_2_2),
    .O_9_0_0(n65_O_9_0_0),
    .O_9_0_1(n65_O_9_0_1),
    .O_9_0_2(n65_O_9_0_2),
    .O_9_1_0(n65_O_9_1_0),
    .O_9_1_1(n65_O_9_1_1),
    .O_9_1_2(n65_O_9_1_2),
    .O_9_2_0(n65_O_9_2_0),
    .O_9_2_1(n65_O_9_2_1),
    .O_9_2_2(n65_O_9_2_2),
    .O_10_0_0(n65_O_10_0_0),
    .O_10_0_1(n65_O_10_0_1),
    .O_10_0_2(n65_O_10_0_2),
    .O_10_1_0(n65_O_10_1_0),
    .O_10_1_1(n65_O_10_1_1),
    .O_10_1_2(n65_O_10_1_2),
    .O_10_2_0(n65_O_10_2_0),
    .O_10_2_1(n65_O_10_2_1),
    .O_10_2_2(n65_O_10_2_2),
    .O_11_0_0(n65_O_11_0_0),
    .O_11_0_1(n65_O_11_0_1),
    .O_11_0_2(n65_O_11_0_2),
    .O_11_1_0(n65_O_11_1_0),
    .O_11_1_1(n65_O_11_1_1),
    .O_11_1_2(n65_O_11_1_2),
    .O_11_2_0(n65_O_11_2_0),
    .O_11_2_1(n65_O_11_2_1),
    .O_11_2_2(n65_O_11_2_2),
    .O_12_0_0(n65_O_12_0_0),
    .O_12_0_1(n65_O_12_0_1),
    .O_12_0_2(n65_O_12_0_2),
    .O_12_1_0(n65_O_12_1_0),
    .O_12_1_1(n65_O_12_1_1),
    .O_12_1_2(n65_O_12_1_2),
    .O_12_2_0(n65_O_12_2_0),
    .O_12_2_1(n65_O_12_2_1),
    .O_12_2_2(n65_O_12_2_2),
    .O_13_0_0(n65_O_13_0_0),
    .O_13_0_1(n65_O_13_0_1),
    .O_13_0_2(n65_O_13_0_2),
    .O_13_1_0(n65_O_13_1_0),
    .O_13_1_1(n65_O_13_1_1),
    .O_13_1_2(n65_O_13_1_2),
    .O_13_2_0(n65_O_13_2_0),
    .O_13_2_1(n65_O_13_2_1),
    .O_13_2_2(n65_O_13_2_2),
    .O_14_0_0(n65_O_14_0_0),
    .O_14_0_1(n65_O_14_0_1),
    .O_14_0_2(n65_O_14_0_2),
    .O_14_1_0(n65_O_14_1_0),
    .O_14_1_1(n65_O_14_1_1),
    .O_14_1_2(n65_O_14_1_2),
    .O_14_2_0(n65_O_14_2_0),
    .O_14_2_1(n65_O_14_2_1),
    .O_14_2_2(n65_O_14_2_2),
    .O_15_0_0(n65_O_15_0_0),
    .O_15_0_1(n65_O_15_0_1),
    .O_15_0_2(n65_O_15_0_2),
    .O_15_1_0(n65_O_15_1_0),
    .O_15_1_1(n65_O_15_1_1),
    .O_15_1_2(n65_O_15_1_2),
    .O_15_2_0(n65_O_15_2_0),
    .O_15_2_1(n65_O_15_2_1),
    .O_15_2_2(n65_O_15_2_2)
  );
  MapS_9 n105 ( // @[Top.scala 199:22]
    .clock(n105_clock),
    .reset(n105_reset),
    .valid_up(n105_valid_up),
    .valid_down(n105_valid_down),
    .I_0_0_0(n105_I_0_0_0),
    .I_0_0_1(n105_I_0_0_1),
    .I_0_0_2(n105_I_0_0_2),
    .I_0_1_0(n105_I_0_1_0),
    .I_0_1_1(n105_I_0_1_1),
    .I_0_1_2(n105_I_0_1_2),
    .I_0_2_0(n105_I_0_2_0),
    .I_0_2_1(n105_I_0_2_1),
    .I_0_2_2(n105_I_0_2_2),
    .I_1_0_0(n105_I_1_0_0),
    .I_1_0_1(n105_I_1_0_1),
    .I_1_0_2(n105_I_1_0_2),
    .I_1_1_0(n105_I_1_1_0),
    .I_1_1_1(n105_I_1_1_1),
    .I_1_1_2(n105_I_1_1_2),
    .I_1_2_0(n105_I_1_2_0),
    .I_1_2_1(n105_I_1_2_1),
    .I_1_2_2(n105_I_1_2_2),
    .I_2_0_0(n105_I_2_0_0),
    .I_2_0_1(n105_I_2_0_1),
    .I_2_0_2(n105_I_2_0_2),
    .I_2_1_0(n105_I_2_1_0),
    .I_2_1_1(n105_I_2_1_1),
    .I_2_1_2(n105_I_2_1_2),
    .I_2_2_0(n105_I_2_2_0),
    .I_2_2_1(n105_I_2_2_1),
    .I_2_2_2(n105_I_2_2_2),
    .I_3_0_0(n105_I_3_0_0),
    .I_3_0_1(n105_I_3_0_1),
    .I_3_0_2(n105_I_3_0_2),
    .I_3_1_0(n105_I_3_1_0),
    .I_3_1_1(n105_I_3_1_1),
    .I_3_1_2(n105_I_3_1_2),
    .I_3_2_0(n105_I_3_2_0),
    .I_3_2_1(n105_I_3_2_1),
    .I_3_2_2(n105_I_3_2_2),
    .I_4_0_0(n105_I_4_0_0),
    .I_4_0_1(n105_I_4_0_1),
    .I_4_0_2(n105_I_4_0_2),
    .I_4_1_0(n105_I_4_1_0),
    .I_4_1_1(n105_I_4_1_1),
    .I_4_1_2(n105_I_4_1_2),
    .I_4_2_0(n105_I_4_2_0),
    .I_4_2_1(n105_I_4_2_1),
    .I_4_2_2(n105_I_4_2_2),
    .I_5_0_0(n105_I_5_0_0),
    .I_5_0_1(n105_I_5_0_1),
    .I_5_0_2(n105_I_5_0_2),
    .I_5_1_0(n105_I_5_1_0),
    .I_5_1_1(n105_I_5_1_1),
    .I_5_1_2(n105_I_5_1_2),
    .I_5_2_0(n105_I_5_2_0),
    .I_5_2_1(n105_I_5_2_1),
    .I_5_2_2(n105_I_5_2_2),
    .I_6_0_0(n105_I_6_0_0),
    .I_6_0_1(n105_I_6_0_1),
    .I_6_0_2(n105_I_6_0_2),
    .I_6_1_0(n105_I_6_1_0),
    .I_6_1_1(n105_I_6_1_1),
    .I_6_1_2(n105_I_6_1_2),
    .I_6_2_0(n105_I_6_2_0),
    .I_6_2_1(n105_I_6_2_1),
    .I_6_2_2(n105_I_6_2_2),
    .I_7_0_0(n105_I_7_0_0),
    .I_7_0_1(n105_I_7_0_1),
    .I_7_0_2(n105_I_7_0_2),
    .I_7_1_0(n105_I_7_1_0),
    .I_7_1_1(n105_I_7_1_1),
    .I_7_1_2(n105_I_7_1_2),
    .I_7_2_0(n105_I_7_2_0),
    .I_7_2_1(n105_I_7_2_1),
    .I_7_2_2(n105_I_7_2_2),
    .I_8_0_0(n105_I_8_0_0),
    .I_8_0_1(n105_I_8_0_1),
    .I_8_0_2(n105_I_8_0_2),
    .I_8_1_0(n105_I_8_1_0),
    .I_8_1_1(n105_I_8_1_1),
    .I_8_1_2(n105_I_8_1_2),
    .I_8_2_0(n105_I_8_2_0),
    .I_8_2_1(n105_I_8_2_1),
    .I_8_2_2(n105_I_8_2_2),
    .I_9_0_0(n105_I_9_0_0),
    .I_9_0_1(n105_I_9_0_1),
    .I_9_0_2(n105_I_9_0_2),
    .I_9_1_0(n105_I_9_1_0),
    .I_9_1_1(n105_I_9_1_1),
    .I_9_1_2(n105_I_9_1_2),
    .I_9_2_0(n105_I_9_2_0),
    .I_9_2_1(n105_I_9_2_1),
    .I_9_2_2(n105_I_9_2_2),
    .I_10_0_0(n105_I_10_0_0),
    .I_10_0_1(n105_I_10_0_1),
    .I_10_0_2(n105_I_10_0_2),
    .I_10_1_0(n105_I_10_1_0),
    .I_10_1_1(n105_I_10_1_1),
    .I_10_1_2(n105_I_10_1_2),
    .I_10_2_0(n105_I_10_2_0),
    .I_10_2_1(n105_I_10_2_1),
    .I_10_2_2(n105_I_10_2_2),
    .I_11_0_0(n105_I_11_0_0),
    .I_11_0_1(n105_I_11_0_1),
    .I_11_0_2(n105_I_11_0_2),
    .I_11_1_0(n105_I_11_1_0),
    .I_11_1_1(n105_I_11_1_1),
    .I_11_1_2(n105_I_11_1_2),
    .I_11_2_0(n105_I_11_2_0),
    .I_11_2_1(n105_I_11_2_1),
    .I_11_2_2(n105_I_11_2_2),
    .I_12_0_0(n105_I_12_0_0),
    .I_12_0_1(n105_I_12_0_1),
    .I_12_0_2(n105_I_12_0_2),
    .I_12_1_0(n105_I_12_1_0),
    .I_12_1_1(n105_I_12_1_1),
    .I_12_1_2(n105_I_12_1_2),
    .I_12_2_0(n105_I_12_2_0),
    .I_12_2_1(n105_I_12_2_1),
    .I_12_2_2(n105_I_12_2_2),
    .I_13_0_0(n105_I_13_0_0),
    .I_13_0_1(n105_I_13_0_1),
    .I_13_0_2(n105_I_13_0_2),
    .I_13_1_0(n105_I_13_1_0),
    .I_13_1_1(n105_I_13_1_1),
    .I_13_1_2(n105_I_13_1_2),
    .I_13_2_0(n105_I_13_2_0),
    .I_13_2_1(n105_I_13_2_1),
    .I_13_2_2(n105_I_13_2_2),
    .I_14_0_0(n105_I_14_0_0),
    .I_14_0_1(n105_I_14_0_1),
    .I_14_0_2(n105_I_14_0_2),
    .I_14_1_0(n105_I_14_1_0),
    .I_14_1_1(n105_I_14_1_1),
    .I_14_1_2(n105_I_14_1_2),
    .I_14_2_0(n105_I_14_2_0),
    .I_14_2_1(n105_I_14_2_1),
    .I_14_2_2(n105_I_14_2_2),
    .I_15_0_0(n105_I_15_0_0),
    .I_15_0_1(n105_I_15_0_1),
    .I_15_0_2(n105_I_15_0_2),
    .I_15_1_0(n105_I_15_1_0),
    .I_15_1_1(n105_I_15_1_1),
    .I_15_1_2(n105_I_15_1_2),
    .I_15_2_0(n105_I_15_2_0),
    .I_15_2_1(n105_I_15_2_1),
    .I_15_2_2(n105_I_15_2_2),
    .O_0_0_0(n105_O_0_0_0),
    .O_1_0_0(n105_O_1_0_0),
    .O_2_0_0(n105_O_2_0_0),
    .O_3_0_0(n105_O_3_0_0),
    .O_4_0_0(n105_O_4_0_0),
    .O_5_0_0(n105_O_5_0_0),
    .O_6_0_0(n105_O_6_0_0),
    .O_7_0_0(n105_O_7_0_0),
    .O_8_0_0(n105_O_8_0_0),
    .O_9_0_0(n105_O_9_0_0),
    .O_10_0_0(n105_O_10_0_0),
    .O_11_0_0(n105_O_11_0_0),
    .O_12_0_0(n105_O_12_0_0),
    .O_13_0_0(n105_O_13_0_0),
    .O_14_0_0(n105_O_14_0_0),
    .O_15_0_0(n105_O_15_0_0)
  );
  UnpartitionS n106 ( // @[Top.scala 202:22]
    .valid_up(n106_valid_up),
    .valid_down(n106_valid_down),
    .I_0_0_0(n106_I_0_0_0),
    .I_1_0_0(n106_I_1_0_0),
    .I_2_0_0(n106_I_2_0_0),
    .I_3_0_0(n106_I_3_0_0),
    .I_4_0_0(n106_I_4_0_0),
    .I_5_0_0(n106_I_5_0_0),
    .I_6_0_0(n106_I_6_0_0),
    .I_7_0_0(n106_I_7_0_0),
    .I_8_0_0(n106_I_8_0_0),
    .I_9_0_0(n106_I_9_0_0),
    .I_10_0_0(n106_I_10_0_0),
    .I_11_0_0(n106_I_11_0_0),
    .I_12_0_0(n106_I_12_0_0),
    .I_13_0_0(n106_I_13_0_0),
    .I_14_0_0(n106_I_14_0_0),
    .I_15_0_0(n106_I_15_0_0),
    .O_0_0(n106_O_0_0),
    .O_1_0(n106_O_1_0),
    .O_2_0(n106_O_2_0),
    .O_3_0(n106_O_3_0),
    .O_4_0(n106_O_4_0),
    .O_5_0(n106_O_5_0),
    .O_6_0(n106_O_6_0),
    .O_7_0(n106_O_7_0),
    .O_8_0(n106_O_8_0),
    .O_9_0(n106_O_9_0),
    .O_10_0(n106_O_10_0),
    .O_11_0(n106_O_11_0),
    .O_12_0(n106_O_12_0),
    .O_13_0(n106_O_13_0),
    .O_14_0(n106_O_14_0),
    .O_15_0(n106_O_15_0)
  );
  UnpartitionS_1 n107 ( // @[Top.scala 205:22]
    .valid_up(n107_valid_up),
    .valid_down(n107_valid_down),
    .I_0_0(n107_I_0_0),
    .I_1_0(n107_I_1_0),
    .I_2_0(n107_I_2_0),
    .I_3_0(n107_I_3_0),
    .I_4_0(n107_I_4_0),
    .I_5_0(n107_I_5_0),
    .I_6_0(n107_I_6_0),
    .I_7_0(n107_I_7_0),
    .I_8_0(n107_I_8_0),
    .I_9_0(n107_I_9_0),
    .I_10_0(n107_I_10_0),
    .I_11_0(n107_I_11_0),
    .I_12_0(n107_I_12_0),
    .I_13_0(n107_I_13_0),
    .I_14_0(n107_I_14_0),
    .I_15_0(n107_I_15_0),
    .O_0(n107_O_0),
    .O_1(n107_O_1),
    .O_2(n107_O_2),
    .O_3(n107_O_3),
    .O_4(n107_O_4),
    .O_5(n107_O_5),
    .O_6(n107_O_6),
    .O_7(n107_O_7),
    .O_8(n107_O_8),
    .O_9(n107_O_9),
    .O_10(n107_O_10),
    .O_11(n107_O_11),
    .O_12(n107_O_12),
    .O_13(n107_O_13),
    .O_14(n107_O_14),
    .O_15(n107_O_15)
  );
  FIFO_1 n108 ( // @[Top.scala 208:22]
    .clock(n108_clock),
    .reset(n108_reset),
    .valid_up(n108_valid_up),
    .valid_down(n108_valid_down),
    .I_0(n108_I_0),
    .I_1(n108_I_1),
    .I_2(n108_I_2),
    .I_3(n108_I_3),
    .I_4(n108_I_4),
    .I_5(n108_I_5),
    .I_6(n108_I_6),
    .I_7(n108_I_7),
    .I_8(n108_I_8),
    .I_9(n108_I_9),
    .I_10(n108_I_10),
    .I_11(n108_I_11),
    .I_12(n108_I_12),
    .I_13(n108_I_13),
    .I_14(n108_I_14),
    .I_15(n108_I_15),
    .O_0(n108_O_0),
    .O_1(n108_O_1),
    .O_2(n108_O_2),
    .O_3(n108_O_3),
    .O_4(n108_O_4),
    .O_5(n108_O_5),
    .O_6(n108_O_6),
    .O_7(n108_O_7),
    .O_8(n108_O_8),
    .O_9(n108_O_9),
    .O_10(n108_O_10),
    .O_11(n108_O_11),
    .O_12(n108_O_12),
    .O_13(n108_O_13),
    .O_14(n108_O_14),
    .O_15(n108_O_15)
  );
  Map2S_12 n109 ( // @[Top.scala 211:22]
    .clock(n109_clock),
    .reset(n109_reset),
    .valid_up(n109_valid_up),
    .valid_down(n109_valid_down),
    .I0_0(n109_I0_0),
    .I0_1(n109_I0_1),
    .I0_2(n109_I0_2),
    .I0_3(n109_I0_3),
    .I0_4(n109_I0_4),
    .I0_5(n109_I0_5),
    .I0_6(n109_I0_6),
    .I0_7(n109_I0_7),
    .I0_8(n109_I0_8),
    .I0_9(n109_I0_9),
    .I0_10(n109_I0_10),
    .I0_11(n109_I0_11),
    .I0_12(n109_I0_12),
    .I0_13(n109_I0_13),
    .I0_14(n109_I0_14),
    .I0_15(n109_I0_15),
    .I1_0(n109_I1_0),
    .I1_1(n109_I1_1),
    .I1_2(n109_I1_2),
    .I1_3(n109_I1_3),
    .I1_4(n109_I1_4),
    .I1_5(n109_I1_5),
    .I1_6(n109_I1_6),
    .I1_7(n109_I1_7),
    .I1_8(n109_I1_8),
    .I1_9(n109_I1_9),
    .I1_10(n109_I1_10),
    .I1_11(n109_I1_11),
    .I1_12(n109_I1_12),
    .I1_13(n109_I1_13),
    .I1_14(n109_I1_14),
    .I1_15(n109_I1_15),
    .O_0(n109_O_0),
    .O_1(n109_O_1),
    .O_2(n109_O_2),
    .O_3(n109_O_3),
    .O_4(n109_O_4),
    .O_5(n109_O_5),
    .O_6(n109_O_6),
    .O_7(n109_O_7),
    .O_8(n109_O_8),
    .O_9(n109_O_9),
    .O_10(n109_O_10),
    .O_11(n109_O_11),
    .O_12(n109_O_12),
    .O_13(n109_O_13),
    .O_14(n109_O_14),
    .O_15(n109_O_15)
  );
  FIFO n136 ( // @[Top.scala 215:22]
    .clock(n136_clock),
    .reset(n136_reset),
    .valid_up(n136_valid_up),
    .valid_down(n136_valid_down),
    .I_0(n136_I_0),
    .I_1(n136_I_1),
    .I_2(n136_I_2),
    .I_3(n136_I_3),
    .I_4(n136_I_4),
    .I_5(n136_I_5),
    .I_6(n136_I_6),
    .I_7(n136_I_7),
    .I_8(n136_I_8),
    .I_9(n136_I_9),
    .I_10(n136_I_10),
    .I_11(n136_I_11),
    .I_12(n136_I_12),
    .I_13(n136_I_13),
    .I_14(n136_I_14),
    .I_15(n136_I_15),
    .O_0(n136_O_0),
    .O_1(n136_O_1),
    .O_2(n136_O_2),
    .O_3(n136_O_3),
    .O_4(n136_O_4),
    .O_5(n136_O_5),
    .O_6(n136_O_6),
    .O_7(n136_O_7),
    .O_8(n136_O_8),
    .O_9(n136_O_9),
    .O_10(n136_O_10),
    .O_11(n136_O_11),
    .O_12(n136_O_12),
    .O_13(n136_O_13),
    .O_14(n136_O_14),
    .O_15(n136_O_15)
  );
  FIFO n137 ( // @[Top.scala 218:22]
    .clock(n137_clock),
    .reset(n137_reset),
    .valid_up(n137_valid_up),
    .valid_down(n137_valid_down),
    .I_0(n137_I_0),
    .I_1(n137_I_1),
    .I_2(n137_I_2),
    .I_3(n137_I_3),
    .I_4(n137_I_4),
    .I_5(n137_I_5),
    .I_6(n137_I_6),
    .I_7(n137_I_7),
    .I_8(n137_I_8),
    .I_9(n137_I_9),
    .I_10(n137_I_10),
    .I_11(n137_I_11),
    .I_12(n137_I_12),
    .I_13(n137_I_13),
    .I_14(n137_I_14),
    .I_15(n137_I_15),
    .O_0(n137_O_0),
    .O_1(n137_O_1),
    .O_2(n137_O_2),
    .O_3(n137_O_3),
    .O_4(n137_O_4),
    .O_5(n137_O_5),
    .O_6(n137_O_6),
    .O_7(n137_O_7),
    .O_8(n137_O_8),
    .O_9(n137_O_9),
    .O_10(n137_O_10),
    .O_11(n137_O_11),
    .O_12(n137_O_12),
    .O_13(n137_O_13),
    .O_14(n137_O_14),
    .O_15(n137_O_15)
  );
  FIFO n138 ( // @[Top.scala 221:22]
    .clock(n138_clock),
    .reset(n138_reset),
    .valid_up(n138_valid_up),
    .valid_down(n138_valid_down),
    .I_0(n138_I_0),
    .I_1(n138_I_1),
    .I_2(n138_I_2),
    .I_3(n138_I_3),
    .I_4(n138_I_4),
    .I_5(n138_I_5),
    .I_6(n138_I_6),
    .I_7(n138_I_7),
    .I_8(n138_I_8),
    .I_9(n138_I_9),
    .I_10(n138_I_10),
    .I_11(n138_I_11),
    .I_12(n138_I_12),
    .I_13(n138_I_13),
    .I_14(n138_I_14),
    .I_15(n138_I_15),
    .O_0(n138_O_0),
    .O_1(n138_O_1),
    .O_2(n138_O_2),
    .O_3(n138_O_3),
    .O_4(n138_O_4),
    .O_5(n138_O_5),
    .O_6(n138_O_6),
    .O_7(n138_O_7),
    .O_8(n138_O_8),
    .O_9(n138_O_9),
    .O_10(n138_O_10),
    .O_11(n138_O_11),
    .O_12(n138_O_12),
    .O_13(n138_O_13),
    .O_14(n138_O_14),
    .O_15(n138_O_15)
  );
  assign valid_down = n138_valid_down; // @[Top.scala 225:16]
  assign O_0 = n138_O_0; // @[Top.scala 224:7]
  assign O_1 = n138_O_1; // @[Top.scala 224:7]
  assign O_2 = n138_O_2; // @[Top.scala 224:7]
  assign O_3 = n138_O_3; // @[Top.scala 224:7]
  assign O_4 = n138_O_4; // @[Top.scala 224:7]
  assign O_5 = n138_O_5; // @[Top.scala 224:7]
  assign O_6 = n138_O_6; // @[Top.scala 224:7]
  assign O_7 = n138_O_7; // @[Top.scala 224:7]
  assign O_8 = n138_O_8; // @[Top.scala 224:7]
  assign O_9 = n138_O_9; // @[Top.scala 224:7]
  assign O_10 = n138_O_10; // @[Top.scala 224:7]
  assign O_11 = n138_O_11; // @[Top.scala 224:7]
  assign O_12 = n138_O_12; // @[Top.scala 224:7]
  assign O_13 = n138_O_13; // @[Top.scala 224:7]
  assign O_14 = n138_O_14; // @[Top.scala 224:7]
  assign O_15 = n138_O_15; // @[Top.scala 224:7]
  assign n1_clock = clock;
  assign n1_reset = reset;
  assign n1_valid_up = valid_up; // @[Top.scala 118:17]
  assign n1_I_0 = I_0; // @[Top.scala 117:10]
  assign n1_I_1 = I_1; // @[Top.scala 117:10]
  assign n1_I_2 = I_2; // @[Top.scala 117:10]
  assign n1_I_3 = I_3; // @[Top.scala 117:10]
  assign n1_I_4 = I_4; // @[Top.scala 117:10]
  assign n1_I_5 = I_5; // @[Top.scala 117:10]
  assign n1_I_6 = I_6; // @[Top.scala 117:10]
  assign n1_I_7 = I_7; // @[Top.scala 117:10]
  assign n1_I_8 = I_8; // @[Top.scala 117:10]
  assign n1_I_9 = I_9; // @[Top.scala 117:10]
  assign n1_I_10 = I_10; // @[Top.scala 117:10]
  assign n1_I_11 = I_11; // @[Top.scala 117:10]
  assign n1_I_12 = I_12; // @[Top.scala 117:10]
  assign n1_I_13 = I_13; // @[Top.scala 117:10]
  assign n1_I_14 = I_14; // @[Top.scala 117:10]
  assign n1_I_15 = I_15; // @[Top.scala 117:10]
  assign n2_valid_up = n1_valid_down; // @[Top.scala 121:17]
  assign n2_I_0 = n1_O_0; // @[Top.scala 120:10]
  assign n2_I_1 = n1_O_1; // @[Top.scala 120:10]
  assign n2_I_2 = n1_O_2; // @[Top.scala 120:10]
  assign n2_I_3 = n1_O_3; // @[Top.scala 120:10]
  assign n2_I_4 = n1_O_4; // @[Top.scala 120:10]
  assign n2_I_5 = n1_O_5; // @[Top.scala 120:10]
  assign n2_I_6 = n1_O_6; // @[Top.scala 120:10]
  assign n2_I_7 = n1_O_7; // @[Top.scala 120:10]
  assign n2_I_8 = n1_O_8; // @[Top.scala 120:10]
  assign n2_I_9 = n1_O_9; // @[Top.scala 120:10]
  assign n2_I_10 = n1_O_10; // @[Top.scala 120:10]
  assign n2_I_11 = n1_O_11; // @[Top.scala 120:10]
  assign n2_I_12 = n1_O_12; // @[Top.scala 120:10]
  assign n2_I_13 = n1_O_13; // @[Top.scala 120:10]
  assign n2_I_14 = n1_O_14; // @[Top.scala 120:10]
  assign n2_I_15 = n1_O_15; // @[Top.scala 120:10]
  assign n3_valid_up = n2_valid_down; // @[Top.scala 124:17]
  assign n3_I_0 = n2_O_0; // @[Top.scala 123:10]
  assign n3_I_1 = n2_O_1; // @[Top.scala 123:10]
  assign n3_I_2 = n2_O_2; // @[Top.scala 123:10]
  assign n3_I_3 = n2_O_3; // @[Top.scala 123:10]
  assign n3_I_4 = n2_O_4; // @[Top.scala 123:10]
  assign n3_I_5 = n2_O_5; // @[Top.scala 123:10]
  assign n3_I_6 = n2_O_6; // @[Top.scala 123:10]
  assign n3_I_7 = n2_O_7; // @[Top.scala 123:10]
  assign n3_I_8 = n2_O_8; // @[Top.scala 123:10]
  assign n3_I_9 = n2_O_9; // @[Top.scala 123:10]
  assign n3_I_10 = n2_O_10; // @[Top.scala 123:10]
  assign n3_I_11 = n2_O_11; // @[Top.scala 123:10]
  assign n3_I_12 = n2_O_12; // @[Top.scala 123:10]
  assign n3_I_13 = n2_O_13; // @[Top.scala 123:10]
  assign n3_I_14 = n2_O_14; // @[Top.scala 123:10]
  assign n3_I_15 = n2_O_15; // @[Top.scala 123:10]
  assign n4_valid_up = n3_valid_down; // @[Top.scala 127:17]
  assign n4_I_0 = n3_O_0; // @[Top.scala 126:10]
  assign n4_I_1 = n3_O_1; // @[Top.scala 126:10]
  assign n4_I_2 = n3_O_2; // @[Top.scala 126:10]
  assign n4_I_3 = n3_O_3; // @[Top.scala 126:10]
  assign n4_I_4 = n3_O_4; // @[Top.scala 126:10]
  assign n4_I_5 = n3_O_5; // @[Top.scala 126:10]
  assign n4_I_6 = n3_O_6; // @[Top.scala 126:10]
  assign n4_I_7 = n3_O_7; // @[Top.scala 126:10]
  assign n4_I_8 = n3_O_8; // @[Top.scala 126:10]
  assign n4_I_9 = n3_O_9; // @[Top.scala 126:10]
  assign n4_I_10 = n3_O_10; // @[Top.scala 126:10]
  assign n4_I_11 = n3_O_11; // @[Top.scala 126:10]
  assign n4_I_12 = n3_O_12; // @[Top.scala 126:10]
  assign n4_I_13 = n3_O_13; // @[Top.scala 126:10]
  assign n4_I_14 = n3_O_14; // @[Top.scala 126:10]
  assign n4_I_15 = n3_O_15; // @[Top.scala 126:10]
  assign n5_valid_up = n4_valid_down; // @[Top.scala 130:17]
  assign n5_I_0 = n4_O_0; // @[Top.scala 129:10]
  assign n5_I_1 = n4_O_1; // @[Top.scala 129:10]
  assign n5_I_2 = n4_O_2; // @[Top.scala 129:10]
  assign n5_I_3 = n4_O_3; // @[Top.scala 129:10]
  assign n5_I_4 = n4_O_4; // @[Top.scala 129:10]
  assign n5_I_5 = n4_O_5; // @[Top.scala 129:10]
  assign n5_I_6 = n4_O_6; // @[Top.scala 129:10]
  assign n5_I_7 = n4_O_7; // @[Top.scala 129:10]
  assign n5_I_8 = n4_O_8; // @[Top.scala 129:10]
  assign n5_I_9 = n4_O_9; // @[Top.scala 129:10]
  assign n5_I_10 = n4_O_10; // @[Top.scala 129:10]
  assign n5_I_11 = n4_O_11; // @[Top.scala 129:10]
  assign n5_I_12 = n4_O_12; // @[Top.scala 129:10]
  assign n5_I_13 = n4_O_13; // @[Top.scala 129:10]
  assign n5_I_14 = n4_O_14; // @[Top.scala 129:10]
  assign n5_I_15 = n4_O_15; // @[Top.scala 129:10]
  assign n6_valid_up = n5_valid_down & n4_valid_down; // @[Top.scala 134:17]
  assign n6_I0_0 = n5_O_0; // @[Top.scala 132:11]
  assign n6_I0_1 = n5_O_1; // @[Top.scala 132:11]
  assign n6_I0_2 = n5_O_2; // @[Top.scala 132:11]
  assign n6_I0_3 = n5_O_3; // @[Top.scala 132:11]
  assign n6_I0_4 = n5_O_4; // @[Top.scala 132:11]
  assign n6_I0_5 = n5_O_5; // @[Top.scala 132:11]
  assign n6_I0_6 = n5_O_6; // @[Top.scala 132:11]
  assign n6_I0_7 = n5_O_7; // @[Top.scala 132:11]
  assign n6_I0_8 = n5_O_8; // @[Top.scala 132:11]
  assign n6_I0_9 = n5_O_9; // @[Top.scala 132:11]
  assign n6_I0_10 = n5_O_10; // @[Top.scala 132:11]
  assign n6_I0_11 = n5_O_11; // @[Top.scala 132:11]
  assign n6_I0_12 = n5_O_12; // @[Top.scala 132:11]
  assign n6_I0_13 = n5_O_13; // @[Top.scala 132:11]
  assign n6_I0_14 = n5_O_14; // @[Top.scala 132:11]
  assign n6_I0_15 = n5_O_15; // @[Top.scala 132:11]
  assign n6_I1_0 = n4_O_0; // @[Top.scala 133:11]
  assign n6_I1_1 = n4_O_1; // @[Top.scala 133:11]
  assign n6_I1_2 = n4_O_2; // @[Top.scala 133:11]
  assign n6_I1_3 = n4_O_3; // @[Top.scala 133:11]
  assign n6_I1_4 = n4_O_4; // @[Top.scala 133:11]
  assign n6_I1_5 = n4_O_5; // @[Top.scala 133:11]
  assign n6_I1_6 = n4_O_6; // @[Top.scala 133:11]
  assign n6_I1_7 = n4_O_7; // @[Top.scala 133:11]
  assign n6_I1_8 = n4_O_8; // @[Top.scala 133:11]
  assign n6_I1_9 = n4_O_9; // @[Top.scala 133:11]
  assign n6_I1_10 = n4_O_10; // @[Top.scala 133:11]
  assign n6_I1_11 = n4_O_11; // @[Top.scala 133:11]
  assign n6_I1_12 = n4_O_12; // @[Top.scala 133:11]
  assign n6_I1_13 = n4_O_13; // @[Top.scala 133:11]
  assign n6_I1_14 = n4_O_14; // @[Top.scala 133:11]
  assign n6_I1_15 = n4_O_15; // @[Top.scala 133:11]
  assign n10_valid_up = n6_valid_down & n3_valid_down; // @[Top.scala 138:18]
  assign n10_I0_0_0 = n6_O_0_0; // @[Top.scala 136:12]
  assign n10_I0_0_1 = n6_O_0_1; // @[Top.scala 136:12]
  assign n10_I0_1_0 = n6_O_1_0; // @[Top.scala 136:12]
  assign n10_I0_1_1 = n6_O_1_1; // @[Top.scala 136:12]
  assign n10_I0_2_0 = n6_O_2_0; // @[Top.scala 136:12]
  assign n10_I0_2_1 = n6_O_2_1; // @[Top.scala 136:12]
  assign n10_I0_3_0 = n6_O_3_0; // @[Top.scala 136:12]
  assign n10_I0_3_1 = n6_O_3_1; // @[Top.scala 136:12]
  assign n10_I0_4_0 = n6_O_4_0; // @[Top.scala 136:12]
  assign n10_I0_4_1 = n6_O_4_1; // @[Top.scala 136:12]
  assign n10_I0_5_0 = n6_O_5_0; // @[Top.scala 136:12]
  assign n10_I0_5_1 = n6_O_5_1; // @[Top.scala 136:12]
  assign n10_I0_6_0 = n6_O_6_0; // @[Top.scala 136:12]
  assign n10_I0_6_1 = n6_O_6_1; // @[Top.scala 136:12]
  assign n10_I0_7_0 = n6_O_7_0; // @[Top.scala 136:12]
  assign n10_I0_7_1 = n6_O_7_1; // @[Top.scala 136:12]
  assign n10_I0_8_0 = n6_O_8_0; // @[Top.scala 136:12]
  assign n10_I0_8_1 = n6_O_8_1; // @[Top.scala 136:12]
  assign n10_I0_9_0 = n6_O_9_0; // @[Top.scala 136:12]
  assign n10_I0_9_1 = n6_O_9_1; // @[Top.scala 136:12]
  assign n10_I0_10_0 = n6_O_10_0; // @[Top.scala 136:12]
  assign n10_I0_10_1 = n6_O_10_1; // @[Top.scala 136:12]
  assign n10_I0_11_0 = n6_O_11_0; // @[Top.scala 136:12]
  assign n10_I0_11_1 = n6_O_11_1; // @[Top.scala 136:12]
  assign n10_I0_12_0 = n6_O_12_0; // @[Top.scala 136:12]
  assign n10_I0_12_1 = n6_O_12_1; // @[Top.scala 136:12]
  assign n10_I0_13_0 = n6_O_13_0; // @[Top.scala 136:12]
  assign n10_I0_13_1 = n6_O_13_1; // @[Top.scala 136:12]
  assign n10_I0_14_0 = n6_O_14_0; // @[Top.scala 136:12]
  assign n10_I0_14_1 = n6_O_14_1; // @[Top.scala 136:12]
  assign n10_I0_15_0 = n6_O_15_0; // @[Top.scala 136:12]
  assign n10_I0_15_1 = n6_O_15_1; // @[Top.scala 136:12]
  assign n10_I1_0 = n3_O_0; // @[Top.scala 137:12]
  assign n10_I1_1 = n3_O_1; // @[Top.scala 137:12]
  assign n10_I1_2 = n3_O_2; // @[Top.scala 137:12]
  assign n10_I1_3 = n3_O_3; // @[Top.scala 137:12]
  assign n10_I1_4 = n3_O_4; // @[Top.scala 137:12]
  assign n10_I1_5 = n3_O_5; // @[Top.scala 137:12]
  assign n10_I1_6 = n3_O_6; // @[Top.scala 137:12]
  assign n10_I1_7 = n3_O_7; // @[Top.scala 137:12]
  assign n10_I1_8 = n3_O_8; // @[Top.scala 137:12]
  assign n10_I1_9 = n3_O_9; // @[Top.scala 137:12]
  assign n10_I1_10 = n3_O_10; // @[Top.scala 137:12]
  assign n10_I1_11 = n3_O_11; // @[Top.scala 137:12]
  assign n10_I1_12 = n3_O_12; // @[Top.scala 137:12]
  assign n10_I1_13 = n3_O_13; // @[Top.scala 137:12]
  assign n10_I1_14 = n3_O_14; // @[Top.scala 137:12]
  assign n10_I1_15 = n3_O_15; // @[Top.scala 137:12]
  assign n14_valid_up = n10_valid_down; // @[Top.scala 141:18]
  assign n14_I_0_0 = n10_O_0_0; // @[Top.scala 140:11]
  assign n14_I_0_1 = n10_O_0_1; // @[Top.scala 140:11]
  assign n14_I_0_2 = n10_O_0_2; // @[Top.scala 140:11]
  assign n14_I_1_0 = n10_O_1_0; // @[Top.scala 140:11]
  assign n14_I_1_1 = n10_O_1_1; // @[Top.scala 140:11]
  assign n14_I_1_2 = n10_O_1_2; // @[Top.scala 140:11]
  assign n14_I_2_0 = n10_O_2_0; // @[Top.scala 140:11]
  assign n14_I_2_1 = n10_O_2_1; // @[Top.scala 140:11]
  assign n14_I_2_2 = n10_O_2_2; // @[Top.scala 140:11]
  assign n14_I_3_0 = n10_O_3_0; // @[Top.scala 140:11]
  assign n14_I_3_1 = n10_O_3_1; // @[Top.scala 140:11]
  assign n14_I_3_2 = n10_O_3_2; // @[Top.scala 140:11]
  assign n14_I_4_0 = n10_O_4_0; // @[Top.scala 140:11]
  assign n14_I_4_1 = n10_O_4_1; // @[Top.scala 140:11]
  assign n14_I_4_2 = n10_O_4_2; // @[Top.scala 140:11]
  assign n14_I_5_0 = n10_O_5_0; // @[Top.scala 140:11]
  assign n14_I_5_1 = n10_O_5_1; // @[Top.scala 140:11]
  assign n14_I_5_2 = n10_O_5_2; // @[Top.scala 140:11]
  assign n14_I_6_0 = n10_O_6_0; // @[Top.scala 140:11]
  assign n14_I_6_1 = n10_O_6_1; // @[Top.scala 140:11]
  assign n14_I_6_2 = n10_O_6_2; // @[Top.scala 140:11]
  assign n14_I_7_0 = n10_O_7_0; // @[Top.scala 140:11]
  assign n14_I_7_1 = n10_O_7_1; // @[Top.scala 140:11]
  assign n14_I_7_2 = n10_O_7_2; // @[Top.scala 140:11]
  assign n14_I_8_0 = n10_O_8_0; // @[Top.scala 140:11]
  assign n14_I_8_1 = n10_O_8_1; // @[Top.scala 140:11]
  assign n14_I_8_2 = n10_O_8_2; // @[Top.scala 140:11]
  assign n14_I_9_0 = n10_O_9_0; // @[Top.scala 140:11]
  assign n14_I_9_1 = n10_O_9_1; // @[Top.scala 140:11]
  assign n14_I_9_2 = n10_O_9_2; // @[Top.scala 140:11]
  assign n14_I_10_0 = n10_O_10_0; // @[Top.scala 140:11]
  assign n14_I_10_1 = n10_O_10_1; // @[Top.scala 140:11]
  assign n14_I_10_2 = n10_O_10_2; // @[Top.scala 140:11]
  assign n14_I_11_0 = n10_O_11_0; // @[Top.scala 140:11]
  assign n14_I_11_1 = n10_O_11_1; // @[Top.scala 140:11]
  assign n14_I_11_2 = n10_O_11_2; // @[Top.scala 140:11]
  assign n14_I_12_0 = n10_O_12_0; // @[Top.scala 140:11]
  assign n14_I_12_1 = n10_O_12_1; // @[Top.scala 140:11]
  assign n14_I_12_2 = n10_O_12_2; // @[Top.scala 140:11]
  assign n14_I_13_0 = n10_O_13_0; // @[Top.scala 140:11]
  assign n14_I_13_1 = n10_O_13_1; // @[Top.scala 140:11]
  assign n14_I_13_2 = n10_O_13_2; // @[Top.scala 140:11]
  assign n14_I_14_0 = n10_O_14_0; // @[Top.scala 140:11]
  assign n14_I_14_1 = n10_O_14_1; // @[Top.scala 140:11]
  assign n14_I_14_2 = n10_O_14_2; // @[Top.scala 140:11]
  assign n14_I_15_0 = n10_O_15_0; // @[Top.scala 140:11]
  assign n14_I_15_1 = n10_O_15_1; // @[Top.scala 140:11]
  assign n14_I_15_2 = n10_O_15_2; // @[Top.scala 140:11]
  assign n19_valid_up = n14_valid_down; // @[Top.scala 144:18]
  assign n19_I_0_0_0 = n14_O_0_0_0; // @[Top.scala 143:11]
  assign n19_I_0_0_1 = n14_O_0_0_1; // @[Top.scala 143:11]
  assign n19_I_0_0_2 = n14_O_0_0_2; // @[Top.scala 143:11]
  assign n19_I_1_0_0 = n14_O_1_0_0; // @[Top.scala 143:11]
  assign n19_I_1_0_1 = n14_O_1_0_1; // @[Top.scala 143:11]
  assign n19_I_1_0_2 = n14_O_1_0_2; // @[Top.scala 143:11]
  assign n19_I_2_0_0 = n14_O_2_0_0; // @[Top.scala 143:11]
  assign n19_I_2_0_1 = n14_O_2_0_1; // @[Top.scala 143:11]
  assign n19_I_2_0_2 = n14_O_2_0_2; // @[Top.scala 143:11]
  assign n19_I_3_0_0 = n14_O_3_0_0; // @[Top.scala 143:11]
  assign n19_I_3_0_1 = n14_O_3_0_1; // @[Top.scala 143:11]
  assign n19_I_3_0_2 = n14_O_3_0_2; // @[Top.scala 143:11]
  assign n19_I_4_0_0 = n14_O_4_0_0; // @[Top.scala 143:11]
  assign n19_I_4_0_1 = n14_O_4_0_1; // @[Top.scala 143:11]
  assign n19_I_4_0_2 = n14_O_4_0_2; // @[Top.scala 143:11]
  assign n19_I_5_0_0 = n14_O_5_0_0; // @[Top.scala 143:11]
  assign n19_I_5_0_1 = n14_O_5_0_1; // @[Top.scala 143:11]
  assign n19_I_5_0_2 = n14_O_5_0_2; // @[Top.scala 143:11]
  assign n19_I_6_0_0 = n14_O_6_0_0; // @[Top.scala 143:11]
  assign n19_I_6_0_1 = n14_O_6_0_1; // @[Top.scala 143:11]
  assign n19_I_6_0_2 = n14_O_6_0_2; // @[Top.scala 143:11]
  assign n19_I_7_0_0 = n14_O_7_0_0; // @[Top.scala 143:11]
  assign n19_I_7_0_1 = n14_O_7_0_1; // @[Top.scala 143:11]
  assign n19_I_7_0_2 = n14_O_7_0_2; // @[Top.scala 143:11]
  assign n19_I_8_0_0 = n14_O_8_0_0; // @[Top.scala 143:11]
  assign n19_I_8_0_1 = n14_O_8_0_1; // @[Top.scala 143:11]
  assign n19_I_8_0_2 = n14_O_8_0_2; // @[Top.scala 143:11]
  assign n19_I_9_0_0 = n14_O_9_0_0; // @[Top.scala 143:11]
  assign n19_I_9_0_1 = n14_O_9_0_1; // @[Top.scala 143:11]
  assign n19_I_9_0_2 = n14_O_9_0_2; // @[Top.scala 143:11]
  assign n19_I_10_0_0 = n14_O_10_0_0; // @[Top.scala 143:11]
  assign n19_I_10_0_1 = n14_O_10_0_1; // @[Top.scala 143:11]
  assign n19_I_10_0_2 = n14_O_10_0_2; // @[Top.scala 143:11]
  assign n19_I_11_0_0 = n14_O_11_0_0; // @[Top.scala 143:11]
  assign n19_I_11_0_1 = n14_O_11_0_1; // @[Top.scala 143:11]
  assign n19_I_11_0_2 = n14_O_11_0_2; // @[Top.scala 143:11]
  assign n19_I_12_0_0 = n14_O_12_0_0; // @[Top.scala 143:11]
  assign n19_I_12_0_1 = n14_O_12_0_1; // @[Top.scala 143:11]
  assign n19_I_12_0_2 = n14_O_12_0_2; // @[Top.scala 143:11]
  assign n19_I_13_0_0 = n14_O_13_0_0; // @[Top.scala 143:11]
  assign n19_I_13_0_1 = n14_O_13_0_1; // @[Top.scala 143:11]
  assign n19_I_13_0_2 = n14_O_13_0_2; // @[Top.scala 143:11]
  assign n19_I_14_0_0 = n14_O_14_0_0; // @[Top.scala 143:11]
  assign n19_I_14_0_1 = n14_O_14_0_1; // @[Top.scala 143:11]
  assign n19_I_14_0_2 = n14_O_14_0_2; // @[Top.scala 143:11]
  assign n19_I_15_0_0 = n14_O_15_0_0; // @[Top.scala 143:11]
  assign n19_I_15_0_1 = n14_O_15_0_1; // @[Top.scala 143:11]
  assign n19_I_15_0_2 = n14_O_15_0_2; // @[Top.scala 143:11]
  assign n20_valid_up = n2_valid_down; // @[Top.scala 147:18]
  assign n20_I_0 = n2_O_0; // @[Top.scala 146:11]
  assign n20_I_1 = n2_O_1; // @[Top.scala 146:11]
  assign n20_I_2 = n2_O_2; // @[Top.scala 146:11]
  assign n20_I_3 = n2_O_3; // @[Top.scala 146:11]
  assign n20_I_4 = n2_O_4; // @[Top.scala 146:11]
  assign n20_I_5 = n2_O_5; // @[Top.scala 146:11]
  assign n20_I_6 = n2_O_6; // @[Top.scala 146:11]
  assign n20_I_7 = n2_O_7; // @[Top.scala 146:11]
  assign n20_I_8 = n2_O_8; // @[Top.scala 146:11]
  assign n20_I_9 = n2_O_9; // @[Top.scala 146:11]
  assign n20_I_10 = n2_O_10; // @[Top.scala 146:11]
  assign n20_I_11 = n2_O_11; // @[Top.scala 146:11]
  assign n20_I_12 = n2_O_12; // @[Top.scala 146:11]
  assign n20_I_13 = n2_O_13; // @[Top.scala 146:11]
  assign n20_I_14 = n2_O_14; // @[Top.scala 146:11]
  assign n20_I_15 = n2_O_15; // @[Top.scala 146:11]
  assign n21_valid_up = n20_valid_down; // @[Top.scala 150:18]
  assign n21_I_0 = n20_O_0; // @[Top.scala 149:11]
  assign n21_I_1 = n20_O_1; // @[Top.scala 149:11]
  assign n21_I_2 = n20_O_2; // @[Top.scala 149:11]
  assign n21_I_3 = n20_O_3; // @[Top.scala 149:11]
  assign n21_I_4 = n20_O_4; // @[Top.scala 149:11]
  assign n21_I_5 = n20_O_5; // @[Top.scala 149:11]
  assign n21_I_6 = n20_O_6; // @[Top.scala 149:11]
  assign n21_I_7 = n20_O_7; // @[Top.scala 149:11]
  assign n21_I_8 = n20_O_8; // @[Top.scala 149:11]
  assign n21_I_9 = n20_O_9; // @[Top.scala 149:11]
  assign n21_I_10 = n20_O_10; // @[Top.scala 149:11]
  assign n21_I_11 = n20_O_11; // @[Top.scala 149:11]
  assign n21_I_12 = n20_O_12; // @[Top.scala 149:11]
  assign n21_I_13 = n20_O_13; // @[Top.scala 149:11]
  assign n21_I_14 = n20_O_14; // @[Top.scala 149:11]
  assign n21_I_15 = n20_O_15; // @[Top.scala 149:11]
  assign n22_valid_up = n21_valid_down & n20_valid_down; // @[Top.scala 154:18]
  assign n22_I0_0 = n21_O_0; // @[Top.scala 152:12]
  assign n22_I0_1 = n21_O_1; // @[Top.scala 152:12]
  assign n22_I0_2 = n21_O_2; // @[Top.scala 152:12]
  assign n22_I0_3 = n21_O_3; // @[Top.scala 152:12]
  assign n22_I0_4 = n21_O_4; // @[Top.scala 152:12]
  assign n22_I0_5 = n21_O_5; // @[Top.scala 152:12]
  assign n22_I0_6 = n21_O_6; // @[Top.scala 152:12]
  assign n22_I0_7 = n21_O_7; // @[Top.scala 152:12]
  assign n22_I0_8 = n21_O_8; // @[Top.scala 152:12]
  assign n22_I0_9 = n21_O_9; // @[Top.scala 152:12]
  assign n22_I0_10 = n21_O_10; // @[Top.scala 152:12]
  assign n22_I0_11 = n21_O_11; // @[Top.scala 152:12]
  assign n22_I0_12 = n21_O_12; // @[Top.scala 152:12]
  assign n22_I0_13 = n21_O_13; // @[Top.scala 152:12]
  assign n22_I0_14 = n21_O_14; // @[Top.scala 152:12]
  assign n22_I0_15 = n21_O_15; // @[Top.scala 152:12]
  assign n22_I1_0 = n20_O_0; // @[Top.scala 153:12]
  assign n22_I1_1 = n20_O_1; // @[Top.scala 153:12]
  assign n22_I1_2 = n20_O_2; // @[Top.scala 153:12]
  assign n22_I1_3 = n20_O_3; // @[Top.scala 153:12]
  assign n22_I1_4 = n20_O_4; // @[Top.scala 153:12]
  assign n22_I1_5 = n20_O_5; // @[Top.scala 153:12]
  assign n22_I1_6 = n20_O_6; // @[Top.scala 153:12]
  assign n22_I1_7 = n20_O_7; // @[Top.scala 153:12]
  assign n22_I1_8 = n20_O_8; // @[Top.scala 153:12]
  assign n22_I1_9 = n20_O_9; // @[Top.scala 153:12]
  assign n22_I1_10 = n20_O_10; // @[Top.scala 153:12]
  assign n22_I1_11 = n20_O_11; // @[Top.scala 153:12]
  assign n22_I1_12 = n20_O_12; // @[Top.scala 153:12]
  assign n22_I1_13 = n20_O_13; // @[Top.scala 153:12]
  assign n22_I1_14 = n20_O_14; // @[Top.scala 153:12]
  assign n22_I1_15 = n20_O_15; // @[Top.scala 153:12]
  assign n26_valid_up = n22_valid_down & n2_valid_down; // @[Top.scala 158:18]
  assign n26_I0_0_0 = n22_O_0_0; // @[Top.scala 156:12]
  assign n26_I0_0_1 = n22_O_0_1; // @[Top.scala 156:12]
  assign n26_I0_1_0 = n22_O_1_0; // @[Top.scala 156:12]
  assign n26_I0_1_1 = n22_O_1_1; // @[Top.scala 156:12]
  assign n26_I0_2_0 = n22_O_2_0; // @[Top.scala 156:12]
  assign n26_I0_2_1 = n22_O_2_1; // @[Top.scala 156:12]
  assign n26_I0_3_0 = n22_O_3_0; // @[Top.scala 156:12]
  assign n26_I0_3_1 = n22_O_3_1; // @[Top.scala 156:12]
  assign n26_I0_4_0 = n22_O_4_0; // @[Top.scala 156:12]
  assign n26_I0_4_1 = n22_O_4_1; // @[Top.scala 156:12]
  assign n26_I0_5_0 = n22_O_5_0; // @[Top.scala 156:12]
  assign n26_I0_5_1 = n22_O_5_1; // @[Top.scala 156:12]
  assign n26_I0_6_0 = n22_O_6_0; // @[Top.scala 156:12]
  assign n26_I0_6_1 = n22_O_6_1; // @[Top.scala 156:12]
  assign n26_I0_7_0 = n22_O_7_0; // @[Top.scala 156:12]
  assign n26_I0_7_1 = n22_O_7_1; // @[Top.scala 156:12]
  assign n26_I0_8_0 = n22_O_8_0; // @[Top.scala 156:12]
  assign n26_I0_8_1 = n22_O_8_1; // @[Top.scala 156:12]
  assign n26_I0_9_0 = n22_O_9_0; // @[Top.scala 156:12]
  assign n26_I0_9_1 = n22_O_9_1; // @[Top.scala 156:12]
  assign n26_I0_10_0 = n22_O_10_0; // @[Top.scala 156:12]
  assign n26_I0_10_1 = n22_O_10_1; // @[Top.scala 156:12]
  assign n26_I0_11_0 = n22_O_11_0; // @[Top.scala 156:12]
  assign n26_I0_11_1 = n22_O_11_1; // @[Top.scala 156:12]
  assign n26_I0_12_0 = n22_O_12_0; // @[Top.scala 156:12]
  assign n26_I0_12_1 = n22_O_12_1; // @[Top.scala 156:12]
  assign n26_I0_13_0 = n22_O_13_0; // @[Top.scala 156:12]
  assign n26_I0_13_1 = n22_O_13_1; // @[Top.scala 156:12]
  assign n26_I0_14_0 = n22_O_14_0; // @[Top.scala 156:12]
  assign n26_I0_14_1 = n22_O_14_1; // @[Top.scala 156:12]
  assign n26_I0_15_0 = n22_O_15_0; // @[Top.scala 156:12]
  assign n26_I0_15_1 = n22_O_15_1; // @[Top.scala 156:12]
  assign n26_I1_0 = n2_O_0; // @[Top.scala 157:12]
  assign n26_I1_1 = n2_O_1; // @[Top.scala 157:12]
  assign n26_I1_2 = n2_O_2; // @[Top.scala 157:12]
  assign n26_I1_3 = n2_O_3; // @[Top.scala 157:12]
  assign n26_I1_4 = n2_O_4; // @[Top.scala 157:12]
  assign n26_I1_5 = n2_O_5; // @[Top.scala 157:12]
  assign n26_I1_6 = n2_O_6; // @[Top.scala 157:12]
  assign n26_I1_7 = n2_O_7; // @[Top.scala 157:12]
  assign n26_I1_8 = n2_O_8; // @[Top.scala 157:12]
  assign n26_I1_9 = n2_O_9; // @[Top.scala 157:12]
  assign n26_I1_10 = n2_O_10; // @[Top.scala 157:12]
  assign n26_I1_11 = n2_O_11; // @[Top.scala 157:12]
  assign n26_I1_12 = n2_O_12; // @[Top.scala 157:12]
  assign n26_I1_13 = n2_O_13; // @[Top.scala 157:12]
  assign n26_I1_14 = n2_O_14; // @[Top.scala 157:12]
  assign n26_I1_15 = n2_O_15; // @[Top.scala 157:12]
  assign n30_valid_up = n26_valid_down; // @[Top.scala 161:18]
  assign n30_I_0_0 = n26_O_0_0; // @[Top.scala 160:11]
  assign n30_I_0_1 = n26_O_0_1; // @[Top.scala 160:11]
  assign n30_I_0_2 = n26_O_0_2; // @[Top.scala 160:11]
  assign n30_I_1_0 = n26_O_1_0; // @[Top.scala 160:11]
  assign n30_I_1_1 = n26_O_1_1; // @[Top.scala 160:11]
  assign n30_I_1_2 = n26_O_1_2; // @[Top.scala 160:11]
  assign n30_I_2_0 = n26_O_2_0; // @[Top.scala 160:11]
  assign n30_I_2_1 = n26_O_2_1; // @[Top.scala 160:11]
  assign n30_I_2_2 = n26_O_2_2; // @[Top.scala 160:11]
  assign n30_I_3_0 = n26_O_3_0; // @[Top.scala 160:11]
  assign n30_I_3_1 = n26_O_3_1; // @[Top.scala 160:11]
  assign n30_I_3_2 = n26_O_3_2; // @[Top.scala 160:11]
  assign n30_I_4_0 = n26_O_4_0; // @[Top.scala 160:11]
  assign n30_I_4_1 = n26_O_4_1; // @[Top.scala 160:11]
  assign n30_I_4_2 = n26_O_4_2; // @[Top.scala 160:11]
  assign n30_I_5_0 = n26_O_5_0; // @[Top.scala 160:11]
  assign n30_I_5_1 = n26_O_5_1; // @[Top.scala 160:11]
  assign n30_I_5_2 = n26_O_5_2; // @[Top.scala 160:11]
  assign n30_I_6_0 = n26_O_6_0; // @[Top.scala 160:11]
  assign n30_I_6_1 = n26_O_6_1; // @[Top.scala 160:11]
  assign n30_I_6_2 = n26_O_6_2; // @[Top.scala 160:11]
  assign n30_I_7_0 = n26_O_7_0; // @[Top.scala 160:11]
  assign n30_I_7_1 = n26_O_7_1; // @[Top.scala 160:11]
  assign n30_I_7_2 = n26_O_7_2; // @[Top.scala 160:11]
  assign n30_I_8_0 = n26_O_8_0; // @[Top.scala 160:11]
  assign n30_I_8_1 = n26_O_8_1; // @[Top.scala 160:11]
  assign n30_I_8_2 = n26_O_8_2; // @[Top.scala 160:11]
  assign n30_I_9_0 = n26_O_9_0; // @[Top.scala 160:11]
  assign n30_I_9_1 = n26_O_9_1; // @[Top.scala 160:11]
  assign n30_I_9_2 = n26_O_9_2; // @[Top.scala 160:11]
  assign n30_I_10_0 = n26_O_10_0; // @[Top.scala 160:11]
  assign n30_I_10_1 = n26_O_10_1; // @[Top.scala 160:11]
  assign n30_I_10_2 = n26_O_10_2; // @[Top.scala 160:11]
  assign n30_I_11_0 = n26_O_11_0; // @[Top.scala 160:11]
  assign n30_I_11_1 = n26_O_11_1; // @[Top.scala 160:11]
  assign n30_I_11_2 = n26_O_11_2; // @[Top.scala 160:11]
  assign n30_I_12_0 = n26_O_12_0; // @[Top.scala 160:11]
  assign n30_I_12_1 = n26_O_12_1; // @[Top.scala 160:11]
  assign n30_I_12_2 = n26_O_12_2; // @[Top.scala 160:11]
  assign n30_I_13_0 = n26_O_13_0; // @[Top.scala 160:11]
  assign n30_I_13_1 = n26_O_13_1; // @[Top.scala 160:11]
  assign n30_I_13_2 = n26_O_13_2; // @[Top.scala 160:11]
  assign n30_I_14_0 = n26_O_14_0; // @[Top.scala 160:11]
  assign n30_I_14_1 = n26_O_14_1; // @[Top.scala 160:11]
  assign n30_I_14_2 = n26_O_14_2; // @[Top.scala 160:11]
  assign n30_I_15_0 = n26_O_15_0; // @[Top.scala 160:11]
  assign n30_I_15_1 = n26_O_15_1; // @[Top.scala 160:11]
  assign n30_I_15_2 = n26_O_15_2; // @[Top.scala 160:11]
  assign n35_valid_up = n30_valid_down; // @[Top.scala 164:18]
  assign n35_I_0_0_0 = n30_O_0_0_0; // @[Top.scala 163:11]
  assign n35_I_0_0_1 = n30_O_0_0_1; // @[Top.scala 163:11]
  assign n35_I_0_0_2 = n30_O_0_0_2; // @[Top.scala 163:11]
  assign n35_I_1_0_0 = n30_O_1_0_0; // @[Top.scala 163:11]
  assign n35_I_1_0_1 = n30_O_1_0_1; // @[Top.scala 163:11]
  assign n35_I_1_0_2 = n30_O_1_0_2; // @[Top.scala 163:11]
  assign n35_I_2_0_0 = n30_O_2_0_0; // @[Top.scala 163:11]
  assign n35_I_2_0_1 = n30_O_2_0_1; // @[Top.scala 163:11]
  assign n35_I_2_0_2 = n30_O_2_0_2; // @[Top.scala 163:11]
  assign n35_I_3_0_0 = n30_O_3_0_0; // @[Top.scala 163:11]
  assign n35_I_3_0_1 = n30_O_3_0_1; // @[Top.scala 163:11]
  assign n35_I_3_0_2 = n30_O_3_0_2; // @[Top.scala 163:11]
  assign n35_I_4_0_0 = n30_O_4_0_0; // @[Top.scala 163:11]
  assign n35_I_4_0_1 = n30_O_4_0_1; // @[Top.scala 163:11]
  assign n35_I_4_0_2 = n30_O_4_0_2; // @[Top.scala 163:11]
  assign n35_I_5_0_0 = n30_O_5_0_0; // @[Top.scala 163:11]
  assign n35_I_5_0_1 = n30_O_5_0_1; // @[Top.scala 163:11]
  assign n35_I_5_0_2 = n30_O_5_0_2; // @[Top.scala 163:11]
  assign n35_I_6_0_0 = n30_O_6_0_0; // @[Top.scala 163:11]
  assign n35_I_6_0_1 = n30_O_6_0_1; // @[Top.scala 163:11]
  assign n35_I_6_0_2 = n30_O_6_0_2; // @[Top.scala 163:11]
  assign n35_I_7_0_0 = n30_O_7_0_0; // @[Top.scala 163:11]
  assign n35_I_7_0_1 = n30_O_7_0_1; // @[Top.scala 163:11]
  assign n35_I_7_0_2 = n30_O_7_0_2; // @[Top.scala 163:11]
  assign n35_I_8_0_0 = n30_O_8_0_0; // @[Top.scala 163:11]
  assign n35_I_8_0_1 = n30_O_8_0_1; // @[Top.scala 163:11]
  assign n35_I_8_0_2 = n30_O_8_0_2; // @[Top.scala 163:11]
  assign n35_I_9_0_0 = n30_O_9_0_0; // @[Top.scala 163:11]
  assign n35_I_9_0_1 = n30_O_9_0_1; // @[Top.scala 163:11]
  assign n35_I_9_0_2 = n30_O_9_0_2; // @[Top.scala 163:11]
  assign n35_I_10_0_0 = n30_O_10_0_0; // @[Top.scala 163:11]
  assign n35_I_10_0_1 = n30_O_10_0_1; // @[Top.scala 163:11]
  assign n35_I_10_0_2 = n30_O_10_0_2; // @[Top.scala 163:11]
  assign n35_I_11_0_0 = n30_O_11_0_0; // @[Top.scala 163:11]
  assign n35_I_11_0_1 = n30_O_11_0_1; // @[Top.scala 163:11]
  assign n35_I_11_0_2 = n30_O_11_0_2; // @[Top.scala 163:11]
  assign n35_I_12_0_0 = n30_O_12_0_0; // @[Top.scala 163:11]
  assign n35_I_12_0_1 = n30_O_12_0_1; // @[Top.scala 163:11]
  assign n35_I_12_0_2 = n30_O_12_0_2; // @[Top.scala 163:11]
  assign n35_I_13_0_0 = n30_O_13_0_0; // @[Top.scala 163:11]
  assign n35_I_13_0_1 = n30_O_13_0_1; // @[Top.scala 163:11]
  assign n35_I_13_0_2 = n30_O_13_0_2; // @[Top.scala 163:11]
  assign n35_I_14_0_0 = n30_O_14_0_0; // @[Top.scala 163:11]
  assign n35_I_14_0_1 = n30_O_14_0_1; // @[Top.scala 163:11]
  assign n35_I_14_0_2 = n30_O_14_0_2; // @[Top.scala 163:11]
  assign n35_I_15_0_0 = n30_O_15_0_0; // @[Top.scala 163:11]
  assign n35_I_15_0_1 = n30_O_15_0_1; // @[Top.scala 163:11]
  assign n35_I_15_0_2 = n30_O_15_0_2; // @[Top.scala 163:11]
  assign n36_valid_up = n19_valid_down & n35_valid_down; // @[Top.scala 168:18]
  assign n36_I0_0_0 = n19_O_0_0; // @[Top.scala 166:12]
  assign n36_I0_0_1 = n19_O_0_1; // @[Top.scala 166:12]
  assign n36_I0_0_2 = n19_O_0_2; // @[Top.scala 166:12]
  assign n36_I0_1_0 = n19_O_1_0; // @[Top.scala 166:12]
  assign n36_I0_1_1 = n19_O_1_1; // @[Top.scala 166:12]
  assign n36_I0_1_2 = n19_O_1_2; // @[Top.scala 166:12]
  assign n36_I0_2_0 = n19_O_2_0; // @[Top.scala 166:12]
  assign n36_I0_2_1 = n19_O_2_1; // @[Top.scala 166:12]
  assign n36_I0_2_2 = n19_O_2_2; // @[Top.scala 166:12]
  assign n36_I0_3_0 = n19_O_3_0; // @[Top.scala 166:12]
  assign n36_I0_3_1 = n19_O_3_1; // @[Top.scala 166:12]
  assign n36_I0_3_2 = n19_O_3_2; // @[Top.scala 166:12]
  assign n36_I0_4_0 = n19_O_4_0; // @[Top.scala 166:12]
  assign n36_I0_4_1 = n19_O_4_1; // @[Top.scala 166:12]
  assign n36_I0_4_2 = n19_O_4_2; // @[Top.scala 166:12]
  assign n36_I0_5_0 = n19_O_5_0; // @[Top.scala 166:12]
  assign n36_I0_5_1 = n19_O_5_1; // @[Top.scala 166:12]
  assign n36_I0_5_2 = n19_O_5_2; // @[Top.scala 166:12]
  assign n36_I0_6_0 = n19_O_6_0; // @[Top.scala 166:12]
  assign n36_I0_6_1 = n19_O_6_1; // @[Top.scala 166:12]
  assign n36_I0_6_2 = n19_O_6_2; // @[Top.scala 166:12]
  assign n36_I0_7_0 = n19_O_7_0; // @[Top.scala 166:12]
  assign n36_I0_7_1 = n19_O_7_1; // @[Top.scala 166:12]
  assign n36_I0_7_2 = n19_O_7_2; // @[Top.scala 166:12]
  assign n36_I0_8_0 = n19_O_8_0; // @[Top.scala 166:12]
  assign n36_I0_8_1 = n19_O_8_1; // @[Top.scala 166:12]
  assign n36_I0_8_2 = n19_O_8_2; // @[Top.scala 166:12]
  assign n36_I0_9_0 = n19_O_9_0; // @[Top.scala 166:12]
  assign n36_I0_9_1 = n19_O_9_1; // @[Top.scala 166:12]
  assign n36_I0_9_2 = n19_O_9_2; // @[Top.scala 166:12]
  assign n36_I0_10_0 = n19_O_10_0; // @[Top.scala 166:12]
  assign n36_I0_10_1 = n19_O_10_1; // @[Top.scala 166:12]
  assign n36_I0_10_2 = n19_O_10_2; // @[Top.scala 166:12]
  assign n36_I0_11_0 = n19_O_11_0; // @[Top.scala 166:12]
  assign n36_I0_11_1 = n19_O_11_1; // @[Top.scala 166:12]
  assign n36_I0_11_2 = n19_O_11_2; // @[Top.scala 166:12]
  assign n36_I0_12_0 = n19_O_12_0; // @[Top.scala 166:12]
  assign n36_I0_12_1 = n19_O_12_1; // @[Top.scala 166:12]
  assign n36_I0_12_2 = n19_O_12_2; // @[Top.scala 166:12]
  assign n36_I0_13_0 = n19_O_13_0; // @[Top.scala 166:12]
  assign n36_I0_13_1 = n19_O_13_1; // @[Top.scala 166:12]
  assign n36_I0_13_2 = n19_O_13_2; // @[Top.scala 166:12]
  assign n36_I0_14_0 = n19_O_14_0; // @[Top.scala 166:12]
  assign n36_I0_14_1 = n19_O_14_1; // @[Top.scala 166:12]
  assign n36_I0_14_2 = n19_O_14_2; // @[Top.scala 166:12]
  assign n36_I0_15_0 = n19_O_15_0; // @[Top.scala 166:12]
  assign n36_I0_15_1 = n19_O_15_1; // @[Top.scala 166:12]
  assign n36_I0_15_2 = n19_O_15_2; // @[Top.scala 166:12]
  assign n36_I1_0_0 = n35_O_0_0; // @[Top.scala 167:12]
  assign n36_I1_0_1 = n35_O_0_1; // @[Top.scala 167:12]
  assign n36_I1_0_2 = n35_O_0_2; // @[Top.scala 167:12]
  assign n36_I1_1_0 = n35_O_1_0; // @[Top.scala 167:12]
  assign n36_I1_1_1 = n35_O_1_1; // @[Top.scala 167:12]
  assign n36_I1_1_2 = n35_O_1_2; // @[Top.scala 167:12]
  assign n36_I1_2_0 = n35_O_2_0; // @[Top.scala 167:12]
  assign n36_I1_2_1 = n35_O_2_1; // @[Top.scala 167:12]
  assign n36_I1_2_2 = n35_O_2_2; // @[Top.scala 167:12]
  assign n36_I1_3_0 = n35_O_3_0; // @[Top.scala 167:12]
  assign n36_I1_3_1 = n35_O_3_1; // @[Top.scala 167:12]
  assign n36_I1_3_2 = n35_O_3_2; // @[Top.scala 167:12]
  assign n36_I1_4_0 = n35_O_4_0; // @[Top.scala 167:12]
  assign n36_I1_4_1 = n35_O_4_1; // @[Top.scala 167:12]
  assign n36_I1_4_2 = n35_O_4_2; // @[Top.scala 167:12]
  assign n36_I1_5_0 = n35_O_5_0; // @[Top.scala 167:12]
  assign n36_I1_5_1 = n35_O_5_1; // @[Top.scala 167:12]
  assign n36_I1_5_2 = n35_O_5_2; // @[Top.scala 167:12]
  assign n36_I1_6_0 = n35_O_6_0; // @[Top.scala 167:12]
  assign n36_I1_6_1 = n35_O_6_1; // @[Top.scala 167:12]
  assign n36_I1_6_2 = n35_O_6_2; // @[Top.scala 167:12]
  assign n36_I1_7_0 = n35_O_7_0; // @[Top.scala 167:12]
  assign n36_I1_7_1 = n35_O_7_1; // @[Top.scala 167:12]
  assign n36_I1_7_2 = n35_O_7_2; // @[Top.scala 167:12]
  assign n36_I1_8_0 = n35_O_8_0; // @[Top.scala 167:12]
  assign n36_I1_8_1 = n35_O_8_1; // @[Top.scala 167:12]
  assign n36_I1_8_2 = n35_O_8_2; // @[Top.scala 167:12]
  assign n36_I1_9_0 = n35_O_9_0; // @[Top.scala 167:12]
  assign n36_I1_9_1 = n35_O_9_1; // @[Top.scala 167:12]
  assign n36_I1_9_2 = n35_O_9_2; // @[Top.scala 167:12]
  assign n36_I1_10_0 = n35_O_10_0; // @[Top.scala 167:12]
  assign n36_I1_10_1 = n35_O_10_1; // @[Top.scala 167:12]
  assign n36_I1_10_2 = n35_O_10_2; // @[Top.scala 167:12]
  assign n36_I1_11_0 = n35_O_11_0; // @[Top.scala 167:12]
  assign n36_I1_11_1 = n35_O_11_1; // @[Top.scala 167:12]
  assign n36_I1_11_2 = n35_O_11_2; // @[Top.scala 167:12]
  assign n36_I1_12_0 = n35_O_12_0; // @[Top.scala 167:12]
  assign n36_I1_12_1 = n35_O_12_1; // @[Top.scala 167:12]
  assign n36_I1_12_2 = n35_O_12_2; // @[Top.scala 167:12]
  assign n36_I1_13_0 = n35_O_13_0; // @[Top.scala 167:12]
  assign n36_I1_13_1 = n35_O_13_1; // @[Top.scala 167:12]
  assign n36_I1_13_2 = n35_O_13_2; // @[Top.scala 167:12]
  assign n36_I1_14_0 = n35_O_14_0; // @[Top.scala 167:12]
  assign n36_I1_14_1 = n35_O_14_1; // @[Top.scala 167:12]
  assign n36_I1_14_2 = n35_O_14_2; // @[Top.scala 167:12]
  assign n36_I1_15_0 = n35_O_15_0; // @[Top.scala 167:12]
  assign n36_I1_15_1 = n35_O_15_1; // @[Top.scala 167:12]
  assign n36_I1_15_2 = n35_O_15_2; // @[Top.scala 167:12]
  assign n40_valid_up = n1_valid_down; // @[Top.scala 171:18]
  assign n40_I_0 = n1_O_0; // @[Top.scala 170:11]
  assign n40_I_1 = n1_O_1; // @[Top.scala 170:11]
  assign n40_I_2 = n1_O_2; // @[Top.scala 170:11]
  assign n40_I_3 = n1_O_3; // @[Top.scala 170:11]
  assign n40_I_4 = n1_O_4; // @[Top.scala 170:11]
  assign n40_I_5 = n1_O_5; // @[Top.scala 170:11]
  assign n40_I_6 = n1_O_6; // @[Top.scala 170:11]
  assign n40_I_7 = n1_O_7; // @[Top.scala 170:11]
  assign n40_I_8 = n1_O_8; // @[Top.scala 170:11]
  assign n40_I_9 = n1_O_9; // @[Top.scala 170:11]
  assign n40_I_10 = n1_O_10; // @[Top.scala 170:11]
  assign n40_I_11 = n1_O_11; // @[Top.scala 170:11]
  assign n40_I_12 = n1_O_12; // @[Top.scala 170:11]
  assign n40_I_13 = n1_O_13; // @[Top.scala 170:11]
  assign n40_I_14 = n1_O_14; // @[Top.scala 170:11]
  assign n40_I_15 = n1_O_15; // @[Top.scala 170:11]
  assign n41_valid_up = n40_valid_down; // @[Top.scala 174:18]
  assign n41_I_0 = n40_O_0; // @[Top.scala 173:11]
  assign n41_I_1 = n40_O_1; // @[Top.scala 173:11]
  assign n41_I_2 = n40_O_2; // @[Top.scala 173:11]
  assign n41_I_3 = n40_O_3; // @[Top.scala 173:11]
  assign n41_I_4 = n40_O_4; // @[Top.scala 173:11]
  assign n41_I_5 = n40_O_5; // @[Top.scala 173:11]
  assign n41_I_6 = n40_O_6; // @[Top.scala 173:11]
  assign n41_I_7 = n40_O_7; // @[Top.scala 173:11]
  assign n41_I_8 = n40_O_8; // @[Top.scala 173:11]
  assign n41_I_9 = n40_O_9; // @[Top.scala 173:11]
  assign n41_I_10 = n40_O_10; // @[Top.scala 173:11]
  assign n41_I_11 = n40_O_11; // @[Top.scala 173:11]
  assign n41_I_12 = n40_O_12; // @[Top.scala 173:11]
  assign n41_I_13 = n40_O_13; // @[Top.scala 173:11]
  assign n41_I_14 = n40_O_14; // @[Top.scala 173:11]
  assign n41_I_15 = n40_O_15; // @[Top.scala 173:11]
  assign n42_valid_up = n41_valid_down & n40_valid_down; // @[Top.scala 178:18]
  assign n42_I0_0 = n41_O_0; // @[Top.scala 176:12]
  assign n42_I0_1 = n41_O_1; // @[Top.scala 176:12]
  assign n42_I0_2 = n41_O_2; // @[Top.scala 176:12]
  assign n42_I0_3 = n41_O_3; // @[Top.scala 176:12]
  assign n42_I0_4 = n41_O_4; // @[Top.scala 176:12]
  assign n42_I0_5 = n41_O_5; // @[Top.scala 176:12]
  assign n42_I0_6 = n41_O_6; // @[Top.scala 176:12]
  assign n42_I0_7 = n41_O_7; // @[Top.scala 176:12]
  assign n42_I0_8 = n41_O_8; // @[Top.scala 176:12]
  assign n42_I0_9 = n41_O_9; // @[Top.scala 176:12]
  assign n42_I0_10 = n41_O_10; // @[Top.scala 176:12]
  assign n42_I0_11 = n41_O_11; // @[Top.scala 176:12]
  assign n42_I0_12 = n41_O_12; // @[Top.scala 176:12]
  assign n42_I0_13 = n41_O_13; // @[Top.scala 176:12]
  assign n42_I0_14 = n41_O_14; // @[Top.scala 176:12]
  assign n42_I0_15 = n41_O_15; // @[Top.scala 176:12]
  assign n42_I1_0 = n40_O_0; // @[Top.scala 177:12]
  assign n42_I1_1 = n40_O_1; // @[Top.scala 177:12]
  assign n42_I1_2 = n40_O_2; // @[Top.scala 177:12]
  assign n42_I1_3 = n40_O_3; // @[Top.scala 177:12]
  assign n42_I1_4 = n40_O_4; // @[Top.scala 177:12]
  assign n42_I1_5 = n40_O_5; // @[Top.scala 177:12]
  assign n42_I1_6 = n40_O_6; // @[Top.scala 177:12]
  assign n42_I1_7 = n40_O_7; // @[Top.scala 177:12]
  assign n42_I1_8 = n40_O_8; // @[Top.scala 177:12]
  assign n42_I1_9 = n40_O_9; // @[Top.scala 177:12]
  assign n42_I1_10 = n40_O_10; // @[Top.scala 177:12]
  assign n42_I1_11 = n40_O_11; // @[Top.scala 177:12]
  assign n42_I1_12 = n40_O_12; // @[Top.scala 177:12]
  assign n42_I1_13 = n40_O_13; // @[Top.scala 177:12]
  assign n42_I1_14 = n40_O_14; // @[Top.scala 177:12]
  assign n42_I1_15 = n40_O_15; // @[Top.scala 177:12]
  assign n46_valid_up = n42_valid_down & n1_valid_down; // @[Top.scala 182:18]
  assign n46_I0_0_0 = n42_O_0_0; // @[Top.scala 180:12]
  assign n46_I0_0_1 = n42_O_0_1; // @[Top.scala 180:12]
  assign n46_I0_1_0 = n42_O_1_0; // @[Top.scala 180:12]
  assign n46_I0_1_1 = n42_O_1_1; // @[Top.scala 180:12]
  assign n46_I0_2_0 = n42_O_2_0; // @[Top.scala 180:12]
  assign n46_I0_2_1 = n42_O_2_1; // @[Top.scala 180:12]
  assign n46_I0_3_0 = n42_O_3_0; // @[Top.scala 180:12]
  assign n46_I0_3_1 = n42_O_3_1; // @[Top.scala 180:12]
  assign n46_I0_4_0 = n42_O_4_0; // @[Top.scala 180:12]
  assign n46_I0_4_1 = n42_O_4_1; // @[Top.scala 180:12]
  assign n46_I0_5_0 = n42_O_5_0; // @[Top.scala 180:12]
  assign n46_I0_5_1 = n42_O_5_1; // @[Top.scala 180:12]
  assign n46_I0_6_0 = n42_O_6_0; // @[Top.scala 180:12]
  assign n46_I0_6_1 = n42_O_6_1; // @[Top.scala 180:12]
  assign n46_I0_7_0 = n42_O_7_0; // @[Top.scala 180:12]
  assign n46_I0_7_1 = n42_O_7_1; // @[Top.scala 180:12]
  assign n46_I0_8_0 = n42_O_8_0; // @[Top.scala 180:12]
  assign n46_I0_8_1 = n42_O_8_1; // @[Top.scala 180:12]
  assign n46_I0_9_0 = n42_O_9_0; // @[Top.scala 180:12]
  assign n46_I0_9_1 = n42_O_9_1; // @[Top.scala 180:12]
  assign n46_I0_10_0 = n42_O_10_0; // @[Top.scala 180:12]
  assign n46_I0_10_1 = n42_O_10_1; // @[Top.scala 180:12]
  assign n46_I0_11_0 = n42_O_11_0; // @[Top.scala 180:12]
  assign n46_I0_11_1 = n42_O_11_1; // @[Top.scala 180:12]
  assign n46_I0_12_0 = n42_O_12_0; // @[Top.scala 180:12]
  assign n46_I0_12_1 = n42_O_12_1; // @[Top.scala 180:12]
  assign n46_I0_13_0 = n42_O_13_0; // @[Top.scala 180:12]
  assign n46_I0_13_1 = n42_O_13_1; // @[Top.scala 180:12]
  assign n46_I0_14_0 = n42_O_14_0; // @[Top.scala 180:12]
  assign n46_I0_14_1 = n42_O_14_1; // @[Top.scala 180:12]
  assign n46_I0_15_0 = n42_O_15_0; // @[Top.scala 180:12]
  assign n46_I0_15_1 = n42_O_15_1; // @[Top.scala 180:12]
  assign n46_I1_0 = n1_O_0; // @[Top.scala 181:12]
  assign n46_I1_1 = n1_O_1; // @[Top.scala 181:12]
  assign n46_I1_2 = n1_O_2; // @[Top.scala 181:12]
  assign n46_I1_3 = n1_O_3; // @[Top.scala 181:12]
  assign n46_I1_4 = n1_O_4; // @[Top.scala 181:12]
  assign n46_I1_5 = n1_O_5; // @[Top.scala 181:12]
  assign n46_I1_6 = n1_O_6; // @[Top.scala 181:12]
  assign n46_I1_7 = n1_O_7; // @[Top.scala 181:12]
  assign n46_I1_8 = n1_O_8; // @[Top.scala 181:12]
  assign n46_I1_9 = n1_O_9; // @[Top.scala 181:12]
  assign n46_I1_10 = n1_O_10; // @[Top.scala 181:12]
  assign n46_I1_11 = n1_O_11; // @[Top.scala 181:12]
  assign n46_I1_12 = n1_O_12; // @[Top.scala 181:12]
  assign n46_I1_13 = n1_O_13; // @[Top.scala 181:12]
  assign n46_I1_14 = n1_O_14; // @[Top.scala 181:12]
  assign n46_I1_15 = n1_O_15; // @[Top.scala 181:12]
  assign n50_valid_up = n46_valid_down; // @[Top.scala 185:18]
  assign n50_I_0_0 = n46_O_0_0; // @[Top.scala 184:11]
  assign n50_I_0_1 = n46_O_0_1; // @[Top.scala 184:11]
  assign n50_I_0_2 = n46_O_0_2; // @[Top.scala 184:11]
  assign n50_I_1_0 = n46_O_1_0; // @[Top.scala 184:11]
  assign n50_I_1_1 = n46_O_1_1; // @[Top.scala 184:11]
  assign n50_I_1_2 = n46_O_1_2; // @[Top.scala 184:11]
  assign n50_I_2_0 = n46_O_2_0; // @[Top.scala 184:11]
  assign n50_I_2_1 = n46_O_2_1; // @[Top.scala 184:11]
  assign n50_I_2_2 = n46_O_2_2; // @[Top.scala 184:11]
  assign n50_I_3_0 = n46_O_3_0; // @[Top.scala 184:11]
  assign n50_I_3_1 = n46_O_3_1; // @[Top.scala 184:11]
  assign n50_I_3_2 = n46_O_3_2; // @[Top.scala 184:11]
  assign n50_I_4_0 = n46_O_4_0; // @[Top.scala 184:11]
  assign n50_I_4_1 = n46_O_4_1; // @[Top.scala 184:11]
  assign n50_I_4_2 = n46_O_4_2; // @[Top.scala 184:11]
  assign n50_I_5_0 = n46_O_5_0; // @[Top.scala 184:11]
  assign n50_I_5_1 = n46_O_5_1; // @[Top.scala 184:11]
  assign n50_I_5_2 = n46_O_5_2; // @[Top.scala 184:11]
  assign n50_I_6_0 = n46_O_6_0; // @[Top.scala 184:11]
  assign n50_I_6_1 = n46_O_6_1; // @[Top.scala 184:11]
  assign n50_I_6_2 = n46_O_6_2; // @[Top.scala 184:11]
  assign n50_I_7_0 = n46_O_7_0; // @[Top.scala 184:11]
  assign n50_I_7_1 = n46_O_7_1; // @[Top.scala 184:11]
  assign n50_I_7_2 = n46_O_7_2; // @[Top.scala 184:11]
  assign n50_I_8_0 = n46_O_8_0; // @[Top.scala 184:11]
  assign n50_I_8_1 = n46_O_8_1; // @[Top.scala 184:11]
  assign n50_I_8_2 = n46_O_8_2; // @[Top.scala 184:11]
  assign n50_I_9_0 = n46_O_9_0; // @[Top.scala 184:11]
  assign n50_I_9_1 = n46_O_9_1; // @[Top.scala 184:11]
  assign n50_I_9_2 = n46_O_9_2; // @[Top.scala 184:11]
  assign n50_I_10_0 = n46_O_10_0; // @[Top.scala 184:11]
  assign n50_I_10_1 = n46_O_10_1; // @[Top.scala 184:11]
  assign n50_I_10_2 = n46_O_10_2; // @[Top.scala 184:11]
  assign n50_I_11_0 = n46_O_11_0; // @[Top.scala 184:11]
  assign n50_I_11_1 = n46_O_11_1; // @[Top.scala 184:11]
  assign n50_I_11_2 = n46_O_11_2; // @[Top.scala 184:11]
  assign n50_I_12_0 = n46_O_12_0; // @[Top.scala 184:11]
  assign n50_I_12_1 = n46_O_12_1; // @[Top.scala 184:11]
  assign n50_I_12_2 = n46_O_12_2; // @[Top.scala 184:11]
  assign n50_I_13_0 = n46_O_13_0; // @[Top.scala 184:11]
  assign n50_I_13_1 = n46_O_13_1; // @[Top.scala 184:11]
  assign n50_I_13_2 = n46_O_13_2; // @[Top.scala 184:11]
  assign n50_I_14_0 = n46_O_14_0; // @[Top.scala 184:11]
  assign n50_I_14_1 = n46_O_14_1; // @[Top.scala 184:11]
  assign n50_I_14_2 = n46_O_14_2; // @[Top.scala 184:11]
  assign n50_I_15_0 = n46_O_15_0; // @[Top.scala 184:11]
  assign n50_I_15_1 = n46_O_15_1; // @[Top.scala 184:11]
  assign n50_I_15_2 = n46_O_15_2; // @[Top.scala 184:11]
  assign n55_valid_up = n50_valid_down; // @[Top.scala 188:18]
  assign n55_I_0_0_0 = n50_O_0_0_0; // @[Top.scala 187:11]
  assign n55_I_0_0_1 = n50_O_0_0_1; // @[Top.scala 187:11]
  assign n55_I_0_0_2 = n50_O_0_0_2; // @[Top.scala 187:11]
  assign n55_I_1_0_0 = n50_O_1_0_0; // @[Top.scala 187:11]
  assign n55_I_1_0_1 = n50_O_1_0_1; // @[Top.scala 187:11]
  assign n55_I_1_0_2 = n50_O_1_0_2; // @[Top.scala 187:11]
  assign n55_I_2_0_0 = n50_O_2_0_0; // @[Top.scala 187:11]
  assign n55_I_2_0_1 = n50_O_2_0_1; // @[Top.scala 187:11]
  assign n55_I_2_0_2 = n50_O_2_0_2; // @[Top.scala 187:11]
  assign n55_I_3_0_0 = n50_O_3_0_0; // @[Top.scala 187:11]
  assign n55_I_3_0_1 = n50_O_3_0_1; // @[Top.scala 187:11]
  assign n55_I_3_0_2 = n50_O_3_0_2; // @[Top.scala 187:11]
  assign n55_I_4_0_0 = n50_O_4_0_0; // @[Top.scala 187:11]
  assign n55_I_4_0_1 = n50_O_4_0_1; // @[Top.scala 187:11]
  assign n55_I_4_0_2 = n50_O_4_0_2; // @[Top.scala 187:11]
  assign n55_I_5_0_0 = n50_O_5_0_0; // @[Top.scala 187:11]
  assign n55_I_5_0_1 = n50_O_5_0_1; // @[Top.scala 187:11]
  assign n55_I_5_0_2 = n50_O_5_0_2; // @[Top.scala 187:11]
  assign n55_I_6_0_0 = n50_O_6_0_0; // @[Top.scala 187:11]
  assign n55_I_6_0_1 = n50_O_6_0_1; // @[Top.scala 187:11]
  assign n55_I_6_0_2 = n50_O_6_0_2; // @[Top.scala 187:11]
  assign n55_I_7_0_0 = n50_O_7_0_0; // @[Top.scala 187:11]
  assign n55_I_7_0_1 = n50_O_7_0_1; // @[Top.scala 187:11]
  assign n55_I_7_0_2 = n50_O_7_0_2; // @[Top.scala 187:11]
  assign n55_I_8_0_0 = n50_O_8_0_0; // @[Top.scala 187:11]
  assign n55_I_8_0_1 = n50_O_8_0_1; // @[Top.scala 187:11]
  assign n55_I_8_0_2 = n50_O_8_0_2; // @[Top.scala 187:11]
  assign n55_I_9_0_0 = n50_O_9_0_0; // @[Top.scala 187:11]
  assign n55_I_9_0_1 = n50_O_9_0_1; // @[Top.scala 187:11]
  assign n55_I_9_0_2 = n50_O_9_0_2; // @[Top.scala 187:11]
  assign n55_I_10_0_0 = n50_O_10_0_0; // @[Top.scala 187:11]
  assign n55_I_10_0_1 = n50_O_10_0_1; // @[Top.scala 187:11]
  assign n55_I_10_0_2 = n50_O_10_0_2; // @[Top.scala 187:11]
  assign n55_I_11_0_0 = n50_O_11_0_0; // @[Top.scala 187:11]
  assign n55_I_11_0_1 = n50_O_11_0_1; // @[Top.scala 187:11]
  assign n55_I_11_0_2 = n50_O_11_0_2; // @[Top.scala 187:11]
  assign n55_I_12_0_0 = n50_O_12_0_0; // @[Top.scala 187:11]
  assign n55_I_12_0_1 = n50_O_12_0_1; // @[Top.scala 187:11]
  assign n55_I_12_0_2 = n50_O_12_0_2; // @[Top.scala 187:11]
  assign n55_I_13_0_0 = n50_O_13_0_0; // @[Top.scala 187:11]
  assign n55_I_13_0_1 = n50_O_13_0_1; // @[Top.scala 187:11]
  assign n55_I_13_0_2 = n50_O_13_0_2; // @[Top.scala 187:11]
  assign n55_I_14_0_0 = n50_O_14_0_0; // @[Top.scala 187:11]
  assign n55_I_14_0_1 = n50_O_14_0_1; // @[Top.scala 187:11]
  assign n55_I_14_0_2 = n50_O_14_0_2; // @[Top.scala 187:11]
  assign n55_I_15_0_0 = n50_O_15_0_0; // @[Top.scala 187:11]
  assign n55_I_15_0_1 = n50_O_15_0_1; // @[Top.scala 187:11]
  assign n55_I_15_0_2 = n50_O_15_0_2; // @[Top.scala 187:11]
  assign n56_valid_up = n36_valid_down & n55_valid_down; // @[Top.scala 192:18]
  assign n56_I0_0_0_0 = n36_O_0_0_0; // @[Top.scala 190:12]
  assign n56_I0_0_0_1 = n36_O_0_0_1; // @[Top.scala 190:12]
  assign n56_I0_0_0_2 = n36_O_0_0_2; // @[Top.scala 190:12]
  assign n56_I0_0_1_0 = n36_O_0_1_0; // @[Top.scala 190:12]
  assign n56_I0_0_1_1 = n36_O_0_1_1; // @[Top.scala 190:12]
  assign n56_I0_0_1_2 = n36_O_0_1_2; // @[Top.scala 190:12]
  assign n56_I0_1_0_0 = n36_O_1_0_0; // @[Top.scala 190:12]
  assign n56_I0_1_0_1 = n36_O_1_0_1; // @[Top.scala 190:12]
  assign n56_I0_1_0_2 = n36_O_1_0_2; // @[Top.scala 190:12]
  assign n56_I0_1_1_0 = n36_O_1_1_0; // @[Top.scala 190:12]
  assign n56_I0_1_1_1 = n36_O_1_1_1; // @[Top.scala 190:12]
  assign n56_I0_1_1_2 = n36_O_1_1_2; // @[Top.scala 190:12]
  assign n56_I0_2_0_0 = n36_O_2_0_0; // @[Top.scala 190:12]
  assign n56_I0_2_0_1 = n36_O_2_0_1; // @[Top.scala 190:12]
  assign n56_I0_2_0_2 = n36_O_2_0_2; // @[Top.scala 190:12]
  assign n56_I0_2_1_0 = n36_O_2_1_0; // @[Top.scala 190:12]
  assign n56_I0_2_1_1 = n36_O_2_1_1; // @[Top.scala 190:12]
  assign n56_I0_2_1_2 = n36_O_2_1_2; // @[Top.scala 190:12]
  assign n56_I0_3_0_0 = n36_O_3_0_0; // @[Top.scala 190:12]
  assign n56_I0_3_0_1 = n36_O_3_0_1; // @[Top.scala 190:12]
  assign n56_I0_3_0_2 = n36_O_3_0_2; // @[Top.scala 190:12]
  assign n56_I0_3_1_0 = n36_O_3_1_0; // @[Top.scala 190:12]
  assign n56_I0_3_1_1 = n36_O_3_1_1; // @[Top.scala 190:12]
  assign n56_I0_3_1_2 = n36_O_3_1_2; // @[Top.scala 190:12]
  assign n56_I0_4_0_0 = n36_O_4_0_0; // @[Top.scala 190:12]
  assign n56_I0_4_0_1 = n36_O_4_0_1; // @[Top.scala 190:12]
  assign n56_I0_4_0_2 = n36_O_4_0_2; // @[Top.scala 190:12]
  assign n56_I0_4_1_0 = n36_O_4_1_0; // @[Top.scala 190:12]
  assign n56_I0_4_1_1 = n36_O_4_1_1; // @[Top.scala 190:12]
  assign n56_I0_4_1_2 = n36_O_4_1_2; // @[Top.scala 190:12]
  assign n56_I0_5_0_0 = n36_O_5_0_0; // @[Top.scala 190:12]
  assign n56_I0_5_0_1 = n36_O_5_0_1; // @[Top.scala 190:12]
  assign n56_I0_5_0_2 = n36_O_5_0_2; // @[Top.scala 190:12]
  assign n56_I0_5_1_0 = n36_O_5_1_0; // @[Top.scala 190:12]
  assign n56_I0_5_1_1 = n36_O_5_1_1; // @[Top.scala 190:12]
  assign n56_I0_5_1_2 = n36_O_5_1_2; // @[Top.scala 190:12]
  assign n56_I0_6_0_0 = n36_O_6_0_0; // @[Top.scala 190:12]
  assign n56_I0_6_0_1 = n36_O_6_0_1; // @[Top.scala 190:12]
  assign n56_I0_6_0_2 = n36_O_6_0_2; // @[Top.scala 190:12]
  assign n56_I0_6_1_0 = n36_O_6_1_0; // @[Top.scala 190:12]
  assign n56_I0_6_1_1 = n36_O_6_1_1; // @[Top.scala 190:12]
  assign n56_I0_6_1_2 = n36_O_6_1_2; // @[Top.scala 190:12]
  assign n56_I0_7_0_0 = n36_O_7_0_0; // @[Top.scala 190:12]
  assign n56_I0_7_0_1 = n36_O_7_0_1; // @[Top.scala 190:12]
  assign n56_I0_7_0_2 = n36_O_7_0_2; // @[Top.scala 190:12]
  assign n56_I0_7_1_0 = n36_O_7_1_0; // @[Top.scala 190:12]
  assign n56_I0_7_1_1 = n36_O_7_1_1; // @[Top.scala 190:12]
  assign n56_I0_7_1_2 = n36_O_7_1_2; // @[Top.scala 190:12]
  assign n56_I0_8_0_0 = n36_O_8_0_0; // @[Top.scala 190:12]
  assign n56_I0_8_0_1 = n36_O_8_0_1; // @[Top.scala 190:12]
  assign n56_I0_8_0_2 = n36_O_8_0_2; // @[Top.scala 190:12]
  assign n56_I0_8_1_0 = n36_O_8_1_0; // @[Top.scala 190:12]
  assign n56_I0_8_1_1 = n36_O_8_1_1; // @[Top.scala 190:12]
  assign n56_I0_8_1_2 = n36_O_8_1_2; // @[Top.scala 190:12]
  assign n56_I0_9_0_0 = n36_O_9_0_0; // @[Top.scala 190:12]
  assign n56_I0_9_0_1 = n36_O_9_0_1; // @[Top.scala 190:12]
  assign n56_I0_9_0_2 = n36_O_9_0_2; // @[Top.scala 190:12]
  assign n56_I0_9_1_0 = n36_O_9_1_0; // @[Top.scala 190:12]
  assign n56_I0_9_1_1 = n36_O_9_1_1; // @[Top.scala 190:12]
  assign n56_I0_9_1_2 = n36_O_9_1_2; // @[Top.scala 190:12]
  assign n56_I0_10_0_0 = n36_O_10_0_0; // @[Top.scala 190:12]
  assign n56_I0_10_0_1 = n36_O_10_0_1; // @[Top.scala 190:12]
  assign n56_I0_10_0_2 = n36_O_10_0_2; // @[Top.scala 190:12]
  assign n56_I0_10_1_0 = n36_O_10_1_0; // @[Top.scala 190:12]
  assign n56_I0_10_1_1 = n36_O_10_1_1; // @[Top.scala 190:12]
  assign n56_I0_10_1_2 = n36_O_10_1_2; // @[Top.scala 190:12]
  assign n56_I0_11_0_0 = n36_O_11_0_0; // @[Top.scala 190:12]
  assign n56_I0_11_0_1 = n36_O_11_0_1; // @[Top.scala 190:12]
  assign n56_I0_11_0_2 = n36_O_11_0_2; // @[Top.scala 190:12]
  assign n56_I0_11_1_0 = n36_O_11_1_0; // @[Top.scala 190:12]
  assign n56_I0_11_1_1 = n36_O_11_1_1; // @[Top.scala 190:12]
  assign n56_I0_11_1_2 = n36_O_11_1_2; // @[Top.scala 190:12]
  assign n56_I0_12_0_0 = n36_O_12_0_0; // @[Top.scala 190:12]
  assign n56_I0_12_0_1 = n36_O_12_0_1; // @[Top.scala 190:12]
  assign n56_I0_12_0_2 = n36_O_12_0_2; // @[Top.scala 190:12]
  assign n56_I0_12_1_0 = n36_O_12_1_0; // @[Top.scala 190:12]
  assign n56_I0_12_1_1 = n36_O_12_1_1; // @[Top.scala 190:12]
  assign n56_I0_12_1_2 = n36_O_12_1_2; // @[Top.scala 190:12]
  assign n56_I0_13_0_0 = n36_O_13_0_0; // @[Top.scala 190:12]
  assign n56_I0_13_0_1 = n36_O_13_0_1; // @[Top.scala 190:12]
  assign n56_I0_13_0_2 = n36_O_13_0_2; // @[Top.scala 190:12]
  assign n56_I0_13_1_0 = n36_O_13_1_0; // @[Top.scala 190:12]
  assign n56_I0_13_1_1 = n36_O_13_1_1; // @[Top.scala 190:12]
  assign n56_I0_13_1_2 = n36_O_13_1_2; // @[Top.scala 190:12]
  assign n56_I0_14_0_0 = n36_O_14_0_0; // @[Top.scala 190:12]
  assign n56_I0_14_0_1 = n36_O_14_0_1; // @[Top.scala 190:12]
  assign n56_I0_14_0_2 = n36_O_14_0_2; // @[Top.scala 190:12]
  assign n56_I0_14_1_0 = n36_O_14_1_0; // @[Top.scala 190:12]
  assign n56_I0_14_1_1 = n36_O_14_1_1; // @[Top.scala 190:12]
  assign n56_I0_14_1_2 = n36_O_14_1_2; // @[Top.scala 190:12]
  assign n56_I0_15_0_0 = n36_O_15_0_0; // @[Top.scala 190:12]
  assign n56_I0_15_0_1 = n36_O_15_0_1; // @[Top.scala 190:12]
  assign n56_I0_15_0_2 = n36_O_15_0_2; // @[Top.scala 190:12]
  assign n56_I0_15_1_0 = n36_O_15_1_0; // @[Top.scala 190:12]
  assign n56_I0_15_1_1 = n36_O_15_1_1; // @[Top.scala 190:12]
  assign n56_I0_15_1_2 = n36_O_15_1_2; // @[Top.scala 190:12]
  assign n56_I1_0_0 = n55_O_0_0; // @[Top.scala 191:12]
  assign n56_I1_0_1 = n55_O_0_1; // @[Top.scala 191:12]
  assign n56_I1_0_2 = n55_O_0_2; // @[Top.scala 191:12]
  assign n56_I1_1_0 = n55_O_1_0; // @[Top.scala 191:12]
  assign n56_I1_1_1 = n55_O_1_1; // @[Top.scala 191:12]
  assign n56_I1_1_2 = n55_O_1_2; // @[Top.scala 191:12]
  assign n56_I1_2_0 = n55_O_2_0; // @[Top.scala 191:12]
  assign n56_I1_2_1 = n55_O_2_1; // @[Top.scala 191:12]
  assign n56_I1_2_2 = n55_O_2_2; // @[Top.scala 191:12]
  assign n56_I1_3_0 = n55_O_3_0; // @[Top.scala 191:12]
  assign n56_I1_3_1 = n55_O_3_1; // @[Top.scala 191:12]
  assign n56_I1_3_2 = n55_O_3_2; // @[Top.scala 191:12]
  assign n56_I1_4_0 = n55_O_4_0; // @[Top.scala 191:12]
  assign n56_I1_4_1 = n55_O_4_1; // @[Top.scala 191:12]
  assign n56_I1_4_2 = n55_O_4_2; // @[Top.scala 191:12]
  assign n56_I1_5_0 = n55_O_5_0; // @[Top.scala 191:12]
  assign n56_I1_5_1 = n55_O_5_1; // @[Top.scala 191:12]
  assign n56_I1_5_2 = n55_O_5_2; // @[Top.scala 191:12]
  assign n56_I1_6_0 = n55_O_6_0; // @[Top.scala 191:12]
  assign n56_I1_6_1 = n55_O_6_1; // @[Top.scala 191:12]
  assign n56_I1_6_2 = n55_O_6_2; // @[Top.scala 191:12]
  assign n56_I1_7_0 = n55_O_7_0; // @[Top.scala 191:12]
  assign n56_I1_7_1 = n55_O_7_1; // @[Top.scala 191:12]
  assign n56_I1_7_2 = n55_O_7_2; // @[Top.scala 191:12]
  assign n56_I1_8_0 = n55_O_8_0; // @[Top.scala 191:12]
  assign n56_I1_8_1 = n55_O_8_1; // @[Top.scala 191:12]
  assign n56_I1_8_2 = n55_O_8_2; // @[Top.scala 191:12]
  assign n56_I1_9_0 = n55_O_9_0; // @[Top.scala 191:12]
  assign n56_I1_9_1 = n55_O_9_1; // @[Top.scala 191:12]
  assign n56_I1_9_2 = n55_O_9_2; // @[Top.scala 191:12]
  assign n56_I1_10_0 = n55_O_10_0; // @[Top.scala 191:12]
  assign n56_I1_10_1 = n55_O_10_1; // @[Top.scala 191:12]
  assign n56_I1_10_2 = n55_O_10_2; // @[Top.scala 191:12]
  assign n56_I1_11_0 = n55_O_11_0; // @[Top.scala 191:12]
  assign n56_I1_11_1 = n55_O_11_1; // @[Top.scala 191:12]
  assign n56_I1_11_2 = n55_O_11_2; // @[Top.scala 191:12]
  assign n56_I1_12_0 = n55_O_12_0; // @[Top.scala 191:12]
  assign n56_I1_12_1 = n55_O_12_1; // @[Top.scala 191:12]
  assign n56_I1_12_2 = n55_O_12_2; // @[Top.scala 191:12]
  assign n56_I1_13_0 = n55_O_13_0; // @[Top.scala 191:12]
  assign n56_I1_13_1 = n55_O_13_1; // @[Top.scala 191:12]
  assign n56_I1_13_2 = n55_O_13_2; // @[Top.scala 191:12]
  assign n56_I1_14_0 = n55_O_14_0; // @[Top.scala 191:12]
  assign n56_I1_14_1 = n55_O_14_1; // @[Top.scala 191:12]
  assign n56_I1_14_2 = n55_O_14_2; // @[Top.scala 191:12]
  assign n56_I1_15_0 = n55_O_15_0; // @[Top.scala 191:12]
  assign n56_I1_15_1 = n55_O_15_1; // @[Top.scala 191:12]
  assign n56_I1_15_2 = n55_O_15_2; // @[Top.scala 191:12]
  assign n60_valid_up = n56_valid_down; // @[Top.scala 195:18]
  assign n60_I_0_0_0 = n56_O_0_0_0; // @[Top.scala 194:11]
  assign n60_I_0_0_1 = n56_O_0_0_1; // @[Top.scala 194:11]
  assign n60_I_0_0_2 = n56_O_0_0_2; // @[Top.scala 194:11]
  assign n60_I_0_1_0 = n56_O_0_1_0; // @[Top.scala 194:11]
  assign n60_I_0_1_1 = n56_O_0_1_1; // @[Top.scala 194:11]
  assign n60_I_0_1_2 = n56_O_0_1_2; // @[Top.scala 194:11]
  assign n60_I_0_2_0 = n56_O_0_2_0; // @[Top.scala 194:11]
  assign n60_I_0_2_1 = n56_O_0_2_1; // @[Top.scala 194:11]
  assign n60_I_0_2_2 = n56_O_0_2_2; // @[Top.scala 194:11]
  assign n60_I_1_0_0 = n56_O_1_0_0; // @[Top.scala 194:11]
  assign n60_I_1_0_1 = n56_O_1_0_1; // @[Top.scala 194:11]
  assign n60_I_1_0_2 = n56_O_1_0_2; // @[Top.scala 194:11]
  assign n60_I_1_1_0 = n56_O_1_1_0; // @[Top.scala 194:11]
  assign n60_I_1_1_1 = n56_O_1_1_1; // @[Top.scala 194:11]
  assign n60_I_1_1_2 = n56_O_1_1_2; // @[Top.scala 194:11]
  assign n60_I_1_2_0 = n56_O_1_2_0; // @[Top.scala 194:11]
  assign n60_I_1_2_1 = n56_O_1_2_1; // @[Top.scala 194:11]
  assign n60_I_1_2_2 = n56_O_1_2_2; // @[Top.scala 194:11]
  assign n60_I_2_0_0 = n56_O_2_0_0; // @[Top.scala 194:11]
  assign n60_I_2_0_1 = n56_O_2_0_1; // @[Top.scala 194:11]
  assign n60_I_2_0_2 = n56_O_2_0_2; // @[Top.scala 194:11]
  assign n60_I_2_1_0 = n56_O_2_1_0; // @[Top.scala 194:11]
  assign n60_I_2_1_1 = n56_O_2_1_1; // @[Top.scala 194:11]
  assign n60_I_2_1_2 = n56_O_2_1_2; // @[Top.scala 194:11]
  assign n60_I_2_2_0 = n56_O_2_2_0; // @[Top.scala 194:11]
  assign n60_I_2_2_1 = n56_O_2_2_1; // @[Top.scala 194:11]
  assign n60_I_2_2_2 = n56_O_2_2_2; // @[Top.scala 194:11]
  assign n60_I_3_0_0 = n56_O_3_0_0; // @[Top.scala 194:11]
  assign n60_I_3_0_1 = n56_O_3_0_1; // @[Top.scala 194:11]
  assign n60_I_3_0_2 = n56_O_3_0_2; // @[Top.scala 194:11]
  assign n60_I_3_1_0 = n56_O_3_1_0; // @[Top.scala 194:11]
  assign n60_I_3_1_1 = n56_O_3_1_1; // @[Top.scala 194:11]
  assign n60_I_3_1_2 = n56_O_3_1_2; // @[Top.scala 194:11]
  assign n60_I_3_2_0 = n56_O_3_2_0; // @[Top.scala 194:11]
  assign n60_I_3_2_1 = n56_O_3_2_1; // @[Top.scala 194:11]
  assign n60_I_3_2_2 = n56_O_3_2_2; // @[Top.scala 194:11]
  assign n60_I_4_0_0 = n56_O_4_0_0; // @[Top.scala 194:11]
  assign n60_I_4_0_1 = n56_O_4_0_1; // @[Top.scala 194:11]
  assign n60_I_4_0_2 = n56_O_4_0_2; // @[Top.scala 194:11]
  assign n60_I_4_1_0 = n56_O_4_1_0; // @[Top.scala 194:11]
  assign n60_I_4_1_1 = n56_O_4_1_1; // @[Top.scala 194:11]
  assign n60_I_4_1_2 = n56_O_4_1_2; // @[Top.scala 194:11]
  assign n60_I_4_2_0 = n56_O_4_2_0; // @[Top.scala 194:11]
  assign n60_I_4_2_1 = n56_O_4_2_1; // @[Top.scala 194:11]
  assign n60_I_4_2_2 = n56_O_4_2_2; // @[Top.scala 194:11]
  assign n60_I_5_0_0 = n56_O_5_0_0; // @[Top.scala 194:11]
  assign n60_I_5_0_1 = n56_O_5_0_1; // @[Top.scala 194:11]
  assign n60_I_5_0_2 = n56_O_5_0_2; // @[Top.scala 194:11]
  assign n60_I_5_1_0 = n56_O_5_1_0; // @[Top.scala 194:11]
  assign n60_I_5_1_1 = n56_O_5_1_1; // @[Top.scala 194:11]
  assign n60_I_5_1_2 = n56_O_5_1_2; // @[Top.scala 194:11]
  assign n60_I_5_2_0 = n56_O_5_2_0; // @[Top.scala 194:11]
  assign n60_I_5_2_1 = n56_O_5_2_1; // @[Top.scala 194:11]
  assign n60_I_5_2_2 = n56_O_5_2_2; // @[Top.scala 194:11]
  assign n60_I_6_0_0 = n56_O_6_0_0; // @[Top.scala 194:11]
  assign n60_I_6_0_1 = n56_O_6_0_1; // @[Top.scala 194:11]
  assign n60_I_6_0_2 = n56_O_6_0_2; // @[Top.scala 194:11]
  assign n60_I_6_1_0 = n56_O_6_1_0; // @[Top.scala 194:11]
  assign n60_I_6_1_1 = n56_O_6_1_1; // @[Top.scala 194:11]
  assign n60_I_6_1_2 = n56_O_6_1_2; // @[Top.scala 194:11]
  assign n60_I_6_2_0 = n56_O_6_2_0; // @[Top.scala 194:11]
  assign n60_I_6_2_1 = n56_O_6_2_1; // @[Top.scala 194:11]
  assign n60_I_6_2_2 = n56_O_6_2_2; // @[Top.scala 194:11]
  assign n60_I_7_0_0 = n56_O_7_0_0; // @[Top.scala 194:11]
  assign n60_I_7_0_1 = n56_O_7_0_1; // @[Top.scala 194:11]
  assign n60_I_7_0_2 = n56_O_7_0_2; // @[Top.scala 194:11]
  assign n60_I_7_1_0 = n56_O_7_1_0; // @[Top.scala 194:11]
  assign n60_I_7_1_1 = n56_O_7_1_1; // @[Top.scala 194:11]
  assign n60_I_7_1_2 = n56_O_7_1_2; // @[Top.scala 194:11]
  assign n60_I_7_2_0 = n56_O_7_2_0; // @[Top.scala 194:11]
  assign n60_I_7_2_1 = n56_O_7_2_1; // @[Top.scala 194:11]
  assign n60_I_7_2_2 = n56_O_7_2_2; // @[Top.scala 194:11]
  assign n60_I_8_0_0 = n56_O_8_0_0; // @[Top.scala 194:11]
  assign n60_I_8_0_1 = n56_O_8_0_1; // @[Top.scala 194:11]
  assign n60_I_8_0_2 = n56_O_8_0_2; // @[Top.scala 194:11]
  assign n60_I_8_1_0 = n56_O_8_1_0; // @[Top.scala 194:11]
  assign n60_I_8_1_1 = n56_O_8_1_1; // @[Top.scala 194:11]
  assign n60_I_8_1_2 = n56_O_8_1_2; // @[Top.scala 194:11]
  assign n60_I_8_2_0 = n56_O_8_2_0; // @[Top.scala 194:11]
  assign n60_I_8_2_1 = n56_O_8_2_1; // @[Top.scala 194:11]
  assign n60_I_8_2_2 = n56_O_8_2_2; // @[Top.scala 194:11]
  assign n60_I_9_0_0 = n56_O_9_0_0; // @[Top.scala 194:11]
  assign n60_I_9_0_1 = n56_O_9_0_1; // @[Top.scala 194:11]
  assign n60_I_9_0_2 = n56_O_9_0_2; // @[Top.scala 194:11]
  assign n60_I_9_1_0 = n56_O_9_1_0; // @[Top.scala 194:11]
  assign n60_I_9_1_1 = n56_O_9_1_1; // @[Top.scala 194:11]
  assign n60_I_9_1_2 = n56_O_9_1_2; // @[Top.scala 194:11]
  assign n60_I_9_2_0 = n56_O_9_2_0; // @[Top.scala 194:11]
  assign n60_I_9_2_1 = n56_O_9_2_1; // @[Top.scala 194:11]
  assign n60_I_9_2_2 = n56_O_9_2_2; // @[Top.scala 194:11]
  assign n60_I_10_0_0 = n56_O_10_0_0; // @[Top.scala 194:11]
  assign n60_I_10_0_1 = n56_O_10_0_1; // @[Top.scala 194:11]
  assign n60_I_10_0_2 = n56_O_10_0_2; // @[Top.scala 194:11]
  assign n60_I_10_1_0 = n56_O_10_1_0; // @[Top.scala 194:11]
  assign n60_I_10_1_1 = n56_O_10_1_1; // @[Top.scala 194:11]
  assign n60_I_10_1_2 = n56_O_10_1_2; // @[Top.scala 194:11]
  assign n60_I_10_2_0 = n56_O_10_2_0; // @[Top.scala 194:11]
  assign n60_I_10_2_1 = n56_O_10_2_1; // @[Top.scala 194:11]
  assign n60_I_10_2_2 = n56_O_10_2_2; // @[Top.scala 194:11]
  assign n60_I_11_0_0 = n56_O_11_0_0; // @[Top.scala 194:11]
  assign n60_I_11_0_1 = n56_O_11_0_1; // @[Top.scala 194:11]
  assign n60_I_11_0_2 = n56_O_11_0_2; // @[Top.scala 194:11]
  assign n60_I_11_1_0 = n56_O_11_1_0; // @[Top.scala 194:11]
  assign n60_I_11_1_1 = n56_O_11_1_1; // @[Top.scala 194:11]
  assign n60_I_11_1_2 = n56_O_11_1_2; // @[Top.scala 194:11]
  assign n60_I_11_2_0 = n56_O_11_2_0; // @[Top.scala 194:11]
  assign n60_I_11_2_1 = n56_O_11_2_1; // @[Top.scala 194:11]
  assign n60_I_11_2_2 = n56_O_11_2_2; // @[Top.scala 194:11]
  assign n60_I_12_0_0 = n56_O_12_0_0; // @[Top.scala 194:11]
  assign n60_I_12_0_1 = n56_O_12_0_1; // @[Top.scala 194:11]
  assign n60_I_12_0_2 = n56_O_12_0_2; // @[Top.scala 194:11]
  assign n60_I_12_1_0 = n56_O_12_1_0; // @[Top.scala 194:11]
  assign n60_I_12_1_1 = n56_O_12_1_1; // @[Top.scala 194:11]
  assign n60_I_12_1_2 = n56_O_12_1_2; // @[Top.scala 194:11]
  assign n60_I_12_2_0 = n56_O_12_2_0; // @[Top.scala 194:11]
  assign n60_I_12_2_1 = n56_O_12_2_1; // @[Top.scala 194:11]
  assign n60_I_12_2_2 = n56_O_12_2_2; // @[Top.scala 194:11]
  assign n60_I_13_0_0 = n56_O_13_0_0; // @[Top.scala 194:11]
  assign n60_I_13_0_1 = n56_O_13_0_1; // @[Top.scala 194:11]
  assign n60_I_13_0_2 = n56_O_13_0_2; // @[Top.scala 194:11]
  assign n60_I_13_1_0 = n56_O_13_1_0; // @[Top.scala 194:11]
  assign n60_I_13_1_1 = n56_O_13_1_1; // @[Top.scala 194:11]
  assign n60_I_13_1_2 = n56_O_13_1_2; // @[Top.scala 194:11]
  assign n60_I_13_2_0 = n56_O_13_2_0; // @[Top.scala 194:11]
  assign n60_I_13_2_1 = n56_O_13_2_1; // @[Top.scala 194:11]
  assign n60_I_13_2_2 = n56_O_13_2_2; // @[Top.scala 194:11]
  assign n60_I_14_0_0 = n56_O_14_0_0; // @[Top.scala 194:11]
  assign n60_I_14_0_1 = n56_O_14_0_1; // @[Top.scala 194:11]
  assign n60_I_14_0_2 = n56_O_14_0_2; // @[Top.scala 194:11]
  assign n60_I_14_1_0 = n56_O_14_1_0; // @[Top.scala 194:11]
  assign n60_I_14_1_1 = n56_O_14_1_1; // @[Top.scala 194:11]
  assign n60_I_14_1_2 = n56_O_14_1_2; // @[Top.scala 194:11]
  assign n60_I_14_2_0 = n56_O_14_2_0; // @[Top.scala 194:11]
  assign n60_I_14_2_1 = n56_O_14_2_1; // @[Top.scala 194:11]
  assign n60_I_14_2_2 = n56_O_14_2_2; // @[Top.scala 194:11]
  assign n60_I_15_0_0 = n56_O_15_0_0; // @[Top.scala 194:11]
  assign n60_I_15_0_1 = n56_O_15_0_1; // @[Top.scala 194:11]
  assign n60_I_15_0_2 = n56_O_15_0_2; // @[Top.scala 194:11]
  assign n60_I_15_1_0 = n56_O_15_1_0; // @[Top.scala 194:11]
  assign n60_I_15_1_1 = n56_O_15_1_1; // @[Top.scala 194:11]
  assign n60_I_15_1_2 = n56_O_15_1_2; // @[Top.scala 194:11]
  assign n60_I_15_2_0 = n56_O_15_2_0; // @[Top.scala 194:11]
  assign n60_I_15_2_1 = n56_O_15_2_1; // @[Top.scala 194:11]
  assign n60_I_15_2_2 = n56_O_15_2_2; // @[Top.scala 194:11]
  assign n65_valid_up = n60_valid_down; // @[Top.scala 198:18]
  assign n65_I_0_0_0_0 = n60_O_0_0_0_0; // @[Top.scala 197:11]
  assign n65_I_0_0_0_1 = n60_O_0_0_0_1; // @[Top.scala 197:11]
  assign n65_I_0_0_0_2 = n60_O_0_0_0_2; // @[Top.scala 197:11]
  assign n65_I_0_0_1_0 = n60_O_0_0_1_0; // @[Top.scala 197:11]
  assign n65_I_0_0_1_1 = n60_O_0_0_1_1; // @[Top.scala 197:11]
  assign n65_I_0_0_1_2 = n60_O_0_0_1_2; // @[Top.scala 197:11]
  assign n65_I_0_0_2_0 = n60_O_0_0_2_0; // @[Top.scala 197:11]
  assign n65_I_0_0_2_1 = n60_O_0_0_2_1; // @[Top.scala 197:11]
  assign n65_I_0_0_2_2 = n60_O_0_0_2_2; // @[Top.scala 197:11]
  assign n65_I_1_0_0_0 = n60_O_1_0_0_0; // @[Top.scala 197:11]
  assign n65_I_1_0_0_1 = n60_O_1_0_0_1; // @[Top.scala 197:11]
  assign n65_I_1_0_0_2 = n60_O_1_0_0_2; // @[Top.scala 197:11]
  assign n65_I_1_0_1_0 = n60_O_1_0_1_0; // @[Top.scala 197:11]
  assign n65_I_1_0_1_1 = n60_O_1_0_1_1; // @[Top.scala 197:11]
  assign n65_I_1_0_1_2 = n60_O_1_0_1_2; // @[Top.scala 197:11]
  assign n65_I_1_0_2_0 = n60_O_1_0_2_0; // @[Top.scala 197:11]
  assign n65_I_1_0_2_1 = n60_O_1_0_2_1; // @[Top.scala 197:11]
  assign n65_I_1_0_2_2 = n60_O_1_0_2_2; // @[Top.scala 197:11]
  assign n65_I_2_0_0_0 = n60_O_2_0_0_0; // @[Top.scala 197:11]
  assign n65_I_2_0_0_1 = n60_O_2_0_0_1; // @[Top.scala 197:11]
  assign n65_I_2_0_0_2 = n60_O_2_0_0_2; // @[Top.scala 197:11]
  assign n65_I_2_0_1_0 = n60_O_2_0_1_0; // @[Top.scala 197:11]
  assign n65_I_2_0_1_1 = n60_O_2_0_1_1; // @[Top.scala 197:11]
  assign n65_I_2_0_1_2 = n60_O_2_0_1_2; // @[Top.scala 197:11]
  assign n65_I_2_0_2_0 = n60_O_2_0_2_0; // @[Top.scala 197:11]
  assign n65_I_2_0_2_1 = n60_O_2_0_2_1; // @[Top.scala 197:11]
  assign n65_I_2_0_2_2 = n60_O_2_0_2_2; // @[Top.scala 197:11]
  assign n65_I_3_0_0_0 = n60_O_3_0_0_0; // @[Top.scala 197:11]
  assign n65_I_3_0_0_1 = n60_O_3_0_0_1; // @[Top.scala 197:11]
  assign n65_I_3_0_0_2 = n60_O_3_0_0_2; // @[Top.scala 197:11]
  assign n65_I_3_0_1_0 = n60_O_3_0_1_0; // @[Top.scala 197:11]
  assign n65_I_3_0_1_1 = n60_O_3_0_1_1; // @[Top.scala 197:11]
  assign n65_I_3_0_1_2 = n60_O_3_0_1_2; // @[Top.scala 197:11]
  assign n65_I_3_0_2_0 = n60_O_3_0_2_0; // @[Top.scala 197:11]
  assign n65_I_3_0_2_1 = n60_O_3_0_2_1; // @[Top.scala 197:11]
  assign n65_I_3_0_2_2 = n60_O_3_0_2_2; // @[Top.scala 197:11]
  assign n65_I_4_0_0_0 = n60_O_4_0_0_0; // @[Top.scala 197:11]
  assign n65_I_4_0_0_1 = n60_O_4_0_0_1; // @[Top.scala 197:11]
  assign n65_I_4_0_0_2 = n60_O_4_0_0_2; // @[Top.scala 197:11]
  assign n65_I_4_0_1_0 = n60_O_4_0_1_0; // @[Top.scala 197:11]
  assign n65_I_4_0_1_1 = n60_O_4_0_1_1; // @[Top.scala 197:11]
  assign n65_I_4_0_1_2 = n60_O_4_0_1_2; // @[Top.scala 197:11]
  assign n65_I_4_0_2_0 = n60_O_4_0_2_0; // @[Top.scala 197:11]
  assign n65_I_4_0_2_1 = n60_O_4_0_2_1; // @[Top.scala 197:11]
  assign n65_I_4_0_2_2 = n60_O_4_0_2_2; // @[Top.scala 197:11]
  assign n65_I_5_0_0_0 = n60_O_5_0_0_0; // @[Top.scala 197:11]
  assign n65_I_5_0_0_1 = n60_O_5_0_0_1; // @[Top.scala 197:11]
  assign n65_I_5_0_0_2 = n60_O_5_0_0_2; // @[Top.scala 197:11]
  assign n65_I_5_0_1_0 = n60_O_5_0_1_0; // @[Top.scala 197:11]
  assign n65_I_5_0_1_1 = n60_O_5_0_1_1; // @[Top.scala 197:11]
  assign n65_I_5_0_1_2 = n60_O_5_0_1_2; // @[Top.scala 197:11]
  assign n65_I_5_0_2_0 = n60_O_5_0_2_0; // @[Top.scala 197:11]
  assign n65_I_5_0_2_1 = n60_O_5_0_2_1; // @[Top.scala 197:11]
  assign n65_I_5_0_2_2 = n60_O_5_0_2_2; // @[Top.scala 197:11]
  assign n65_I_6_0_0_0 = n60_O_6_0_0_0; // @[Top.scala 197:11]
  assign n65_I_6_0_0_1 = n60_O_6_0_0_1; // @[Top.scala 197:11]
  assign n65_I_6_0_0_2 = n60_O_6_0_0_2; // @[Top.scala 197:11]
  assign n65_I_6_0_1_0 = n60_O_6_0_1_0; // @[Top.scala 197:11]
  assign n65_I_6_0_1_1 = n60_O_6_0_1_1; // @[Top.scala 197:11]
  assign n65_I_6_0_1_2 = n60_O_6_0_1_2; // @[Top.scala 197:11]
  assign n65_I_6_0_2_0 = n60_O_6_0_2_0; // @[Top.scala 197:11]
  assign n65_I_6_0_2_1 = n60_O_6_0_2_1; // @[Top.scala 197:11]
  assign n65_I_6_0_2_2 = n60_O_6_0_2_2; // @[Top.scala 197:11]
  assign n65_I_7_0_0_0 = n60_O_7_0_0_0; // @[Top.scala 197:11]
  assign n65_I_7_0_0_1 = n60_O_7_0_0_1; // @[Top.scala 197:11]
  assign n65_I_7_0_0_2 = n60_O_7_0_0_2; // @[Top.scala 197:11]
  assign n65_I_7_0_1_0 = n60_O_7_0_1_0; // @[Top.scala 197:11]
  assign n65_I_7_0_1_1 = n60_O_7_0_1_1; // @[Top.scala 197:11]
  assign n65_I_7_0_1_2 = n60_O_7_0_1_2; // @[Top.scala 197:11]
  assign n65_I_7_0_2_0 = n60_O_7_0_2_0; // @[Top.scala 197:11]
  assign n65_I_7_0_2_1 = n60_O_7_0_2_1; // @[Top.scala 197:11]
  assign n65_I_7_0_2_2 = n60_O_7_0_2_2; // @[Top.scala 197:11]
  assign n65_I_8_0_0_0 = n60_O_8_0_0_0; // @[Top.scala 197:11]
  assign n65_I_8_0_0_1 = n60_O_8_0_0_1; // @[Top.scala 197:11]
  assign n65_I_8_0_0_2 = n60_O_8_0_0_2; // @[Top.scala 197:11]
  assign n65_I_8_0_1_0 = n60_O_8_0_1_0; // @[Top.scala 197:11]
  assign n65_I_8_0_1_1 = n60_O_8_0_1_1; // @[Top.scala 197:11]
  assign n65_I_8_0_1_2 = n60_O_8_0_1_2; // @[Top.scala 197:11]
  assign n65_I_8_0_2_0 = n60_O_8_0_2_0; // @[Top.scala 197:11]
  assign n65_I_8_0_2_1 = n60_O_8_0_2_1; // @[Top.scala 197:11]
  assign n65_I_8_0_2_2 = n60_O_8_0_2_2; // @[Top.scala 197:11]
  assign n65_I_9_0_0_0 = n60_O_9_0_0_0; // @[Top.scala 197:11]
  assign n65_I_9_0_0_1 = n60_O_9_0_0_1; // @[Top.scala 197:11]
  assign n65_I_9_0_0_2 = n60_O_9_0_0_2; // @[Top.scala 197:11]
  assign n65_I_9_0_1_0 = n60_O_9_0_1_0; // @[Top.scala 197:11]
  assign n65_I_9_0_1_1 = n60_O_9_0_1_1; // @[Top.scala 197:11]
  assign n65_I_9_0_1_2 = n60_O_9_0_1_2; // @[Top.scala 197:11]
  assign n65_I_9_0_2_0 = n60_O_9_0_2_0; // @[Top.scala 197:11]
  assign n65_I_9_0_2_1 = n60_O_9_0_2_1; // @[Top.scala 197:11]
  assign n65_I_9_0_2_2 = n60_O_9_0_2_2; // @[Top.scala 197:11]
  assign n65_I_10_0_0_0 = n60_O_10_0_0_0; // @[Top.scala 197:11]
  assign n65_I_10_0_0_1 = n60_O_10_0_0_1; // @[Top.scala 197:11]
  assign n65_I_10_0_0_2 = n60_O_10_0_0_2; // @[Top.scala 197:11]
  assign n65_I_10_0_1_0 = n60_O_10_0_1_0; // @[Top.scala 197:11]
  assign n65_I_10_0_1_1 = n60_O_10_0_1_1; // @[Top.scala 197:11]
  assign n65_I_10_0_1_2 = n60_O_10_0_1_2; // @[Top.scala 197:11]
  assign n65_I_10_0_2_0 = n60_O_10_0_2_0; // @[Top.scala 197:11]
  assign n65_I_10_0_2_1 = n60_O_10_0_2_1; // @[Top.scala 197:11]
  assign n65_I_10_0_2_2 = n60_O_10_0_2_2; // @[Top.scala 197:11]
  assign n65_I_11_0_0_0 = n60_O_11_0_0_0; // @[Top.scala 197:11]
  assign n65_I_11_0_0_1 = n60_O_11_0_0_1; // @[Top.scala 197:11]
  assign n65_I_11_0_0_2 = n60_O_11_0_0_2; // @[Top.scala 197:11]
  assign n65_I_11_0_1_0 = n60_O_11_0_1_0; // @[Top.scala 197:11]
  assign n65_I_11_0_1_1 = n60_O_11_0_1_1; // @[Top.scala 197:11]
  assign n65_I_11_0_1_2 = n60_O_11_0_1_2; // @[Top.scala 197:11]
  assign n65_I_11_0_2_0 = n60_O_11_0_2_0; // @[Top.scala 197:11]
  assign n65_I_11_0_2_1 = n60_O_11_0_2_1; // @[Top.scala 197:11]
  assign n65_I_11_0_2_2 = n60_O_11_0_2_2; // @[Top.scala 197:11]
  assign n65_I_12_0_0_0 = n60_O_12_0_0_0; // @[Top.scala 197:11]
  assign n65_I_12_0_0_1 = n60_O_12_0_0_1; // @[Top.scala 197:11]
  assign n65_I_12_0_0_2 = n60_O_12_0_0_2; // @[Top.scala 197:11]
  assign n65_I_12_0_1_0 = n60_O_12_0_1_0; // @[Top.scala 197:11]
  assign n65_I_12_0_1_1 = n60_O_12_0_1_1; // @[Top.scala 197:11]
  assign n65_I_12_0_1_2 = n60_O_12_0_1_2; // @[Top.scala 197:11]
  assign n65_I_12_0_2_0 = n60_O_12_0_2_0; // @[Top.scala 197:11]
  assign n65_I_12_0_2_1 = n60_O_12_0_2_1; // @[Top.scala 197:11]
  assign n65_I_12_0_2_2 = n60_O_12_0_2_2; // @[Top.scala 197:11]
  assign n65_I_13_0_0_0 = n60_O_13_0_0_0; // @[Top.scala 197:11]
  assign n65_I_13_0_0_1 = n60_O_13_0_0_1; // @[Top.scala 197:11]
  assign n65_I_13_0_0_2 = n60_O_13_0_0_2; // @[Top.scala 197:11]
  assign n65_I_13_0_1_0 = n60_O_13_0_1_0; // @[Top.scala 197:11]
  assign n65_I_13_0_1_1 = n60_O_13_0_1_1; // @[Top.scala 197:11]
  assign n65_I_13_0_1_2 = n60_O_13_0_1_2; // @[Top.scala 197:11]
  assign n65_I_13_0_2_0 = n60_O_13_0_2_0; // @[Top.scala 197:11]
  assign n65_I_13_0_2_1 = n60_O_13_0_2_1; // @[Top.scala 197:11]
  assign n65_I_13_0_2_2 = n60_O_13_0_2_2; // @[Top.scala 197:11]
  assign n65_I_14_0_0_0 = n60_O_14_0_0_0; // @[Top.scala 197:11]
  assign n65_I_14_0_0_1 = n60_O_14_0_0_1; // @[Top.scala 197:11]
  assign n65_I_14_0_0_2 = n60_O_14_0_0_2; // @[Top.scala 197:11]
  assign n65_I_14_0_1_0 = n60_O_14_0_1_0; // @[Top.scala 197:11]
  assign n65_I_14_0_1_1 = n60_O_14_0_1_1; // @[Top.scala 197:11]
  assign n65_I_14_0_1_2 = n60_O_14_0_1_2; // @[Top.scala 197:11]
  assign n65_I_14_0_2_0 = n60_O_14_0_2_0; // @[Top.scala 197:11]
  assign n65_I_14_0_2_1 = n60_O_14_0_2_1; // @[Top.scala 197:11]
  assign n65_I_14_0_2_2 = n60_O_14_0_2_2; // @[Top.scala 197:11]
  assign n65_I_15_0_0_0 = n60_O_15_0_0_0; // @[Top.scala 197:11]
  assign n65_I_15_0_0_1 = n60_O_15_0_0_1; // @[Top.scala 197:11]
  assign n65_I_15_0_0_2 = n60_O_15_0_0_2; // @[Top.scala 197:11]
  assign n65_I_15_0_1_0 = n60_O_15_0_1_0; // @[Top.scala 197:11]
  assign n65_I_15_0_1_1 = n60_O_15_0_1_1; // @[Top.scala 197:11]
  assign n65_I_15_0_1_2 = n60_O_15_0_1_2; // @[Top.scala 197:11]
  assign n65_I_15_0_2_0 = n60_O_15_0_2_0; // @[Top.scala 197:11]
  assign n65_I_15_0_2_1 = n60_O_15_0_2_1; // @[Top.scala 197:11]
  assign n65_I_15_0_2_2 = n60_O_15_0_2_2; // @[Top.scala 197:11]
  assign n105_clock = clock;
  assign n105_reset = reset;
  assign n105_valid_up = n65_valid_down; // @[Top.scala 201:19]
  assign n105_I_0_0_0 = n65_O_0_0_0; // @[Top.scala 200:12]
  assign n105_I_0_0_1 = n65_O_0_0_1; // @[Top.scala 200:12]
  assign n105_I_0_0_2 = n65_O_0_0_2; // @[Top.scala 200:12]
  assign n105_I_0_1_0 = n65_O_0_1_0; // @[Top.scala 200:12]
  assign n105_I_0_1_1 = n65_O_0_1_1; // @[Top.scala 200:12]
  assign n105_I_0_1_2 = n65_O_0_1_2; // @[Top.scala 200:12]
  assign n105_I_0_2_0 = n65_O_0_2_0; // @[Top.scala 200:12]
  assign n105_I_0_2_1 = n65_O_0_2_1; // @[Top.scala 200:12]
  assign n105_I_0_2_2 = n65_O_0_2_2; // @[Top.scala 200:12]
  assign n105_I_1_0_0 = n65_O_1_0_0; // @[Top.scala 200:12]
  assign n105_I_1_0_1 = n65_O_1_0_1; // @[Top.scala 200:12]
  assign n105_I_1_0_2 = n65_O_1_0_2; // @[Top.scala 200:12]
  assign n105_I_1_1_0 = n65_O_1_1_0; // @[Top.scala 200:12]
  assign n105_I_1_1_1 = n65_O_1_1_1; // @[Top.scala 200:12]
  assign n105_I_1_1_2 = n65_O_1_1_2; // @[Top.scala 200:12]
  assign n105_I_1_2_0 = n65_O_1_2_0; // @[Top.scala 200:12]
  assign n105_I_1_2_1 = n65_O_1_2_1; // @[Top.scala 200:12]
  assign n105_I_1_2_2 = n65_O_1_2_2; // @[Top.scala 200:12]
  assign n105_I_2_0_0 = n65_O_2_0_0; // @[Top.scala 200:12]
  assign n105_I_2_0_1 = n65_O_2_0_1; // @[Top.scala 200:12]
  assign n105_I_2_0_2 = n65_O_2_0_2; // @[Top.scala 200:12]
  assign n105_I_2_1_0 = n65_O_2_1_0; // @[Top.scala 200:12]
  assign n105_I_2_1_1 = n65_O_2_1_1; // @[Top.scala 200:12]
  assign n105_I_2_1_2 = n65_O_2_1_2; // @[Top.scala 200:12]
  assign n105_I_2_2_0 = n65_O_2_2_0; // @[Top.scala 200:12]
  assign n105_I_2_2_1 = n65_O_2_2_1; // @[Top.scala 200:12]
  assign n105_I_2_2_2 = n65_O_2_2_2; // @[Top.scala 200:12]
  assign n105_I_3_0_0 = n65_O_3_0_0; // @[Top.scala 200:12]
  assign n105_I_3_0_1 = n65_O_3_0_1; // @[Top.scala 200:12]
  assign n105_I_3_0_2 = n65_O_3_0_2; // @[Top.scala 200:12]
  assign n105_I_3_1_0 = n65_O_3_1_0; // @[Top.scala 200:12]
  assign n105_I_3_1_1 = n65_O_3_1_1; // @[Top.scala 200:12]
  assign n105_I_3_1_2 = n65_O_3_1_2; // @[Top.scala 200:12]
  assign n105_I_3_2_0 = n65_O_3_2_0; // @[Top.scala 200:12]
  assign n105_I_3_2_1 = n65_O_3_2_1; // @[Top.scala 200:12]
  assign n105_I_3_2_2 = n65_O_3_2_2; // @[Top.scala 200:12]
  assign n105_I_4_0_0 = n65_O_4_0_0; // @[Top.scala 200:12]
  assign n105_I_4_0_1 = n65_O_4_0_1; // @[Top.scala 200:12]
  assign n105_I_4_0_2 = n65_O_4_0_2; // @[Top.scala 200:12]
  assign n105_I_4_1_0 = n65_O_4_1_0; // @[Top.scala 200:12]
  assign n105_I_4_1_1 = n65_O_4_1_1; // @[Top.scala 200:12]
  assign n105_I_4_1_2 = n65_O_4_1_2; // @[Top.scala 200:12]
  assign n105_I_4_2_0 = n65_O_4_2_0; // @[Top.scala 200:12]
  assign n105_I_4_2_1 = n65_O_4_2_1; // @[Top.scala 200:12]
  assign n105_I_4_2_2 = n65_O_4_2_2; // @[Top.scala 200:12]
  assign n105_I_5_0_0 = n65_O_5_0_0; // @[Top.scala 200:12]
  assign n105_I_5_0_1 = n65_O_5_0_1; // @[Top.scala 200:12]
  assign n105_I_5_0_2 = n65_O_5_0_2; // @[Top.scala 200:12]
  assign n105_I_5_1_0 = n65_O_5_1_0; // @[Top.scala 200:12]
  assign n105_I_5_1_1 = n65_O_5_1_1; // @[Top.scala 200:12]
  assign n105_I_5_1_2 = n65_O_5_1_2; // @[Top.scala 200:12]
  assign n105_I_5_2_0 = n65_O_5_2_0; // @[Top.scala 200:12]
  assign n105_I_5_2_1 = n65_O_5_2_1; // @[Top.scala 200:12]
  assign n105_I_5_2_2 = n65_O_5_2_2; // @[Top.scala 200:12]
  assign n105_I_6_0_0 = n65_O_6_0_0; // @[Top.scala 200:12]
  assign n105_I_6_0_1 = n65_O_6_0_1; // @[Top.scala 200:12]
  assign n105_I_6_0_2 = n65_O_6_0_2; // @[Top.scala 200:12]
  assign n105_I_6_1_0 = n65_O_6_1_0; // @[Top.scala 200:12]
  assign n105_I_6_1_1 = n65_O_6_1_1; // @[Top.scala 200:12]
  assign n105_I_6_1_2 = n65_O_6_1_2; // @[Top.scala 200:12]
  assign n105_I_6_2_0 = n65_O_6_2_0; // @[Top.scala 200:12]
  assign n105_I_6_2_1 = n65_O_6_2_1; // @[Top.scala 200:12]
  assign n105_I_6_2_2 = n65_O_6_2_2; // @[Top.scala 200:12]
  assign n105_I_7_0_0 = n65_O_7_0_0; // @[Top.scala 200:12]
  assign n105_I_7_0_1 = n65_O_7_0_1; // @[Top.scala 200:12]
  assign n105_I_7_0_2 = n65_O_7_0_2; // @[Top.scala 200:12]
  assign n105_I_7_1_0 = n65_O_7_1_0; // @[Top.scala 200:12]
  assign n105_I_7_1_1 = n65_O_7_1_1; // @[Top.scala 200:12]
  assign n105_I_7_1_2 = n65_O_7_1_2; // @[Top.scala 200:12]
  assign n105_I_7_2_0 = n65_O_7_2_0; // @[Top.scala 200:12]
  assign n105_I_7_2_1 = n65_O_7_2_1; // @[Top.scala 200:12]
  assign n105_I_7_2_2 = n65_O_7_2_2; // @[Top.scala 200:12]
  assign n105_I_8_0_0 = n65_O_8_0_0; // @[Top.scala 200:12]
  assign n105_I_8_0_1 = n65_O_8_0_1; // @[Top.scala 200:12]
  assign n105_I_8_0_2 = n65_O_8_0_2; // @[Top.scala 200:12]
  assign n105_I_8_1_0 = n65_O_8_1_0; // @[Top.scala 200:12]
  assign n105_I_8_1_1 = n65_O_8_1_1; // @[Top.scala 200:12]
  assign n105_I_8_1_2 = n65_O_8_1_2; // @[Top.scala 200:12]
  assign n105_I_8_2_0 = n65_O_8_2_0; // @[Top.scala 200:12]
  assign n105_I_8_2_1 = n65_O_8_2_1; // @[Top.scala 200:12]
  assign n105_I_8_2_2 = n65_O_8_2_2; // @[Top.scala 200:12]
  assign n105_I_9_0_0 = n65_O_9_0_0; // @[Top.scala 200:12]
  assign n105_I_9_0_1 = n65_O_9_0_1; // @[Top.scala 200:12]
  assign n105_I_9_0_2 = n65_O_9_0_2; // @[Top.scala 200:12]
  assign n105_I_9_1_0 = n65_O_9_1_0; // @[Top.scala 200:12]
  assign n105_I_9_1_1 = n65_O_9_1_1; // @[Top.scala 200:12]
  assign n105_I_9_1_2 = n65_O_9_1_2; // @[Top.scala 200:12]
  assign n105_I_9_2_0 = n65_O_9_2_0; // @[Top.scala 200:12]
  assign n105_I_9_2_1 = n65_O_9_2_1; // @[Top.scala 200:12]
  assign n105_I_9_2_2 = n65_O_9_2_2; // @[Top.scala 200:12]
  assign n105_I_10_0_0 = n65_O_10_0_0; // @[Top.scala 200:12]
  assign n105_I_10_0_1 = n65_O_10_0_1; // @[Top.scala 200:12]
  assign n105_I_10_0_2 = n65_O_10_0_2; // @[Top.scala 200:12]
  assign n105_I_10_1_0 = n65_O_10_1_0; // @[Top.scala 200:12]
  assign n105_I_10_1_1 = n65_O_10_1_1; // @[Top.scala 200:12]
  assign n105_I_10_1_2 = n65_O_10_1_2; // @[Top.scala 200:12]
  assign n105_I_10_2_0 = n65_O_10_2_0; // @[Top.scala 200:12]
  assign n105_I_10_2_1 = n65_O_10_2_1; // @[Top.scala 200:12]
  assign n105_I_10_2_2 = n65_O_10_2_2; // @[Top.scala 200:12]
  assign n105_I_11_0_0 = n65_O_11_0_0; // @[Top.scala 200:12]
  assign n105_I_11_0_1 = n65_O_11_0_1; // @[Top.scala 200:12]
  assign n105_I_11_0_2 = n65_O_11_0_2; // @[Top.scala 200:12]
  assign n105_I_11_1_0 = n65_O_11_1_0; // @[Top.scala 200:12]
  assign n105_I_11_1_1 = n65_O_11_1_1; // @[Top.scala 200:12]
  assign n105_I_11_1_2 = n65_O_11_1_2; // @[Top.scala 200:12]
  assign n105_I_11_2_0 = n65_O_11_2_0; // @[Top.scala 200:12]
  assign n105_I_11_2_1 = n65_O_11_2_1; // @[Top.scala 200:12]
  assign n105_I_11_2_2 = n65_O_11_2_2; // @[Top.scala 200:12]
  assign n105_I_12_0_0 = n65_O_12_0_0; // @[Top.scala 200:12]
  assign n105_I_12_0_1 = n65_O_12_0_1; // @[Top.scala 200:12]
  assign n105_I_12_0_2 = n65_O_12_0_2; // @[Top.scala 200:12]
  assign n105_I_12_1_0 = n65_O_12_1_0; // @[Top.scala 200:12]
  assign n105_I_12_1_1 = n65_O_12_1_1; // @[Top.scala 200:12]
  assign n105_I_12_1_2 = n65_O_12_1_2; // @[Top.scala 200:12]
  assign n105_I_12_2_0 = n65_O_12_2_0; // @[Top.scala 200:12]
  assign n105_I_12_2_1 = n65_O_12_2_1; // @[Top.scala 200:12]
  assign n105_I_12_2_2 = n65_O_12_2_2; // @[Top.scala 200:12]
  assign n105_I_13_0_0 = n65_O_13_0_0; // @[Top.scala 200:12]
  assign n105_I_13_0_1 = n65_O_13_0_1; // @[Top.scala 200:12]
  assign n105_I_13_0_2 = n65_O_13_0_2; // @[Top.scala 200:12]
  assign n105_I_13_1_0 = n65_O_13_1_0; // @[Top.scala 200:12]
  assign n105_I_13_1_1 = n65_O_13_1_1; // @[Top.scala 200:12]
  assign n105_I_13_1_2 = n65_O_13_1_2; // @[Top.scala 200:12]
  assign n105_I_13_2_0 = n65_O_13_2_0; // @[Top.scala 200:12]
  assign n105_I_13_2_1 = n65_O_13_2_1; // @[Top.scala 200:12]
  assign n105_I_13_2_2 = n65_O_13_2_2; // @[Top.scala 200:12]
  assign n105_I_14_0_0 = n65_O_14_0_0; // @[Top.scala 200:12]
  assign n105_I_14_0_1 = n65_O_14_0_1; // @[Top.scala 200:12]
  assign n105_I_14_0_2 = n65_O_14_0_2; // @[Top.scala 200:12]
  assign n105_I_14_1_0 = n65_O_14_1_0; // @[Top.scala 200:12]
  assign n105_I_14_1_1 = n65_O_14_1_1; // @[Top.scala 200:12]
  assign n105_I_14_1_2 = n65_O_14_1_2; // @[Top.scala 200:12]
  assign n105_I_14_2_0 = n65_O_14_2_0; // @[Top.scala 200:12]
  assign n105_I_14_2_1 = n65_O_14_2_1; // @[Top.scala 200:12]
  assign n105_I_14_2_2 = n65_O_14_2_2; // @[Top.scala 200:12]
  assign n105_I_15_0_0 = n65_O_15_0_0; // @[Top.scala 200:12]
  assign n105_I_15_0_1 = n65_O_15_0_1; // @[Top.scala 200:12]
  assign n105_I_15_0_2 = n65_O_15_0_2; // @[Top.scala 200:12]
  assign n105_I_15_1_0 = n65_O_15_1_0; // @[Top.scala 200:12]
  assign n105_I_15_1_1 = n65_O_15_1_1; // @[Top.scala 200:12]
  assign n105_I_15_1_2 = n65_O_15_1_2; // @[Top.scala 200:12]
  assign n105_I_15_2_0 = n65_O_15_2_0; // @[Top.scala 200:12]
  assign n105_I_15_2_1 = n65_O_15_2_1; // @[Top.scala 200:12]
  assign n105_I_15_2_2 = n65_O_15_2_2; // @[Top.scala 200:12]
  assign n106_valid_up = n105_valid_down; // @[Top.scala 204:19]
  assign n106_I_0_0_0 = n105_O_0_0_0; // @[Top.scala 203:12]
  assign n106_I_1_0_0 = n105_O_1_0_0; // @[Top.scala 203:12]
  assign n106_I_2_0_0 = n105_O_2_0_0; // @[Top.scala 203:12]
  assign n106_I_3_0_0 = n105_O_3_0_0; // @[Top.scala 203:12]
  assign n106_I_4_0_0 = n105_O_4_0_0; // @[Top.scala 203:12]
  assign n106_I_5_0_0 = n105_O_5_0_0; // @[Top.scala 203:12]
  assign n106_I_6_0_0 = n105_O_6_0_0; // @[Top.scala 203:12]
  assign n106_I_7_0_0 = n105_O_7_0_0; // @[Top.scala 203:12]
  assign n106_I_8_0_0 = n105_O_8_0_0; // @[Top.scala 203:12]
  assign n106_I_9_0_0 = n105_O_9_0_0; // @[Top.scala 203:12]
  assign n106_I_10_0_0 = n105_O_10_0_0; // @[Top.scala 203:12]
  assign n106_I_11_0_0 = n105_O_11_0_0; // @[Top.scala 203:12]
  assign n106_I_12_0_0 = n105_O_12_0_0; // @[Top.scala 203:12]
  assign n106_I_13_0_0 = n105_O_13_0_0; // @[Top.scala 203:12]
  assign n106_I_14_0_0 = n105_O_14_0_0; // @[Top.scala 203:12]
  assign n106_I_15_0_0 = n105_O_15_0_0; // @[Top.scala 203:12]
  assign n107_valid_up = n106_valid_down; // @[Top.scala 207:19]
  assign n107_I_0_0 = n106_O_0_0; // @[Top.scala 206:12]
  assign n107_I_1_0 = n106_O_1_0; // @[Top.scala 206:12]
  assign n107_I_2_0 = n106_O_2_0; // @[Top.scala 206:12]
  assign n107_I_3_0 = n106_O_3_0; // @[Top.scala 206:12]
  assign n107_I_4_0 = n106_O_4_0; // @[Top.scala 206:12]
  assign n107_I_5_0 = n106_O_5_0; // @[Top.scala 206:12]
  assign n107_I_6_0 = n106_O_6_0; // @[Top.scala 206:12]
  assign n107_I_7_0 = n106_O_7_0; // @[Top.scala 206:12]
  assign n107_I_8_0 = n106_O_8_0; // @[Top.scala 206:12]
  assign n107_I_9_0 = n106_O_9_0; // @[Top.scala 206:12]
  assign n107_I_10_0 = n106_O_10_0; // @[Top.scala 206:12]
  assign n107_I_11_0 = n106_O_11_0; // @[Top.scala 206:12]
  assign n107_I_12_0 = n106_O_12_0; // @[Top.scala 206:12]
  assign n107_I_13_0 = n106_O_13_0; // @[Top.scala 206:12]
  assign n107_I_14_0 = n106_O_14_0; // @[Top.scala 206:12]
  assign n107_I_15_0 = n106_O_15_0; // @[Top.scala 206:12]
  assign n108_clock = clock;
  assign n108_reset = reset;
  assign n108_valid_up = n1_valid_down; // @[Top.scala 210:19]
  assign n108_I_0 = n1_O_0; // @[Top.scala 209:12]
  assign n108_I_1 = n1_O_1; // @[Top.scala 209:12]
  assign n108_I_2 = n1_O_2; // @[Top.scala 209:12]
  assign n108_I_3 = n1_O_3; // @[Top.scala 209:12]
  assign n108_I_4 = n1_O_4; // @[Top.scala 209:12]
  assign n108_I_5 = n1_O_5; // @[Top.scala 209:12]
  assign n108_I_6 = n1_O_6; // @[Top.scala 209:12]
  assign n108_I_7 = n1_O_7; // @[Top.scala 209:12]
  assign n108_I_8 = n1_O_8; // @[Top.scala 209:12]
  assign n108_I_9 = n1_O_9; // @[Top.scala 209:12]
  assign n108_I_10 = n1_O_10; // @[Top.scala 209:12]
  assign n108_I_11 = n1_O_11; // @[Top.scala 209:12]
  assign n108_I_12 = n1_O_12; // @[Top.scala 209:12]
  assign n108_I_13 = n1_O_13; // @[Top.scala 209:12]
  assign n108_I_14 = n1_O_14; // @[Top.scala 209:12]
  assign n108_I_15 = n1_O_15; // @[Top.scala 209:12]
  assign n109_clock = clock;
  assign n109_reset = reset;
  assign n109_valid_up = n107_valid_down & n108_valid_down; // @[Top.scala 214:19]
  assign n109_I0_0 = n107_O_0; // @[Top.scala 212:13]
  assign n109_I0_1 = n107_O_1; // @[Top.scala 212:13]
  assign n109_I0_2 = n107_O_2; // @[Top.scala 212:13]
  assign n109_I0_3 = n107_O_3; // @[Top.scala 212:13]
  assign n109_I0_4 = n107_O_4; // @[Top.scala 212:13]
  assign n109_I0_5 = n107_O_5; // @[Top.scala 212:13]
  assign n109_I0_6 = n107_O_6; // @[Top.scala 212:13]
  assign n109_I0_7 = n107_O_7; // @[Top.scala 212:13]
  assign n109_I0_8 = n107_O_8; // @[Top.scala 212:13]
  assign n109_I0_9 = n107_O_9; // @[Top.scala 212:13]
  assign n109_I0_10 = n107_O_10; // @[Top.scala 212:13]
  assign n109_I0_11 = n107_O_11; // @[Top.scala 212:13]
  assign n109_I0_12 = n107_O_12; // @[Top.scala 212:13]
  assign n109_I0_13 = n107_O_13; // @[Top.scala 212:13]
  assign n109_I0_14 = n107_O_14; // @[Top.scala 212:13]
  assign n109_I0_15 = n107_O_15; // @[Top.scala 212:13]
  assign n109_I1_0 = n108_O_0; // @[Top.scala 213:13]
  assign n109_I1_1 = n108_O_1; // @[Top.scala 213:13]
  assign n109_I1_2 = n108_O_2; // @[Top.scala 213:13]
  assign n109_I1_3 = n108_O_3; // @[Top.scala 213:13]
  assign n109_I1_4 = n108_O_4; // @[Top.scala 213:13]
  assign n109_I1_5 = n108_O_5; // @[Top.scala 213:13]
  assign n109_I1_6 = n108_O_6; // @[Top.scala 213:13]
  assign n109_I1_7 = n108_O_7; // @[Top.scala 213:13]
  assign n109_I1_8 = n108_O_8; // @[Top.scala 213:13]
  assign n109_I1_9 = n108_O_9; // @[Top.scala 213:13]
  assign n109_I1_10 = n108_O_10; // @[Top.scala 213:13]
  assign n109_I1_11 = n108_O_11; // @[Top.scala 213:13]
  assign n109_I1_12 = n108_O_12; // @[Top.scala 213:13]
  assign n109_I1_13 = n108_O_13; // @[Top.scala 213:13]
  assign n109_I1_14 = n108_O_14; // @[Top.scala 213:13]
  assign n109_I1_15 = n108_O_15; // @[Top.scala 213:13]
  assign n136_clock = clock;
  assign n136_reset = reset;
  assign n136_valid_up = n109_valid_down; // @[Top.scala 217:19]
  assign n136_I_0 = n109_O_0; // @[Top.scala 216:12]
  assign n136_I_1 = n109_O_1; // @[Top.scala 216:12]
  assign n136_I_2 = n109_O_2; // @[Top.scala 216:12]
  assign n136_I_3 = n109_O_3; // @[Top.scala 216:12]
  assign n136_I_4 = n109_O_4; // @[Top.scala 216:12]
  assign n136_I_5 = n109_O_5; // @[Top.scala 216:12]
  assign n136_I_6 = n109_O_6; // @[Top.scala 216:12]
  assign n136_I_7 = n109_O_7; // @[Top.scala 216:12]
  assign n136_I_8 = n109_O_8; // @[Top.scala 216:12]
  assign n136_I_9 = n109_O_9; // @[Top.scala 216:12]
  assign n136_I_10 = n109_O_10; // @[Top.scala 216:12]
  assign n136_I_11 = n109_O_11; // @[Top.scala 216:12]
  assign n136_I_12 = n109_O_12; // @[Top.scala 216:12]
  assign n136_I_13 = n109_O_13; // @[Top.scala 216:12]
  assign n136_I_14 = n109_O_14; // @[Top.scala 216:12]
  assign n136_I_15 = n109_O_15; // @[Top.scala 216:12]
  assign n137_clock = clock;
  assign n137_reset = reset;
  assign n137_valid_up = n136_valid_down; // @[Top.scala 220:19]
  assign n137_I_0 = n136_O_0; // @[Top.scala 219:12]
  assign n137_I_1 = n136_O_1; // @[Top.scala 219:12]
  assign n137_I_2 = n136_O_2; // @[Top.scala 219:12]
  assign n137_I_3 = n136_O_3; // @[Top.scala 219:12]
  assign n137_I_4 = n136_O_4; // @[Top.scala 219:12]
  assign n137_I_5 = n136_O_5; // @[Top.scala 219:12]
  assign n137_I_6 = n136_O_6; // @[Top.scala 219:12]
  assign n137_I_7 = n136_O_7; // @[Top.scala 219:12]
  assign n137_I_8 = n136_O_8; // @[Top.scala 219:12]
  assign n137_I_9 = n136_O_9; // @[Top.scala 219:12]
  assign n137_I_10 = n136_O_10; // @[Top.scala 219:12]
  assign n137_I_11 = n136_O_11; // @[Top.scala 219:12]
  assign n137_I_12 = n136_O_12; // @[Top.scala 219:12]
  assign n137_I_13 = n136_O_13; // @[Top.scala 219:12]
  assign n137_I_14 = n136_O_14; // @[Top.scala 219:12]
  assign n137_I_15 = n136_O_15; // @[Top.scala 219:12]
  assign n138_clock = clock;
  assign n138_reset = reset;
  assign n138_valid_up = n137_valid_down; // @[Top.scala 223:19]
  assign n138_I_0 = n137_O_0; // @[Top.scala 222:12]
  assign n138_I_1 = n137_O_1; // @[Top.scala 222:12]
  assign n138_I_2 = n137_O_2; // @[Top.scala 222:12]
  assign n138_I_3 = n137_O_3; // @[Top.scala 222:12]
  assign n138_I_4 = n137_O_4; // @[Top.scala 222:12]
  assign n138_I_5 = n137_O_5; // @[Top.scala 222:12]
  assign n138_I_6 = n137_O_6; // @[Top.scala 222:12]
  assign n138_I_7 = n137_O_7; // @[Top.scala 222:12]
  assign n138_I_8 = n137_O_8; // @[Top.scala 222:12]
  assign n138_I_9 = n137_O_9; // @[Top.scala 222:12]
  assign n138_I_10 = n137_O_10; // @[Top.scala 222:12]
  assign n138_I_11 = n137_O_11; // @[Top.scala 222:12]
  assign n138_I_12 = n137_O_12; // @[Top.scala 222:12]
  assign n138_I_13 = n137_O_13; // @[Top.scala 222:12]
  assign n138_I_14 = n137_O_14; // @[Top.scala 222:12]
  assign n138_I_15 = n137_O_15; // @[Top.scala 222:12]
endmodule
