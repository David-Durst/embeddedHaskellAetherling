// Latency = 4
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  output [7:0] O
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(clock), // @[:@1296.4]
    .reset('b0), // @[:@1297.4]
    .io_in_x278_TREADY(dontcare), // @[:@1298.4]
    .io_in_x278_TDATA(I_0), // @[:@1298.4]
    .io_in_x278_TID(8'h0),
    .io_in_x278_TDEST(8'h0),
    .io_in_x279_TVALID(valid_down), // @[:@1298.4]
    .io_in_x279_TDATA(O), // @[:@1298.4]
    .io_in_x279_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x286_ctrchain cchain ( // @[:@2879.2]
    .clock(clock), // @[:@2880.4]
    .reset(1'b0), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule

module SRAMVerilogSim
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule

module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 311:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 315:12:@24.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : io_wPort_0_data_0; // @[MemPrimitives.scala 315:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 316:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        ff <= io_wPort_0_data_0;
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh34); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh34); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_parentAck, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  _T_81; // @[Controllers.scala 86:43:@328.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_93; // @[Controllers.scala 92:52:@342.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_134; // @[Controllers.scala 129:57:@382.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  wire  _T_167; // @[package.scala 100:41:@414.4]
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign _T_81 = io_rst | done_0_io_output; // @[Controllers.scala 86:43:@328.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_93 = synchronize | io_rst; // @[Controllers.scala 92:52:@342.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_134 = _T_133 | io_parentAck; // @[Controllers.scala 129:57:@382.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign _T_167 = done_0_io_output & _T_166; // @[package.scala 100:41:@414.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_134 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = _T_81 | io_parentAck; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = _T_93 | io_parentAck; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = _T_167 | io_parentAck; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module SRAM( // @[:@507.2]
  input         clock, // @[:@508.4]
  input  [20:0] io_raddr, // @[:@510.4]
  output [7:0]  io_rdata, // @[:@510.4]
  input         io_backpressure // @[:@510.4]
);
  wire [7:0] SRAMVerilogSim_rdata; // @[SRAM.scala 185:23:@512.4]
  wire [7:0] SRAMVerilogSim_wdata; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_backpressure; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_wen; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_waddrEn; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_raddrEn; // @[SRAM.scala 185:23:@512.4]
  wire [20:0] SRAMVerilogSim_waddr; // @[SRAM.scala 185:23:@512.4]
  wire [20:0] SRAMVerilogSim_raddr; // @[SRAM.scala 185:23:@512.4]
  wire  SRAMVerilogSim_clk; // @[SRAM.scala 185:23:@512.4]
  SRAMVerilogSim #(.DWIDTH(8), .WORDS(2073600), .AWIDTH(21)) SRAMVerilogSim ( // @[SRAM.scala 185:23:@512.4]
    .rdata(SRAMVerilogSim_rdata),
    .wdata(SRAMVerilogSim_wdata),
    .backpressure(SRAMVerilogSim_backpressure),
    .wen(SRAMVerilogSim_wen),
    .waddrEn(SRAMVerilogSim_waddrEn),
    .raddrEn(SRAMVerilogSim_raddrEn),
    .waddr(SRAMVerilogSim_waddr),
    .raddr(SRAMVerilogSim_raddr),
    .clk(SRAMVerilogSim_clk)
  );
  assign io_rdata = SRAMVerilogSim_rdata; // @[SRAM.scala 195:16:@532.4]
  assign SRAMVerilogSim_wdata = 8'h0; // @[SRAM.scala 190:20:@526.4]
  assign SRAMVerilogSim_backpressure = io_backpressure; // @[SRAM.scala 191:27:@527.4]
  assign SRAMVerilogSim_wen = 1'h0; // @[SRAM.scala 188:18:@524.4]
  assign SRAMVerilogSim_waddrEn = 1'h1; // @[SRAM.scala 193:22:@529.4]
  assign SRAMVerilogSim_raddrEn = 1'h1; // @[SRAM.scala 192:22:@528.4]
  assign SRAMVerilogSim_waddr = 21'h0; // @[SRAM.scala 189:20:@525.4]
  assign SRAMVerilogSim_raddr = io_raddr; // @[SRAM.scala 187:20:@523.4]
  assign SRAMVerilogSim_clk = clock; // @[SRAM.scala 186:18:@522.4]
endmodule
module RetimeWrapper_5( // @[:@546.2]
  input         clock, // @[:@547.4]
  input         reset, // @[:@548.4]
  input         io_flow, // @[:@549.4]
  input  [20:0] io_in, // @[:@549.4]
  output [20:0] io_out // @[:@549.4]
);
  wire [20:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire [20:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire [20:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@551.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@551.4]
  RetimeShiftRegister #(.WIDTH(21), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@551.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@564.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@563.4]
  assign sr_init = 21'h0; // @[RetimeShiftRegister.scala 19:16:@562.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@561.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@560.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@558.4]
endmodule
module Mem1D( // @[:@566.2]
  input         clock, // @[:@567.4]
  input         reset, // @[:@568.4]
  input  [20:0] io_r_ofs_0, // @[:@569.4]
  input         io_r_backpressure, // @[:@569.4]
  output [7:0]  io_output // @[:@569.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 705:21:@573.4]
  wire [20:0] SRAM_io_raddr; // @[MemPrimitives.scala 705:21:@573.4]
  wire [7:0] SRAM_io_rdata; // @[MemPrimitives.scala 705:21:@573.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 705:21:@573.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@576.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@576.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@576.4]
  wire [20:0] RetimeWrapper_io_in; // @[package.scala 93:22:@576.4]
  wire [20:0] RetimeWrapper_io_out; // @[package.scala 93:22:@576.4]
  SRAM SRAM ( // @[MemPrimitives.scala 705:21:@573.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@576.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 712:17:@589.4]
  assign SRAM_clock = clock; // @[:@574.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 706:37:@583.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 711:30:@588.4]
  assign RetimeWrapper_clock = clock; // @[:@577.4]
  assign RetimeWrapper_reset = reset; // @[:@578.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@580.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@579.4]
endmodule
module StickySelects( // @[:@591.2]
  input   io_ins_0, // @[:@594.4]
  output  io_outs_0 // @[:@594.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 34:26:@596.4]
endmodule
module RetimeWrapper_6( // @[:@610.2]
  input   clock, // @[:@611.4]
  input   reset, // @[:@612.4]
  input   io_flow, // @[:@613.4]
  input   io_in, // @[:@613.4]
  output  io_out // @[:@613.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@615.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@615.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@615.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@628.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@627.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@626.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@625.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@624.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@622.4]
endmodule
module x280_outbuf_0( // @[:@630.2]
  input         clock, // @[:@631.4]
  input         reset, // @[:@632.4]
  input  [20:0] io_rPort_0_ofs_0, // @[:@633.4]
  input         io_rPort_0_en_0, // @[:@633.4]
  input         io_rPort_0_backpressure, // @[:@633.4]
  output [7:0]  io_rPort_0_output_0 // @[:@633.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@648.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@648.4]
  wire [20:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@648.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@648.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@648.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@674.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@674.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@688.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@688.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@688.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@688.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@688.4]
  wire  _T_76; // @[MemPrimitives.scala 123:41:@678.4]
  wire [22:0] _T_78; // @[Cat.scala 30:58:@680.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@648.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 121:29:@674.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@688.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@678.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@680.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 148:13:@695.4]
  assign Mem1D_clock = clock; // @[:@649.4]
  assign Mem1D_reset = reset; // @[:@650.4]
  assign Mem1D_io_r_ofs_0 = _T_78[20:0]; // @[MemPrimitives.scala 127:28:@684.4]
  assign Mem1D_io_r_backpressure = _T_78[21]; // @[MemPrimitives.scala 128:32:@685.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 122:60:@677.4]
  assign RetimeWrapper_clock = clock; // @[:@689.4]
  assign RetimeWrapper_reset = reset; // @[:@690.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@692.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@691.4]
endmodule
module x556_sm( // @[:@839.2]
  input   clock, // @[:@840.4]
  input   reset, // @[:@841.4]
  input   io_enable, // @[:@842.4]
  output  io_done, // @[:@842.4]
  input   io_ctrDone, // @[:@842.4]
  output  io_ctrInc, // @[:@842.4]
  input   io_parentAck, // @[:@842.4]
  input   io_doneIn_0, // @[:@842.4]
  input   io_doneIn_1, // @[:@842.4]
  output  io_enableOut_0, // @[:@842.4]
  output  io_enableOut_1, // @[:@842.4]
  output  io_childAck_0, // @[:@842.4]
  output  io_childAck_1 // @[:@842.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@845.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@845.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@848.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@848.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@851.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@851.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@854.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@854.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@883.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@886.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@886.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@987.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1004.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1004.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1004.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1004.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1004.4]
  wire  allDone; // @[Controllers.scala 80:47:@857.4]
  wire  synchronize; // @[Controllers.scala 146:56:@911.4]
  wire  _T_127; // @[Controllers.scala 150:35:@913.4]
  wire  _T_129; // @[Controllers.scala 150:60:@914.4]
  wire  _T_130; // @[Controllers.scala 150:58:@915.4]
  wire  _T_132; // @[Controllers.scala 150:76:@916.4]
  wire  _T_133; // @[Controllers.scala 150:74:@917.4]
  wire  _T_135; // @[Controllers.scala 150:97:@918.4]
  wire  _T_136; // @[Controllers.scala 150:95:@919.4]
  wire  _T_152; // @[Controllers.scala 150:35:@937.4]
  wire  _T_154; // @[Controllers.scala 150:60:@938.4]
  wire  _T_155; // @[Controllers.scala 150:58:@939.4]
  wire  _T_157; // @[Controllers.scala 150:76:@940.4]
  wire  _T_158; // @[Controllers.scala 150:74:@941.4]
  wire  _T_161; // @[Controllers.scala 150:95:@943.4]
  wire  _T_179; // @[Controllers.scala 213:68:@965.4]
  wire  _T_181; // @[Controllers.scala 213:90:@967.4]
  wire  _T_183; // @[Controllers.scala 213:132:@969.4]
  wire  _T_184; // @[Controllers.scala 213:130:@970.4]
  wire  _T_185; // @[Controllers.scala 213:156:@971.4]
  wire  _T_187; // @[Controllers.scala 213:68:@974.4]
  wire  _T_189; // @[Controllers.scala 213:90:@976.4]
  wire  _T_196; // @[package.scala 100:49:@982.4]
  reg  _T_199; // @[package.scala 48:56:@983.4]
  reg [31:0] _RAND_0;
  wire  _T_200; // @[package.scala 100:41:@985.4]
  reg  _T_213; // @[package.scala 48:56:@1001.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@845.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@848.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@851.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@854.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@883.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@886.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@987.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1004.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@857.4]
  assign synchronize = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 146:56:@911.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 150:35:@913.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 150:60:@914.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 150:58:@915.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 150:76:@916.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 150:74:@917.4]
  assign _T_135 = io_ctrDone == 1'h0; // @[Controllers.scala 150:97:@918.4]
  assign _T_136 = _T_133 & _T_135; // @[Controllers.scala 150:95:@919.4]
  assign _T_152 = ~ iterDone_1_io_output; // @[Controllers.scala 150:35:@937.4]
  assign _T_154 = io_doneIn_1 == 1'h0; // @[Controllers.scala 150:60:@938.4]
  assign _T_155 = _T_152 & _T_154; // @[Controllers.scala 150:58:@939.4]
  assign _T_157 = done_1_io_output == 1'h0; // @[Controllers.scala 150:76:@940.4]
  assign _T_158 = _T_155 & _T_157; // @[Controllers.scala 150:74:@941.4]
  assign _T_161 = _T_158 & _T_135; // @[Controllers.scala 150:95:@943.4]
  assign _T_179 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@965.4]
  assign _T_181 = _T_179 & _T_127; // @[Controllers.scala 213:90:@967.4]
  assign _T_183 = ~ allDone; // @[Controllers.scala 213:132:@969.4]
  assign _T_184 = _T_181 & _T_183; // @[Controllers.scala 213:130:@970.4]
  assign _T_185 = ~ io_ctrDone; // @[Controllers.scala 213:156:@971.4]
  assign _T_187 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@974.4]
  assign _T_189 = _T_187 & _T_152; // @[Controllers.scala 213:90:@976.4]
  assign _T_196 = allDone == 1'h0; // @[package.scala 100:49:@982.4]
  assign _T_200 = allDone & _T_199; // @[package.scala 100:41:@985.4]
  assign io_done = RetimeWrapper_1_io_out; // @[Controllers.scala 245:13:@1011.4]
  assign io_ctrInc = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 143:17:@910.4]
  assign io_enableOut_0 = _T_184 & _T_185; // @[Controllers.scala 213:55:@973.4]
  assign io_enableOut_1 = _T_189 & _T_183; // @[Controllers.scala 213:55:@981.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@962.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@964.4]
  assign active_0_clock = clock; // @[:@846.4]
  assign active_0_reset = reset; // @[:@847.4]
  assign active_0_io_input_set = _T_136 & io_enable; // @[Controllers.scala 150:32:@922.4]
  assign active_0_io_input_reset = io_doneIn_0 | io_parentAck; // @[Controllers.scala 151:34:@926.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@860.4]
  assign active_1_clock = clock; // @[:@849.4]
  assign active_1_reset = reset; // @[:@850.4]
  assign active_1_io_input_set = _T_161 & io_enable; // @[Controllers.scala 150:32:@946.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_parentAck; // @[Controllers.scala 151:34:@950.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@861.4]
  assign done_0_clock = clock; // @[:@852.4]
  assign done_0_reset = reset; // @[:@853.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@936.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@872.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@862.4]
  assign done_1_clock = clock; // @[:@855.4]
  assign done_1_reset = reset; // @[:@856.4]
  assign done_1_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@960.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@881.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@863.4]
  assign iterDone_0_clock = clock; // @[:@884.4]
  assign iterDone_0_reset = reset; // @[:@885.4]
  assign iterDone_0_io_input_set = io_doneIn_0; // @[Controllers.scala 152:34:@932.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@899.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@889.4]
  assign iterDone_1_clock = clock; // @[:@887.4]
  assign iterDone_1_reset = reset; // @[:@888.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 152:34:@956.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@908.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@890.4]
  assign RetimeWrapper_clock = clock; // @[:@988.4]
  assign RetimeWrapper_reset = reset; // @[:@989.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@991.4]
  assign RetimeWrapper_io_in = _T_200 | io_parentAck; // @[package.scala 94:16:@990.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1005.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1006.4]
  assign RetimeWrapper_1_io_flow = io_enable; // @[package.scala 95:18:@1008.4]
  assign RetimeWrapper_1_io_in = allDone & _T_213; // @[package.scala 94:16:@1007.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_199 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_213 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_199 <= 1'h0;
    end else begin
      _T_199 <= _T_196;
    end
    if (reset) begin
      _T_213 <= 1'h0;
    end else begin
      _T_213 <= _T_196;
    end
  end
endmodule
module x418_outr_UnitPipe_sm( // @[:@1428.2]
  input   clock, // @[:@1429.4]
  input   reset, // @[:@1430.4]
  input   io_enable, // @[:@1431.4]
  output  io_done, // @[:@1431.4]
  input   io_parentAck, // @[:@1431.4]
  input   io_doneIn_0, // @[:@1431.4]
  input   io_doneIn_1, // @[:@1431.4]
  output  io_enableOut_0, // @[:@1431.4]
  output  io_enableOut_1, // @[:@1431.4]
  output  io_childAck_0, // @[:@1431.4]
  output  io_childAck_1, // @[:@1431.4]
  input   io_ctrCopyDone_0, // @[:@1431.4]
  input   io_ctrCopyDone_1 // @[:@1431.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@1434.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@1434.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@1437.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@1437.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@1440.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@1440.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1443.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1443.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1472.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1475.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1475.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1516.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1530.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1548.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1585.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1599.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1617.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1664.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1681.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1681.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1681.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1681.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1681.4]
  wire  allDone; // @[Controllers.scala 80:47:@1446.4]
  wire  _T_127; // @[Controllers.scala 165:35:@1500.4]
  wire  _T_129; // @[Controllers.scala 165:60:@1501.4]
  wire  _T_130; // @[Controllers.scala 165:58:@1502.4]
  wire  _T_132; // @[Controllers.scala 165:76:@1503.4]
  wire  _T_133; // @[Controllers.scala 165:74:@1504.4]
  wire  _T_137; // @[Controllers.scala 165:109:@1507.4]
  wire  _T_140; // @[Controllers.scala 165:141:@1509.4]
  wire  _T_148; // @[package.scala 96:25:@1521.4 package.scala 96:25:@1522.4]
  wire  _T_152; // @[Controllers.scala 167:54:@1524.4]
  wire  _T_153; // @[Controllers.scala 167:52:@1525.4]
  wire  _T_160; // @[package.scala 96:25:@1535.4 package.scala 96:25:@1536.4]
  wire  _T_178; // @[package.scala 96:25:@1553.4 package.scala 96:25:@1554.4]
  wire  _T_182; // @[Controllers.scala 169:67:@1556.4]
  wire  _T_183; // @[Controllers.scala 169:86:@1557.4]
  wire  _T_195; // @[Controllers.scala 165:35:@1569.4]
  wire  _T_197; // @[Controllers.scala 165:60:@1570.4]
  wire  _T_198; // @[Controllers.scala 165:58:@1571.4]
  wire  _T_200; // @[Controllers.scala 165:76:@1572.4]
  wire  _T_201; // @[Controllers.scala 165:74:@1573.4]
  wire  _T_205; // @[Controllers.scala 165:109:@1576.4]
  wire  _T_208; // @[Controllers.scala 165:141:@1578.4]
  wire  _T_216; // @[package.scala 96:25:@1590.4 package.scala 96:25:@1591.4]
  wire  _T_220; // @[Controllers.scala 167:54:@1593.4]
  wire  _T_221; // @[Controllers.scala 167:52:@1594.4]
  wire  _T_228; // @[package.scala 96:25:@1604.4 package.scala 96:25:@1605.4]
  wire  _T_246; // @[package.scala 96:25:@1622.4 package.scala 96:25:@1623.4]
  wire  _T_250; // @[Controllers.scala 169:67:@1625.4]
  wire  _T_251; // @[Controllers.scala 169:86:@1626.4]
  wire  _T_265; // @[Controllers.scala 213:68:@1642.4]
  wire  _T_267; // @[Controllers.scala 213:90:@1644.4]
  wire  _T_269; // @[Controllers.scala 213:132:@1646.4]
  wire  _T_273; // @[Controllers.scala 213:68:@1651.4]
  wire  _T_275; // @[Controllers.scala 213:90:@1653.4]
  wire  _T_282; // @[package.scala 100:49:@1659.4]
  reg  _T_285; // @[package.scala 48:56:@1660.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@1662.4]
  reg  _T_299; // @[package.scala 48:56:@1678.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@1434.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@1437.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@1440.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1443.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1472.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1475.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1516.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1530.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1548.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1585.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1599.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1617.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1664.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1681.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1446.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1500.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1501.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@1502.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1503.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@1504.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@1507.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1509.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@1521.4 package.scala 96:25:@1522.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@1524.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@1525.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1535.4 package.scala 96:25:@1536.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1553.4 package.scala 96:25:@1554.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@1556.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@1557.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1569.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1570.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@1571.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1572.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@1573.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@1576.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1578.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1590.4 package.scala 96:25:@1591.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@1593.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@1594.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1604.4 package.scala 96:25:@1605.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1622.4 package.scala 96:25:@1623.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@1625.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@1626.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1642.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@1644.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@1646.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1651.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@1653.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@1659.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@1662.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@1688.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@1650.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@1658.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1639.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1641.4]
  assign active_0_clock = clock; // @[:@1435.4]
  assign active_0_reset = reset; // @[:@1436.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@1511.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1515.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1449.4]
  assign active_1_clock = clock; // @[:@1438.4]
  assign active_1_reset = reset; // @[:@1439.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@1580.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1584.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1450.4]
  assign done_0_clock = clock; // @[:@1441.4]
  assign done_0_reset = reset; // @[:@1442.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@1561.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1461.4 Controllers.scala 170:32:@1568.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1451.4]
  assign done_1_clock = clock; // @[:@1444.4]
  assign done_1_reset = reset; // @[:@1445.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@1630.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1470.4 Controllers.scala 170:32:@1637.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1452.4]
  assign iterDone_0_clock = clock; // @[:@1473.4]
  assign iterDone_0_reset = reset; // @[:@1474.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@1529.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@1488.4 Controllers.scala 168:36:@1545.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1478.4]
  assign iterDone_1_clock = clock; // @[:@1476.4]
  assign iterDone_1_reset = reset; // @[:@1477.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@1598.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@1497.4 Controllers.scala 168:36:@1614.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1479.4]
  assign RetimeWrapper_clock = clock; // @[:@1517.4]
  assign RetimeWrapper_reset = reset; // @[:@1518.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1520.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1519.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1531.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1532.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1534.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1533.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1549.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1550.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1552.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1551.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1586.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1587.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1589.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1588.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1600.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1601.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1603.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1602.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1618.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1619.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1621.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1620.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1665.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1666.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1668.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@1667.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1682.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1683.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@1685.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@1684.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module CompactingIncDincCtr( // @[:@1917.2]
  input   clock, // @[:@1918.4]
  input   reset, // @[:@1919.4]
  input   io_input_inc_en_0, // @[:@1920.4]
  input   io_input_dinc_en_0, // @[:@1920.4]
  output  io_output_full // @[:@1920.4]
);
  reg [31:0] cnt; // @[Counter.scala 170:20:@1922.4]
  reg [31:0] _RAND_0;
  wire [14:0] numPushed; // @[Counter.scala 172:47:@1923.4]
  wire [14:0] numPopped; // @[Counter.scala 173:48:@1924.4]
  wire [31:0] _GEN_0; // @[Counter.scala 174:14:@1925.4]
  wire [32:0] _T_37; // @[Counter.scala 174:14:@1925.4]
  wire [31:0] _T_38; // @[Counter.scala 174:14:@1926.4]
  wire [31:0] _T_39; // @[Counter.scala 174:14:@1927.4]
  wire [31:0] _GEN_1; // @[Counter.scala 174:26:@1928.4]
  wire [32:0] _T_40; // @[Counter.scala 174:26:@1928.4]
  wire [31:0] _T_41; // @[Counter.scala 174:26:@1929.4]
  wire [31:0] _T_42; // @[Counter.scala 174:26:@1930.4]
  assign numPushed = io_input_inc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 172:47:@1923.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 173:48:@1924.4]
  assign _GEN_0 = {{17{numPushed[14]}},numPushed}; // @[Counter.scala 174:14:@1925.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1925.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1926.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 174:14:@1927.4]
  assign _GEN_1 = {{17{numPopped[14]}},numPopped}; // @[Counter.scala 174:26:@1928.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1928.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1929.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 174:26:@1930.4]
  assign io_output_full = $signed(cnt) > $signed(32'sh1dff); // @[Counter.scala 180:18:@1944.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module x281_fifoinraw_0( // @[:@2067.2]
  input   clock, // @[:@2068.4]
  input   reset // @[:@2069.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 382:24:@2114.4]
  wire  elements_reset; // @[MemPrimitives.scala 382:24:@2114.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 382:24:@2114.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 382:24:@2114.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 382:24:@2114.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 382:24:@2114.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign elements_clock = clock; // @[:@2115.4]
  assign elements_reset = reset; // @[:@2116.4]
  assign elements_io_input_inc_en_0 = 1'h0; // @[MemPrimitives.scala 384:79:@2126.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 385:80:@2127.4]
endmodule
module x282_fifoinpacked_0( // @[:@2490.2]
  input   clock, // @[:@2491.4]
  input   reset, // @[:@2492.4]
  input   io_wPort_0_en_0, // @[:@2493.4]
  output  io_full, // @[:@2493.4]
  input   io_active_0_in, // @[:@2493.4]
  output  io_active_0_out // @[:@2493.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 382:24:@2537.4]
  wire  elements_reset; // @[MemPrimitives.scala 382:24:@2537.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 382:24:@2537.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 382:24:@2537.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 382:24:@2537.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 382:24:@2537.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 429:39:@2611.4]
  assign io_active_0_out = io_active_0_in; // @[MemPrimitives.scala 427:129:@2609.4]
  assign elements_clock = clock; // @[:@2538.4]
  assign elements_reset = reset; // @[:@2539.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 384:79:@2549.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 385:80:@2550.4]
endmodule
module FF_7( // @[:@3040.2]
  input         clock, // @[:@3041.4]
  input         reset, // @[:@3042.4]
  output [12:0] io_rPort_0_output_0, // @[:@3043.4]
  input  [12:0] io_wPort_0_data_0, // @[:@3043.4]
  input         io_wPort_0_reset, // @[:@3043.4]
  input         io_wPort_0_en_0 // @[:@3043.4]
);
  reg [12:0] ff; // @[MemPrimitives.scala 311:19:@3058.4]
  reg [31:0] _RAND_0;
  wire [12:0] _T_68; // @[MemPrimitives.scala 315:32:@3060.4]
  wire [12:0] _T_69; // @[MemPrimitives.scala 315:12:@3061.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 315:32:@3060.4]
  assign _T_69 = io_wPort_0_reset ? 13'h0 : _T_68; // @[MemPrimitives.scala 315:12:@3061.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 316:34:@3063.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 13'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 13'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_1( // @[:@3078.2]
  input         clock, // @[:@3079.4]
  input         reset, // @[:@3080.4]
  input         io_setup_saturate, // @[:@3081.4]
  input         io_input_reset, // @[:@3081.4]
  input         io_input_enable, // @[:@3081.4]
  output [12:0] io_output_count_0, // @[:@3081.4]
  output        io_output_oobs_0, // @[:@3081.4]
  output        io_output_done, // @[:@3081.4]
  output        io_output_saturated // @[:@3081.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3094.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3094.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3094.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3094.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3094.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3094.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3110.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3110.4]
  wire  _T_36; // @[Counter.scala 264:45:@3113.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3138.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3139.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3140.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3141.4]
  wire  _T_57; // @[Counter.scala 293:18:@3143.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3151.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3153.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3154.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3155.4]
  wire  _T_75; // @[Counter.scala 322:102:@3159.4]
  wire  _T_77; // @[Counter.scala 322:130:@3160.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3094.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3110.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3113.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3138.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3139.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3140.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3141.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh438); // @[Counter.scala 293:18:@3143.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3151.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3153.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3154.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3155.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3159.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh438); // @[Counter.scala 322:130:@3160.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3158.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3162.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3164.4]
  assign io_output_saturated = io_setup_saturate & _T_57; // @[Counter.scala 340:25:@3167.4]
  assign bases_0_clock = clock; // @[:@3095.4]
  assign bases_0_reset = reset; // @[:@3096.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3157.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3136.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3137.4]
  assign SRFF_clock = clock; // @[:@3111.4]
  assign SRFF_reset = reset; // @[:@3112.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3115.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3117.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3118.4]
endmodule
module SingleCounter_2( // @[:@3207.2]
  input         clock, // @[:@3208.4]
  input         reset, // @[:@3209.4]
  input         io_setup_saturate, // @[:@3210.4]
  input         io_input_reset, // @[:@3210.4]
  input         io_input_enable, // @[:@3210.4]
  output [12:0] io_output_count_0, // @[:@3210.4]
  output        io_output_oobs_0, // @[:@3210.4]
  output        io_output_done // @[:@3210.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3223.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3223.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3223.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3223.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3223.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3223.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3239.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3239.4]
  wire  _T_36; // @[Counter.scala 264:45:@3242.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3267.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3268.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3269.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3270.4]
  wire  _T_57; // @[Counter.scala 293:18:@3272.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3280.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3282.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3283.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3284.4]
  wire  _T_75; // @[Counter.scala 322:102:@3288.4]
  wire  _T_77; // @[Counter.scala 322:130:@3289.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3223.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3239.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3242.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3267.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3268.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3269.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3270.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh780); // @[Counter.scala 293:18:@3272.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3280.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3282.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3283.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3284.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3288.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh780); // @[Counter.scala 322:130:@3289.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3287.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3291.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3293.4]
  assign bases_0_clock = clock; // @[:@3224.4]
  assign bases_0_reset = reset; // @[:@3225.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3286.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3265.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3266.4]
  assign SRFF_clock = clock; // @[:@3240.4]
  assign SRFF_reset = reset; // @[:@3241.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3244.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3246.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3247.4]
endmodule
module x286_ctrchain( // @[:@3298.2]
  input         clock, // @[:@3299.4]
  input         reset, // @[:@3300.4]
  input         io_input_reset, // @[:@3301.4]
  input         io_input_enable, // @[:@3301.4]
  output [12:0] io_output_counts_1, // @[:@3301.4]
  output [12:0] io_output_counts_0, // @[:@3301.4]
  output        io_output_oobs_0, // @[:@3301.4]
  output        io_output_oobs_1, // @[:@3301.4]
  output        io_output_done // @[:@3301.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@3303.4]
  wire [12:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@3303.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@3306.4]
  wire [12:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@3306.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@3306.4]
  wire  isDone; // @[Counter.scala 541:51:@3323.4]
  reg  wasDone; // @[Counter.scala 542:24:@3324.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@3332.4]
  wire  _T_66; // @[Counter.scala 546:80:@3333.4]
  reg  doneLatch; // @[Counter.scala 550:26:@3338.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@3339.4]
  wire  _T_74; // @[Counter.scala 551:19:@3340.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@3303.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@3306.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@3323.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@3332.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@3333.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@3339.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@3340.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@3345.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@3342.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3344.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3347.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@3335.4]
  assign ctrs_0_clock = clock; // @[:@3304.4]
  assign ctrs_0_reset = reset; // @[:@3305.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 530:29:@3320.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3312.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@3319.4]
  assign ctrs_1_clock = clock; // @[:@3307.4]
  assign ctrs_1_reset = reset; // @[:@3308.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@3322.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3316.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@3317.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_21( // @[:@3387.2]
  input   clock, // @[:@3388.4]
  input   reset, // @[:@3389.4]
  input   io_flow, // @[:@3390.4]
  input   io_in, // @[:@3390.4]
  output  io_out // @[:@3390.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3392.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@3392.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3405.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3404.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3403.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3402.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3401.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3399.4]
endmodule
module RetimeWrapper_25( // @[:@3515.2]
  input   clock, // @[:@3516.4]
  input   reset, // @[:@3517.4]
  input   io_flow, // @[:@3518.4]
  input   io_in, // @[:@3518.4]
  output  io_out // @[:@3518.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3520.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@3520.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3533.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3532.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3531.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3530.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3529.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3527.4]
endmodule
module x300_inr_Foreach_sm( // @[:@3535.2]
  input   clock, // @[:@3536.4]
  input   reset, // @[:@3537.4]
  input   io_enable, // @[:@3538.4]
  output  io_done, // @[:@3538.4]
  output  io_doneLatch, // @[:@3538.4]
  input   io_ctrDone, // @[:@3538.4]
  output  io_datapathEn, // @[:@3538.4]
  output  io_ctrInc, // @[:@3538.4]
  output  io_ctrRst, // @[:@3538.4]
  input   io_parentAck, // @[:@3538.4]
  input   io_backpressure, // @[:@3538.4]
  input   io_break // @[:@3538.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3540.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3540.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3540.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3540.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3540.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3540.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3543.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3543.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3543.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3543.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3543.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3543.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3577.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3599.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3611.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3619.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3635.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3635.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3635.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3635.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3635.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3548.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3549.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3550.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3551.4]
  wire  _T_100; // @[package.scala 100:49:@3568.4]
  reg  _T_103; // @[package.scala 48:56:@3569.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3582.4 package.scala 96:25:@3583.4]
  wire  _T_110; // @[package.scala 100:49:@3584.4]
  reg  _T_113; // @[package.scala 48:56:@3585.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3587.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3592.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3593.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3596.4]
  wire  _T_124; // @[package.scala 96:25:@3604.4 package.scala 96:25:@3605.4]
  wire  _T_126; // @[package.scala 100:49:@3606.4]
  reg  _T_129; // @[package.scala 48:56:@3607.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3629.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3631.4]
  reg  _T_153; // @[package.scala 48:56:@3632.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3640.4 package.scala 96:25:@3641.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3642.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3643.4]
  SRFF active ( // @[Controllers.scala 261:22:@3540.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3543.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@3577.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3599.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3611.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3619.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@3635.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3548.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3549.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3550.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3551.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3568.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3582.4 package.scala 96:25:@3583.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3584.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3587.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3592.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3593.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3596.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3604.4 package.scala 96:25:@3605.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3606.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3631.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3640.4 package.scala 96:25:@3641.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3642.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3643.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3610.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3645.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3595.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3598.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3590.4]
  assign active_clock = clock; // @[:@3541.4]
  assign active_reset = reset; // @[:@3542.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3553.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3557.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3558.4]
  assign done_clock = clock; // @[:@3544.4]
  assign done_reset = reset; // @[:@3545.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3573.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3566.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3567.4]
  assign RetimeWrapper_clock = clock; // @[:@3578.4]
  assign RetimeWrapper_reset = reset; // @[:@3579.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3581.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3580.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3600.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3601.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3603.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3602.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3612.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3613.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3615.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3614.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3620.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3621.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3623.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3622.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3636.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3637.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3639.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3638.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module SimBlackBoxesfix2fixBox( // @[:@3752.2]
  input  [31:0] io_a, // @[:@3755.4]
  output [31:0] io_b // @[:@3755.4]
);
  assign io_b = io_a; // @[SimBlackBoxes.scala 99:40:@3768.4]
endmodule
module _( // @[:@3770.2]
  input  [31:0] io_b, // @[:@3773.4]
  output [31:0] io_result // @[:@3773.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3778.4]
  wire [31:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3778.4]
  SimBlackBoxesfix2fixBox SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3778.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3791.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3786.4]
endmodule
module SimBlackBoxesfix2fixBox_2( // @[:@3834.2]
  input  [31:0] io_a, // @[:@3837.4]
  output [32:0] io_b // @[:@3837.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@3847.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@3847.4]
  assign io_b = {_T_20,io_a}; // @[SimBlackBoxes.scala 99:40:@3852.4]
endmodule
module __2( // @[:@3854.2]
  input  [31:0] io_b, // @[:@3857.4]
  output [32:0] io_result // @[:@3857.4]
);
  wire [31:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@3862.4]
  wire [32:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@3862.4]
  SimBlackBoxesfix2fixBox_2 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@3862.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@3875.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@3870.4]
endmodule
module RetimeWrapper_29( // @[:@3932.2]
  input         clock, // @[:@3933.4]
  input         reset, // @[:@3934.4]
  input         io_flow, // @[:@3935.4]
  input  [31:0] io_in, // @[:@3935.4]
  output [31:0] io_out // @[:@3935.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3937.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3937.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3950.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3949.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3948.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3947.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3946.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3944.4]
endmodule
module fix2fixBox( // @[:@3952.2]
  input         clock, // @[:@3953.4]
  input         reset, // @[:@3954.4]
  input  [32:0] io_a, // @[:@3955.4]
  input         io_flow, // @[:@3955.4]
  output [31:0] io_b // @[:@3955.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3968.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3968.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3968.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3968.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3968.4]
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@3968.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@3975.4]
  assign RetimeWrapper_clock = clock; // @[:@3969.4]
  assign RetimeWrapper_reset = reset; // @[:@3970.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@3972.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@3971.4]
endmodule
module x467_sub( // @[:@3977.2]
  input         clock, // @[:@3978.4]
  input         reset, // @[:@3979.4]
  input  [31:0] io_a, // @[:@3980.4]
  input  [31:0] io_b, // @[:@3980.4]
  input         io_flow, // @[:@3980.4]
  output [31:0] io_result // @[:@3980.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@3988.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@3988.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@3995.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@3995.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@4014.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@4014.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@4014.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@4014.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@4014.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@3993.4 Math.scala 713:14:@3994.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@4000.4 Math.scala 713:14:@4001.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@4002.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@4003.4]
  __2 _ ( // @[Math.scala 709:24:@3988.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@3995.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 182:30:@4014.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@3993.4 Math.scala 713:14:@3994.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@4000.4 Math.scala 713:14:@4001.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@4002.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@4003.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@4022.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@3991.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@3998.4]
  assign fix2fixBox_clock = clock; // @[:@4015.4]
  assign fix2fixBox_reset = reset; // @[:@4016.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@4017.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@4020.4]
endmodule
module x292_sum( // @[:@4199.2]
  input         clock, // @[:@4200.4]
  input         reset, // @[:@4201.4]
  input  [31:0] io_a, // @[:@4202.4]
  input  [31:0] io_b, // @[:@4202.4]
  input         io_flow, // @[:@4202.4]
  output [31:0] io_result // @[:@4202.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@4210.4]
  wire [32:0] __io_result; // @[Math.scala 709:24:@4210.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@4217.4]
  wire [32:0] __1_io_result; // @[Math.scala 709:24:@4217.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4235.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4235.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4235.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4235.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4235.4]
  wire [32:0] a_upcast_number; // @[Math.scala 712:22:@4215.4 Math.scala 713:14:@4216.4]
  wire [32:0] b_upcast_number; // @[Math.scala 712:22:@4222.4 Math.scala 713:14:@4223.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@4224.4]
  __2 _ ( // @[Math.scala 709:24:@4210.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 709:24:@4217.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 141:30:@4235.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@4215.4 Math.scala 713:14:@4216.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@4222.4 Math.scala 713:14:@4223.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4224.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4243.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@4213.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@4220.4]
  assign fix2fixBox_clock = clock; // @[:@4236.4]
  assign fix2fixBox_reset = reset; // @[:@4237.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4238.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4241.4]
endmodule
module x300_inr_Foreach_kernelx300_inr_Foreach_concrete1( // @[:@4760.2]
  input         clock, // @[:@4761.4]
  input         reset, // @[:@4762.4]
  output        io_in_x282_fifoinpacked_0_wPort_0_en_0, // @[:@4763.4]
  input         io_in_x282_fifoinpacked_0_full, // @[:@4763.4]
  output        io_in_x282_fifoinpacked_0_active_0_in, // @[:@4763.4]
  input         io_in_x282_fifoinpacked_0_active_0_out, // @[:@4763.4]
  input         io_sigsIn_backpressure, // @[:@4763.4]
  input         io_sigsIn_datapathEn, // @[:@4763.4]
  input         io_sigsIn_break, // @[:@4763.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_1, // @[:@4763.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@4763.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@4763.4]
  input         io_sigsIn_cchainOutputs_0_oobs_1, // @[:@4763.4]
  input         io_rr // @[:@4763.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@4797.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@4797.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@4809.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@4809.4]
  wire  x467_sub_1_clock; // @[Math.scala 191:24:@4836.4]
  wire  x467_sub_1_reset; // @[Math.scala 191:24:@4836.4]
  wire [31:0] x467_sub_1_io_a; // @[Math.scala 191:24:@4836.4]
  wire [31:0] x467_sub_1_io_b; // @[Math.scala 191:24:@4836.4]
  wire  x467_sub_1_io_flow; // @[Math.scala 191:24:@4836.4]
  wire [31:0] x467_sub_1_io_result; // @[Math.scala 191:24:@4836.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4846.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4846.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@4846.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@4846.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@4846.4]
  wire  x292_sum_1_clock; // @[Math.scala 150:24:@4855.4]
  wire  x292_sum_1_reset; // @[Math.scala 150:24:@4855.4]
  wire [31:0] x292_sum_1_io_a; // @[Math.scala 150:24:@4855.4]
  wire [31:0] x292_sum_1_io_b; // @[Math.scala 150:24:@4855.4]
  wire  x292_sum_1_io_flow; // @[Math.scala 150:24:@4855.4]
  wire [31:0] x292_sum_1_io_result; // @[Math.scala 150:24:@4855.4]
  wire  x293_sum_1_clock; // @[Math.scala 150:24:@4867.4]
  wire  x293_sum_1_reset; // @[Math.scala 150:24:@4867.4]
  wire [31:0] x293_sum_1_io_a; // @[Math.scala 150:24:@4867.4]
  wire [31:0] x293_sum_1_io_b; // @[Math.scala 150:24:@4867.4]
  wire  x293_sum_1_io_flow; // @[Math.scala 150:24:@4867.4]
  wire [31:0] x293_sum_1_io_result; // @[Math.scala 150:24:@4867.4]
  wire  x469_sum_1_clock; // @[Math.scala 150:24:@4882.4]
  wire  x469_sum_1_reset; // @[Math.scala 150:24:@4882.4]
  wire [31:0] x469_sum_1_io_a; // @[Math.scala 150:24:@4882.4]
  wire [31:0] x469_sum_1_io_b; // @[Math.scala 150:24:@4882.4]
  wire  x469_sum_1_io_flow; // @[Math.scala 150:24:@4882.4]
  wire [31:0] x469_sum_1_io_result; // @[Math.scala 150:24:@4882.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@4916.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@4916.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@4916.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@4916.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@4916.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@4925.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@4925.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@4925.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@4925.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@4925.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@4936.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@4936.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@4936.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@4936.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@4936.4]
  wire  _T_327; // @[sm_x300_inr_Foreach.scala 62:18:@4822.4]
  wire  _T_328; // @[sm_x300_inr_Foreach.scala 62:55:@4823.4]
  wire [31:0] b287_number; // @[Math.scala 712:22:@4802.4 Math.scala 713:14:@4803.4]
  wire [42:0] _GEN_0; // @[Math.scala 450:32:@4827.4]
  wire [42:0] _T_332; // @[Math.scala 450:32:@4827.4]
  wire [38:0] _GEN_1; // @[Math.scala 450:32:@4832.4]
  wire [38:0] _T_336; // @[Math.scala 450:32:@4832.4]
  wire [31:0] x293_sum_number; // @[Math.scala 154:22:@4873.4 Math.scala 155:14:@4874.4]
  wire [33:0] _GEN_2; // @[Math.scala 450:32:@4878.4]
  wire [33:0] _T_356; // @[Math.scala 450:32:@4878.4]
  wire  _T_388; // @[sm_x300_inr_Foreach.scala 93:131:@4933.4]
  wire  _T_392; // @[package.scala 96:25:@4941.4 package.scala 96:25:@4942.4]
  wire  _T_394; // @[implicits.scala 55:10:@4943.4]
  wire  _T_395; // @[sm_x300_inr_Foreach.scala 93:148:@4944.4]
  wire  _T_397; // @[sm_x300_inr_Foreach.scala 93:236:@4946.4]
  wire  _T_398; // @[sm_x300_inr_Foreach.scala 93:255:@4947.4]
  wire  x560_b289_D4; // @[package.scala 96:25:@4930.4 package.scala 96:25:@4931.4]
  wire  _T_401; // @[sm_x300_inr_Foreach.scala 93:291:@4949.4]
  wire  x559_b290_D4; // @[package.scala 96:25:@4921.4 package.scala 96:25:@4922.4]
  _ _ ( // @[Math.scala 709:24:@4797.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@4809.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x467_sub x467_sub_1 ( // @[Math.scala 191:24:@4836.4]
    .clock(x467_sub_1_clock),
    .reset(x467_sub_1_reset),
    .io_a(x467_sub_1_io_a),
    .io_b(x467_sub_1_io_b),
    .io_flow(x467_sub_1_io_flow),
    .io_result(x467_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@4846.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x292_sum x292_sum_1 ( // @[Math.scala 150:24:@4855.4]
    .clock(x292_sum_1_clock),
    .reset(x292_sum_1_reset),
    .io_a(x292_sum_1_io_a),
    .io_b(x292_sum_1_io_b),
    .io_flow(x292_sum_1_io_flow),
    .io_result(x292_sum_1_io_result)
  );
  x292_sum x293_sum_1 ( // @[Math.scala 150:24:@4867.4]
    .clock(x293_sum_1_clock),
    .reset(x293_sum_1_reset),
    .io_a(x293_sum_1_io_a),
    .io_b(x293_sum_1_io_b),
    .io_flow(x293_sum_1_io_flow),
    .io_result(x293_sum_1_io_result)
  );
  x292_sum x469_sum_1 ( // @[Math.scala 150:24:@4882.4]
    .clock(x469_sum_1_clock),
    .reset(x469_sum_1_reset),
    .io_a(x469_sum_1_io_a),
    .io_b(x469_sum_1_io_b),
    .io_flow(x469_sum_1_io_flow),
    .io_result(x469_sum_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@4916.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_2 ( // @[package.scala 93:22:@4925.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_3 ( // @[package.scala 93:22:@4936.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_327 = ~ io_in_x282_fifoinpacked_0_full; // @[sm_x300_inr_Foreach.scala 62:18:@4822.4]
  assign _T_328 = ~ io_in_x282_fifoinpacked_0_active_0_out; // @[sm_x300_inr_Foreach.scala 62:55:@4823.4]
  assign b287_number = __io_result; // @[Math.scala 712:22:@4802.4 Math.scala 713:14:@4803.4]
  assign _GEN_0 = {{11'd0}, b287_number}; // @[Math.scala 450:32:@4827.4]
  assign _T_332 = _GEN_0 << 11; // @[Math.scala 450:32:@4827.4]
  assign _GEN_1 = {{7'd0}, b287_number}; // @[Math.scala 450:32:@4832.4]
  assign _T_336 = _GEN_1 << 7; // @[Math.scala 450:32:@4832.4]
  assign x293_sum_number = x293_sum_1_io_result; // @[Math.scala 154:22:@4873.4 Math.scala 155:14:@4874.4]
  assign _GEN_2 = {{2'd0}, x293_sum_number}; // @[Math.scala 450:32:@4878.4]
  assign _T_356 = _GEN_2 << 2; // @[Math.scala 450:32:@4878.4]
  assign _T_388 = ~ io_sigsIn_break; // @[sm_x300_inr_Foreach.scala 93:131:@4933.4]
  assign _T_392 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@4941.4 package.scala 96:25:@4942.4]
  assign _T_394 = io_rr ? _T_392 : 1'h0; // @[implicits.scala 55:10:@4943.4]
  assign _T_395 = _T_388 & _T_394; // @[sm_x300_inr_Foreach.scala 93:148:@4944.4]
  assign _T_397 = _T_395 & _T_388; // @[sm_x300_inr_Foreach.scala 93:236:@4946.4]
  assign _T_398 = _T_397 & io_sigsIn_backpressure; // @[sm_x300_inr_Foreach.scala 93:255:@4947.4]
  assign x560_b289_D4 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@4930.4 package.scala 96:25:@4931.4]
  assign _T_401 = _T_398 & x560_b289_D4; // @[sm_x300_inr_Foreach.scala 93:291:@4949.4]
  assign x559_b290_D4 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@4921.4 package.scala 96:25:@4922.4]
  assign io_in_x282_fifoinpacked_0_wPort_0_en_0 = _T_401 & x559_b290_D4; // @[MemInterfaceType.scala 93:57:@4953.4]
  assign io_in_x282_fifoinpacked_0_active_0_in = x560_b289_D4 & x559_b290_D4; // @[MemInterfaceType.scala 147:18:@4956.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@4800.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@4812.4]
  assign x467_sub_1_clock = clock; // @[:@4837.4]
  assign x467_sub_1_reset = reset; // @[:@4838.4]
  assign x467_sub_1_io_a = _T_332[31:0]; // @[Math.scala 192:17:@4839.4]
  assign x467_sub_1_io_b = _T_336[31:0]; // @[Math.scala 193:17:@4840.4]
  assign x467_sub_1_io_flow = _T_327 | _T_328; // @[Math.scala 194:20:@4841.4]
  assign RetimeWrapper_clock = clock; // @[:@4847.4]
  assign RetimeWrapper_reset = reset; // @[:@4848.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4850.4]
  assign RetimeWrapper_io_in = __1_io_result; // @[package.scala 94:16:@4849.4]
  assign x292_sum_1_clock = clock; // @[:@4856.4]
  assign x292_sum_1_reset = reset; // @[:@4857.4]
  assign x292_sum_1_io_a = x467_sub_1_io_result; // @[Math.scala 151:17:@4858.4]
  assign x292_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@4859.4]
  assign x292_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4860.4]
  assign x293_sum_1_clock = clock; // @[:@4868.4]
  assign x293_sum_1_reset = reset; // @[:@4869.4]
  assign x293_sum_1_io_a = x292_sum_1_io_result; // @[Math.scala 151:17:@4870.4]
  assign x293_sum_1_io_b = 32'h1; // @[Math.scala 152:17:@4871.4]
  assign x293_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4872.4]
  assign x469_sum_1_clock = clock; // @[:@4883.4]
  assign x469_sum_1_reset = reset; // @[:@4884.4]
  assign x469_sum_1_io_a = _T_356[31:0]; // @[Math.scala 151:17:@4885.4]
  assign x469_sum_1_io_b = x293_sum_1_io_result; // @[Math.scala 152:17:@4886.4]
  assign x469_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4887.4]
  assign RetimeWrapper_1_clock = clock; // @[:@4917.4]
  assign RetimeWrapper_1_reset = reset; // @[:@4918.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4920.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@4919.4]
  assign RetimeWrapper_2_clock = clock; // @[:@4926.4]
  assign RetimeWrapper_2_reset = reset; // @[:@4927.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4929.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@4928.4]
  assign RetimeWrapper_3_clock = clock; // @[:@4937.4]
  assign RetimeWrapper_3_reset = reset; // @[:@4938.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4940.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@4939.4]
endmodule
module RetimeWrapper_42( // @[:@6074.2]
  input   clock, // @[:@6075.4]
  input   reset, // @[:@6076.4]
  input   io_flow, // @[:@6077.4]
  input   io_in, // @[:@6077.4]
  output  io_out // @[:@6077.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6079.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6079.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6079.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6079.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6079.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6079.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(52)) sr ( // @[RetimeShiftRegister.scala 15:20:@6079.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6092.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6091.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6090.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6089.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6088.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6086.4]
endmodule
module RetimeWrapper_46( // @[:@6202.2]
  input   clock, // @[:@6203.4]
  input   reset, // @[:@6204.4]
  input   io_flow, // @[:@6205.4]
  input   io_in, // @[:@6205.4]
  output  io_out // @[:@6205.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6207.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6207.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6207.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6207.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6207.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6207.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(51)) sr ( // @[RetimeShiftRegister.scala 15:20:@6207.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6220.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6219.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6218.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6217.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6216.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6214.4]
endmodule
module x416_inr_Foreach_SAMPLER_BOX_sm( // @[:@6222.2]
  input   clock, // @[:@6223.4]
  input   reset, // @[:@6224.4]
  input   io_enable, // @[:@6225.4]
  output  io_done, // @[:@6225.4]
  output  io_doneLatch, // @[:@6225.4]
  input   io_ctrDone, // @[:@6225.4]
  output  io_datapathEn, // @[:@6225.4]
  output  io_ctrInc, // @[:@6225.4]
  output  io_ctrRst, // @[:@6225.4]
  input   io_parentAck, // @[:@6225.4]
  input   io_backpressure, // @[:@6225.4]
  input   io_break // @[:@6225.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@6227.4]
  wire  active_reset; // @[Controllers.scala 261:22:@6227.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@6227.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@6227.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@6227.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@6227.4]
  wire  done_clock; // @[Controllers.scala 262:20:@6230.4]
  wire  done_reset; // @[Controllers.scala 262:20:@6230.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@6230.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@6230.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@6230.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@6230.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6264.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6264.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6264.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@6264.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@6264.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6286.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6286.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6286.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6286.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6286.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6298.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6298.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6298.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6298.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6298.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6306.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6306.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6306.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6306.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6306.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@6322.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@6322.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@6322.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@6322.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@6322.4]
  wire  _T_80; // @[Controllers.scala 264:48:@6235.4]
  wire  _T_81; // @[Controllers.scala 264:46:@6236.4]
  wire  _T_82; // @[Controllers.scala 264:62:@6237.4]
  wire  _T_83; // @[Controllers.scala 264:60:@6238.4]
  wire  _T_100; // @[package.scala 100:49:@6255.4]
  reg  _T_103; // @[package.scala 48:56:@6256.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@6269.4 package.scala 96:25:@6270.4]
  wire  _T_110; // @[package.scala 100:49:@6271.4]
  reg  _T_113; // @[package.scala 48:56:@6272.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@6274.4]
  wire  _T_118; // @[Controllers.scala 283:41:@6279.4]
  wire  _T_119; // @[Controllers.scala 283:59:@6280.4]
  wire  _T_121; // @[Controllers.scala 284:37:@6283.4]
  wire  _T_124; // @[package.scala 96:25:@6291.4 package.scala 96:25:@6292.4]
  wire  _T_126; // @[package.scala 100:49:@6293.4]
  reg  _T_129; // @[package.scala 48:56:@6294.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@6316.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@6318.4]
  reg  _T_153; // @[package.scala 48:56:@6319.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@6327.4 package.scala 96:25:@6328.4]
  wire  _T_158; // @[Controllers.scala 292:61:@6329.4]
  wire  _T_159; // @[Controllers.scala 292:24:@6330.4]
  SRFF active ( // @[Controllers.scala 261:22:@6227.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@6230.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_42 RetimeWrapper ( // @[package.scala 93:22:@6264.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_42 RetimeWrapper_1 ( // @[package.scala 93:22:@6286.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@6298.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@6306.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_46 RetimeWrapper_4 ( // @[package.scala 93:22:@6322.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@6235.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@6236.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@6237.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@6238.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@6255.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@6269.4 package.scala 96:25:@6270.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@6271.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@6274.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@6279.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@6280.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@6283.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6291.4 package.scala 96:25:@6292.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@6293.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@6318.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@6327.4 package.scala 96:25:@6328.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@6329.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@6330.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@6297.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@6332.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@6282.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@6285.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@6277.4]
  assign active_clock = clock; // @[:@6228.4]
  assign active_reset = reset; // @[:@6229.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@6240.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@6244.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@6245.4]
  assign done_clock = clock; // @[:@6231.4]
  assign done_reset = reset; // @[:@6232.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@6260.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@6253.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@6254.4]
  assign RetimeWrapper_clock = clock; // @[:@6265.4]
  assign RetimeWrapper_reset = reset; // @[:@6266.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@6268.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@6267.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6287.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6288.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@6290.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@6289.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6299.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6300.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@6302.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@6301.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6307.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6308.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@6310.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@6309.4]
  assign RetimeWrapper_4_clock = clock; // @[:@6323.4]
  assign RetimeWrapper_4_reset = reset; // @[:@6324.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@6326.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@6325.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module RetimeWrapper_50( // @[:@6533.2]
  input        clock, // @[:@6534.4]
  input        reset, // @[:@6535.4]
  input        io_flow, // @[:@6536.4]
  input  [7:0] io_in, // @[:@6536.4]
  output [7:0] io_out // @[:@6536.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@6538.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@6538.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@6538.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6538.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6538.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6538.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@6538.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6551.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6550.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@6549.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6548.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6547.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6545.4]
endmodule
module SRAM_1( // @[:@6569.2]
  input        clock, // @[:@6570.4]
  input  [9:0] io_raddr, // @[:@6572.4]
  input        io_wen, // @[:@6572.4]
  input  [9:0] io_waddr, // @[:@6572.4]
  input  [7:0] io_wdata, // @[:@6572.4]
  output [7:0] io_rdata, // @[:@6572.4]
  input        io_backpressure // @[:@6572.4]
);
  wire [7:0] SRAMVerilogSim_rdata; // @[SRAM.scala 185:23:@6574.4]
  wire [7:0] SRAMVerilogSim_wdata; // @[SRAM.scala 185:23:@6574.4]
  wire  SRAMVerilogSim_backpressure; // @[SRAM.scala 185:23:@6574.4]
  wire  SRAMVerilogSim_wen; // @[SRAM.scala 185:23:@6574.4]
  wire  SRAMVerilogSim_waddrEn; // @[SRAM.scala 185:23:@6574.4]
  wire  SRAMVerilogSim_raddrEn; // @[SRAM.scala 185:23:@6574.4]
  wire [9:0] SRAMVerilogSim_waddr; // @[SRAM.scala 185:23:@6574.4]
  wire [9:0] SRAMVerilogSim_raddr; // @[SRAM.scala 185:23:@6574.4]
  wire  SRAMVerilogSim_clk; // @[SRAM.scala 185:23:@6574.4]
  SRAMVerilogSim #(.DWIDTH(8), .WORDS(640), .AWIDTH(10)) SRAMVerilogSim ( // @[SRAM.scala 185:23:@6574.4]
    .rdata(SRAMVerilogSim_rdata),
    .wdata(SRAMVerilogSim_wdata),
    .backpressure(SRAMVerilogSim_backpressure),
    .wen(SRAMVerilogSim_wen),
    .waddrEn(SRAMVerilogSim_waddrEn),
    .raddrEn(SRAMVerilogSim_raddrEn),
    .waddr(SRAMVerilogSim_waddr),
    .raddr(SRAMVerilogSim_raddr),
    .clk(SRAMVerilogSim_clk)
  );
  assign io_rdata = SRAMVerilogSim_rdata; // @[SRAM.scala 195:16:@6594.4]
  assign SRAMVerilogSim_wdata = io_wdata; // @[SRAM.scala 190:20:@6588.4]
  assign SRAMVerilogSim_backpressure = io_backpressure; // @[SRAM.scala 191:27:@6589.4]
  assign SRAMVerilogSim_wen = io_wen; // @[SRAM.scala 188:18:@6586.4]
  assign SRAMVerilogSim_waddrEn = 1'h1; // @[SRAM.scala 193:22:@6591.4]
  assign SRAMVerilogSim_raddrEn = 1'h1; // @[SRAM.scala 192:22:@6590.4]
  assign SRAMVerilogSim_waddr = io_waddr; // @[SRAM.scala 189:20:@6587.4]
  assign SRAMVerilogSim_raddr = io_raddr; // @[SRAM.scala 187:20:@6585.4]
  assign SRAMVerilogSim_clk = clock; // @[SRAM.scala 186:18:@6584.4]
endmodule
module RetimeWrapper_51( // @[:@6608.2]
  input        clock, // @[:@6609.4]
  input        reset, // @[:@6610.4]
  input        io_flow, // @[:@6611.4]
  input  [9:0] io_in, // @[:@6611.4]
  output [9:0] io_out // @[:@6611.4]
);
  wire [9:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@6613.4]
  wire [9:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@6613.4]
  wire [9:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@6613.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6613.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6613.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6613.4]
  RetimeShiftRegister #(.WIDTH(10), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@6613.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6626.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6625.4]
  assign sr_init = 10'h0; // @[RetimeShiftRegister.scala 19:16:@6624.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6623.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6622.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6620.4]
endmodule
module Mem1D_5( // @[:@6628.2]
  input        clock, // @[:@6629.4]
  input        reset, // @[:@6630.4]
  input  [9:0] io_r_ofs_0, // @[:@6631.4]
  input        io_r_backpressure, // @[:@6631.4]
  input  [9:0] io_w_ofs_0, // @[:@6631.4]
  input  [7:0] io_w_data_0, // @[:@6631.4]
  input        io_w_en_0, // @[:@6631.4]
  output [7:0] io_output // @[:@6631.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 705:21:@6635.4]
  wire [9:0] SRAM_io_raddr; // @[MemPrimitives.scala 705:21:@6635.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 705:21:@6635.4]
  wire [9:0] SRAM_io_waddr; // @[MemPrimitives.scala 705:21:@6635.4]
  wire [7:0] SRAM_io_wdata; // @[MemPrimitives.scala 705:21:@6635.4]
  wire [7:0] SRAM_io_rdata; // @[MemPrimitives.scala 705:21:@6635.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 705:21:@6635.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6638.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6638.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6638.4]
  wire [9:0] RetimeWrapper_io_in; // @[package.scala 93:22:@6638.4]
  wire [9:0] RetimeWrapper_io_out; // @[package.scala 93:22:@6638.4]
  wire  wInBound; // @[MemPrimitives.scala 692:32:@6633.4]
  SRAM_1 SRAM ( // @[MemPrimitives.scala 705:21:@6635.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_51 RetimeWrapper ( // @[package.scala 93:22:@6638.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 10'h280; // @[MemPrimitives.scala 692:32:@6633.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 712:17:@6651.4]
  assign SRAM_clock = clock; // @[:@6636.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 706:37:@6645.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 709:22:@6648.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 708:22:@6646.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 710:22:@6649.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 711:30:@6650.4]
  assign RetimeWrapper_clock = clock; // @[:@6639.4]
  assign RetimeWrapper_reset = reset; // @[:@6640.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@6642.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@6641.4]
endmodule
module StickySelects_1( // @[:@7753.2]
  input   clock, // @[:@7754.4]
  input   reset, // @[:@7755.4]
  input   io_ins_0, // @[:@7756.4]
  input   io_ins_1, // @[:@7756.4]
  input   io_ins_2, // @[:@7756.4]
  input   io_ins_3, // @[:@7756.4]
  input   io_ins_4, // @[:@7756.4]
  input   io_ins_5, // @[:@7756.4]
  input   io_ins_6, // @[:@7756.4]
  input   io_ins_7, // @[:@7756.4]
  input   io_ins_8, // @[:@7756.4]
  output  io_outs_0, // @[:@7756.4]
  output  io_outs_1, // @[:@7756.4]
  output  io_outs_2, // @[:@7756.4]
  output  io_outs_3, // @[:@7756.4]
  output  io_outs_4, // @[:@7756.4]
  output  io_outs_5, // @[:@7756.4]
  output  io_outs_6, // @[:@7756.4]
  output  io_outs_7, // @[:@7756.4]
  output  io_outs_8 // @[:@7756.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@7758.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@7759.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@7760.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@7761.4]
  reg [31:0] _RAND_3;
  reg  _T_31; // @[StickySelects.scala 37:46:@7762.4]
  reg [31:0] _RAND_4;
  reg  _T_34; // @[StickySelects.scala 37:46:@7763.4]
  reg [31:0] _RAND_5;
  reg  _T_37; // @[StickySelects.scala 37:46:@7764.4]
  reg [31:0] _RAND_6;
  reg  _T_40; // @[StickySelects.scala 37:46:@7765.4]
  reg [31:0] _RAND_7;
  reg  _T_43; // @[StickySelects.scala 37:46:@7766.4]
  reg [31:0] _RAND_8;
  wire  _T_44; // @[StickySelects.scala 47:46:@7767.4]
  wire  _T_45; // @[StickySelects.scala 47:46:@7768.4]
  wire  _T_46; // @[StickySelects.scala 47:46:@7769.4]
  wire  _T_47; // @[StickySelects.scala 47:46:@7770.4]
  wire  _T_48; // @[StickySelects.scala 47:46:@7771.4]
  wire  _T_49; // @[StickySelects.scala 47:46:@7772.4]
  wire  _T_50; // @[StickySelects.scala 47:46:@7773.4]
  wire  _T_51; // @[StickySelects.scala 49:53:@7774.4]
  wire  _T_52; // @[StickySelects.scala 49:21:@7775.4]
  wire  _T_53; // @[StickySelects.scala 47:46:@7777.4]
  wire  _T_54; // @[StickySelects.scala 47:46:@7778.4]
  wire  _T_55; // @[StickySelects.scala 47:46:@7779.4]
  wire  _T_56; // @[StickySelects.scala 47:46:@7780.4]
  wire  _T_57; // @[StickySelects.scala 47:46:@7781.4]
  wire  _T_58; // @[StickySelects.scala 47:46:@7782.4]
  wire  _T_59; // @[StickySelects.scala 47:46:@7783.4]
  wire  _T_60; // @[StickySelects.scala 49:53:@7784.4]
  wire  _T_61; // @[StickySelects.scala 49:21:@7785.4]
  wire  _T_62; // @[StickySelects.scala 47:46:@7787.4]
  wire  _T_63; // @[StickySelects.scala 47:46:@7788.4]
  wire  _T_64; // @[StickySelects.scala 47:46:@7789.4]
  wire  _T_65; // @[StickySelects.scala 47:46:@7790.4]
  wire  _T_66; // @[StickySelects.scala 47:46:@7791.4]
  wire  _T_67; // @[StickySelects.scala 47:46:@7792.4]
  wire  _T_68; // @[StickySelects.scala 47:46:@7793.4]
  wire  _T_69; // @[StickySelects.scala 49:53:@7794.4]
  wire  _T_70; // @[StickySelects.scala 49:21:@7795.4]
  wire  _T_72; // @[StickySelects.scala 47:46:@7798.4]
  wire  _T_73; // @[StickySelects.scala 47:46:@7799.4]
  wire  _T_74; // @[StickySelects.scala 47:46:@7800.4]
  wire  _T_75; // @[StickySelects.scala 47:46:@7801.4]
  wire  _T_76; // @[StickySelects.scala 47:46:@7802.4]
  wire  _T_77; // @[StickySelects.scala 47:46:@7803.4]
  wire  _T_78; // @[StickySelects.scala 49:53:@7804.4]
  wire  _T_79; // @[StickySelects.scala 49:21:@7805.4]
  wire  _T_82; // @[StickySelects.scala 47:46:@7809.4]
  wire  _T_83; // @[StickySelects.scala 47:46:@7810.4]
  wire  _T_84; // @[StickySelects.scala 47:46:@7811.4]
  wire  _T_85; // @[StickySelects.scala 47:46:@7812.4]
  wire  _T_86; // @[StickySelects.scala 47:46:@7813.4]
  wire  _T_87; // @[StickySelects.scala 49:53:@7814.4]
  wire  _T_88; // @[StickySelects.scala 49:21:@7815.4]
  wire  _T_92; // @[StickySelects.scala 47:46:@7820.4]
  wire  _T_93; // @[StickySelects.scala 47:46:@7821.4]
  wire  _T_94; // @[StickySelects.scala 47:46:@7822.4]
  wire  _T_95; // @[StickySelects.scala 47:46:@7823.4]
  wire  _T_96; // @[StickySelects.scala 49:53:@7824.4]
  wire  _T_97; // @[StickySelects.scala 49:21:@7825.4]
  wire  _T_102; // @[StickySelects.scala 47:46:@7831.4]
  wire  _T_103; // @[StickySelects.scala 47:46:@7832.4]
  wire  _T_104; // @[StickySelects.scala 47:46:@7833.4]
  wire  _T_105; // @[StickySelects.scala 49:53:@7834.4]
  wire  _T_106; // @[StickySelects.scala 49:21:@7835.4]
  wire  _T_112; // @[StickySelects.scala 47:46:@7842.4]
  wire  _T_113; // @[StickySelects.scala 47:46:@7843.4]
  wire  _T_114; // @[StickySelects.scala 49:53:@7844.4]
  wire  _T_115; // @[StickySelects.scala 49:21:@7845.4]
  wire  _T_122; // @[StickySelects.scala 47:46:@7853.4]
  wire  _T_123; // @[StickySelects.scala 49:53:@7854.4]
  wire  _T_124; // @[StickySelects.scala 49:21:@7855.4]
  assign _T_44 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@7767.4]
  assign _T_45 = _T_44 | io_ins_3; // @[StickySelects.scala 47:46:@7768.4]
  assign _T_46 = _T_45 | io_ins_4; // @[StickySelects.scala 47:46:@7769.4]
  assign _T_47 = _T_46 | io_ins_5; // @[StickySelects.scala 47:46:@7770.4]
  assign _T_48 = _T_47 | io_ins_6; // @[StickySelects.scala 47:46:@7771.4]
  assign _T_49 = _T_48 | io_ins_7; // @[StickySelects.scala 47:46:@7772.4]
  assign _T_50 = _T_49 | io_ins_8; // @[StickySelects.scala 47:46:@7773.4]
  assign _T_51 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@7774.4]
  assign _T_52 = _T_50 ? io_ins_0 : _T_51; // @[StickySelects.scala 49:21:@7775.4]
  assign _T_53 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@7777.4]
  assign _T_54 = _T_53 | io_ins_3; // @[StickySelects.scala 47:46:@7778.4]
  assign _T_55 = _T_54 | io_ins_4; // @[StickySelects.scala 47:46:@7779.4]
  assign _T_56 = _T_55 | io_ins_5; // @[StickySelects.scala 47:46:@7780.4]
  assign _T_57 = _T_56 | io_ins_6; // @[StickySelects.scala 47:46:@7781.4]
  assign _T_58 = _T_57 | io_ins_7; // @[StickySelects.scala 47:46:@7782.4]
  assign _T_59 = _T_58 | io_ins_8; // @[StickySelects.scala 47:46:@7783.4]
  assign _T_60 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@7784.4]
  assign _T_61 = _T_59 ? io_ins_1 : _T_60; // @[StickySelects.scala 49:21:@7785.4]
  assign _T_62 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@7787.4]
  assign _T_63 = _T_62 | io_ins_3; // @[StickySelects.scala 47:46:@7788.4]
  assign _T_64 = _T_63 | io_ins_4; // @[StickySelects.scala 47:46:@7789.4]
  assign _T_65 = _T_64 | io_ins_5; // @[StickySelects.scala 47:46:@7790.4]
  assign _T_66 = _T_65 | io_ins_6; // @[StickySelects.scala 47:46:@7791.4]
  assign _T_67 = _T_66 | io_ins_7; // @[StickySelects.scala 47:46:@7792.4]
  assign _T_68 = _T_67 | io_ins_8; // @[StickySelects.scala 47:46:@7793.4]
  assign _T_69 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@7794.4]
  assign _T_70 = _T_68 ? io_ins_2 : _T_69; // @[StickySelects.scala 49:21:@7795.4]
  assign _T_72 = _T_62 | io_ins_2; // @[StickySelects.scala 47:46:@7798.4]
  assign _T_73 = _T_72 | io_ins_4; // @[StickySelects.scala 47:46:@7799.4]
  assign _T_74 = _T_73 | io_ins_5; // @[StickySelects.scala 47:46:@7800.4]
  assign _T_75 = _T_74 | io_ins_6; // @[StickySelects.scala 47:46:@7801.4]
  assign _T_76 = _T_75 | io_ins_7; // @[StickySelects.scala 47:46:@7802.4]
  assign _T_77 = _T_76 | io_ins_8; // @[StickySelects.scala 47:46:@7803.4]
  assign _T_78 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@7804.4]
  assign _T_79 = _T_77 ? io_ins_3 : _T_78; // @[StickySelects.scala 49:21:@7805.4]
  assign _T_82 = _T_72 | io_ins_3; // @[StickySelects.scala 47:46:@7809.4]
  assign _T_83 = _T_82 | io_ins_5; // @[StickySelects.scala 47:46:@7810.4]
  assign _T_84 = _T_83 | io_ins_6; // @[StickySelects.scala 47:46:@7811.4]
  assign _T_85 = _T_84 | io_ins_7; // @[StickySelects.scala 47:46:@7812.4]
  assign _T_86 = _T_85 | io_ins_8; // @[StickySelects.scala 47:46:@7813.4]
  assign _T_87 = io_ins_4 | _T_31; // @[StickySelects.scala 49:53:@7814.4]
  assign _T_88 = _T_86 ? io_ins_4 : _T_87; // @[StickySelects.scala 49:21:@7815.4]
  assign _T_92 = _T_82 | io_ins_4; // @[StickySelects.scala 47:46:@7820.4]
  assign _T_93 = _T_92 | io_ins_6; // @[StickySelects.scala 47:46:@7821.4]
  assign _T_94 = _T_93 | io_ins_7; // @[StickySelects.scala 47:46:@7822.4]
  assign _T_95 = _T_94 | io_ins_8; // @[StickySelects.scala 47:46:@7823.4]
  assign _T_96 = io_ins_5 | _T_34; // @[StickySelects.scala 49:53:@7824.4]
  assign _T_97 = _T_95 ? io_ins_5 : _T_96; // @[StickySelects.scala 49:21:@7825.4]
  assign _T_102 = _T_92 | io_ins_5; // @[StickySelects.scala 47:46:@7831.4]
  assign _T_103 = _T_102 | io_ins_7; // @[StickySelects.scala 47:46:@7832.4]
  assign _T_104 = _T_103 | io_ins_8; // @[StickySelects.scala 47:46:@7833.4]
  assign _T_105 = io_ins_6 | _T_37; // @[StickySelects.scala 49:53:@7834.4]
  assign _T_106 = _T_104 ? io_ins_6 : _T_105; // @[StickySelects.scala 49:21:@7835.4]
  assign _T_112 = _T_102 | io_ins_6; // @[StickySelects.scala 47:46:@7842.4]
  assign _T_113 = _T_112 | io_ins_8; // @[StickySelects.scala 47:46:@7843.4]
  assign _T_114 = io_ins_7 | _T_40; // @[StickySelects.scala 49:53:@7844.4]
  assign _T_115 = _T_113 ? io_ins_7 : _T_114; // @[StickySelects.scala 49:21:@7845.4]
  assign _T_122 = _T_112 | io_ins_7; // @[StickySelects.scala 47:46:@7853.4]
  assign _T_123 = io_ins_8 | _T_43; // @[StickySelects.scala 49:53:@7854.4]
  assign _T_124 = _T_122 ? io_ins_8 : _T_123; // @[StickySelects.scala 49:21:@7855.4]
  assign io_outs_0 = _T_50 ? io_ins_0 : _T_51; // @[StickySelects.scala 53:57:@7857.4]
  assign io_outs_1 = _T_59 ? io_ins_1 : _T_60; // @[StickySelects.scala 53:57:@7858.4]
  assign io_outs_2 = _T_68 ? io_ins_2 : _T_69; // @[StickySelects.scala 53:57:@7859.4]
  assign io_outs_3 = _T_77 ? io_ins_3 : _T_78; // @[StickySelects.scala 53:57:@7860.4]
  assign io_outs_4 = _T_86 ? io_ins_4 : _T_87; // @[StickySelects.scala 53:57:@7861.4]
  assign io_outs_5 = _T_95 ? io_ins_5 : _T_96; // @[StickySelects.scala 53:57:@7862.4]
  assign io_outs_6 = _T_104 ? io_ins_6 : _T_105; // @[StickySelects.scala 53:57:@7863.4]
  assign io_outs_7 = _T_113 ? io_ins_7 : _T_114; // @[StickySelects.scala 53:57:@7864.4]
  assign io_outs_8 = _T_122 ? io_ins_8 : _T_123; // @[StickySelects.scala 53:57:@7865.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_31 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_37 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_40 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_43 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_50) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_51;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_59) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_60;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_68) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_69;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_77) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_78;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_86) begin
        _T_31 <= io_ins_4;
      end else begin
        _T_31 <= _T_87;
      end
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (_T_95) begin
        _T_34 <= io_ins_5;
      end else begin
        _T_34 <= _T_96;
      end
    end
    if (reset) begin
      _T_37 <= 1'h0;
    end else begin
      if (_T_104) begin
        _T_37 <= io_ins_6;
      end else begin
        _T_37 <= _T_105;
      end
    end
    if (reset) begin
      _T_40 <= 1'h0;
    end else begin
      if (_T_113) begin
        _T_40 <= io_ins_7;
      end else begin
        _T_40 <= _T_114;
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_122) begin
        _T_43 <= io_ins_8;
      end else begin
        _T_43 <= _T_123;
      end
    end
  end
endmodule
module x311_lb_0( // @[:@12577.2]
  input        clock, // @[:@12578.4]
  input        reset, // @[:@12579.4]
  input  [1:0] io_rPort_8_banks_1, // @[:@12580.4]
  input  [2:0] io_rPort_8_banks_0, // @[:@12580.4]
  input  [9:0] io_rPort_8_ofs_0, // @[:@12580.4]
  input        io_rPort_8_en_0, // @[:@12580.4]
  input        io_rPort_8_backpressure, // @[:@12580.4]
  output [7:0] io_rPort_8_output_0, // @[:@12580.4]
  input  [1:0] io_rPort_7_banks_1, // @[:@12580.4]
  input  [2:0] io_rPort_7_banks_0, // @[:@12580.4]
  input  [9:0] io_rPort_7_ofs_0, // @[:@12580.4]
  input        io_rPort_7_en_0, // @[:@12580.4]
  input        io_rPort_7_backpressure, // @[:@12580.4]
  output [7:0] io_rPort_7_output_0, // @[:@12580.4]
  input  [1:0] io_rPort_6_banks_1, // @[:@12580.4]
  input  [2:0] io_rPort_6_banks_0, // @[:@12580.4]
  input  [9:0] io_rPort_6_ofs_0, // @[:@12580.4]
  input        io_rPort_6_en_0, // @[:@12580.4]
  input        io_rPort_6_backpressure, // @[:@12580.4]
  output [7:0] io_rPort_6_output_0, // @[:@12580.4]
  input  [1:0] io_rPort_5_banks_1, // @[:@12580.4]
  input  [2:0] io_rPort_5_banks_0, // @[:@12580.4]
  input  [9:0] io_rPort_5_ofs_0, // @[:@12580.4]
  input        io_rPort_5_en_0, // @[:@12580.4]
  input        io_rPort_5_backpressure, // @[:@12580.4]
  output [7:0] io_rPort_5_output_0, // @[:@12580.4]
  input  [1:0] io_rPort_4_banks_1, // @[:@12580.4]
  input  [2:0] io_rPort_4_banks_0, // @[:@12580.4]
  input  [9:0] io_rPort_4_ofs_0, // @[:@12580.4]
  input        io_rPort_4_en_0, // @[:@12580.4]
  input        io_rPort_4_backpressure, // @[:@12580.4]
  output [7:0] io_rPort_4_output_0, // @[:@12580.4]
  input  [1:0] io_rPort_3_banks_1, // @[:@12580.4]
  input  [2:0] io_rPort_3_banks_0, // @[:@12580.4]
  input  [9:0] io_rPort_3_ofs_0, // @[:@12580.4]
  input        io_rPort_3_en_0, // @[:@12580.4]
  input        io_rPort_3_backpressure, // @[:@12580.4]
  output [7:0] io_rPort_3_output_0, // @[:@12580.4]
  input  [1:0] io_rPort_2_banks_1, // @[:@12580.4]
  input  [2:0] io_rPort_2_banks_0, // @[:@12580.4]
  input  [9:0] io_rPort_2_ofs_0, // @[:@12580.4]
  input        io_rPort_2_en_0, // @[:@12580.4]
  input        io_rPort_2_backpressure, // @[:@12580.4]
  output [7:0] io_rPort_2_output_0, // @[:@12580.4]
  input  [1:0] io_rPort_1_banks_1, // @[:@12580.4]
  input  [2:0] io_rPort_1_banks_0, // @[:@12580.4]
  input  [9:0] io_rPort_1_ofs_0, // @[:@12580.4]
  input        io_rPort_1_en_0, // @[:@12580.4]
  input        io_rPort_1_backpressure, // @[:@12580.4]
  output [7:0] io_rPort_1_output_0, // @[:@12580.4]
  input  [1:0] io_rPort_0_banks_1, // @[:@12580.4]
  input  [2:0] io_rPort_0_banks_0, // @[:@12580.4]
  input  [9:0] io_rPort_0_ofs_0, // @[:@12580.4]
  input        io_rPort_0_en_0, // @[:@12580.4]
  input        io_rPort_0_backpressure, // @[:@12580.4]
  output [7:0] io_rPort_0_output_0, // @[:@12580.4]
  input  [1:0] io_wPort_0_banks_1, // @[:@12580.4]
  input  [2:0] io_wPort_0_banks_0, // @[:@12580.4]
  input  [9:0] io_wPort_0_ofs_0, // @[:@12580.4]
  input  [7:0] io_wPort_0_data_0, // @[:@12580.4]
  input        io_wPort_0_en_0 // @[:@12580.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@12645.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@12645.4]
  wire [9:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12645.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12645.4]
  wire [9:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12645.4]
  wire [7:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@12645.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@12645.4]
  wire [7:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@12645.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@12661.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@12661.4]
  wire [9:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12661.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12661.4]
  wire [9:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12661.4]
  wire [7:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@12661.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@12661.4]
  wire [7:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@12661.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@12677.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@12677.4]
  wire [9:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12677.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12677.4]
  wire [9:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12677.4]
  wire [7:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@12677.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@12677.4]
  wire [7:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@12677.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@12693.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@12693.4]
  wire [9:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12693.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12693.4]
  wire [9:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12693.4]
  wire [7:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@12693.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@12693.4]
  wire [7:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@12693.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@12709.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@12709.4]
  wire [9:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12709.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12709.4]
  wire [9:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12709.4]
  wire [7:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@12709.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@12709.4]
  wire [7:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@12709.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@12725.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@12725.4]
  wire [9:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12725.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12725.4]
  wire [9:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12725.4]
  wire [7:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@12725.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@12725.4]
  wire [7:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@12725.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@12741.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@12741.4]
  wire [9:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12741.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12741.4]
  wire [9:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12741.4]
  wire [7:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@12741.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@12741.4]
  wire [7:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@12741.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@12757.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@12757.4]
  wire [9:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12757.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12757.4]
  wire [9:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12757.4]
  wire [7:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@12757.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@12757.4]
  wire [7:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@12757.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@12773.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@12773.4]
  wire [9:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12773.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12773.4]
  wire [9:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12773.4]
  wire [7:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@12773.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@12773.4]
  wire [7:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@12773.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@12789.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@12789.4]
  wire [9:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12789.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12789.4]
  wire [9:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12789.4]
  wire [7:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@12789.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@12789.4]
  wire [7:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@12789.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@12805.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@12805.4]
  wire [9:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12805.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12805.4]
  wire [9:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12805.4]
  wire [7:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@12805.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@12805.4]
  wire [7:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@12805.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@12821.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@12821.4]
  wire [9:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12821.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12821.4]
  wire [9:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12821.4]
  wire [7:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@12821.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@12821.4]
  wire [7:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@12821.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_io_ins_6; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_io_ins_7; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_io_ins_8; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_io_outs_6; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_io_outs_7; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_io_outs_8; // @[MemPrimitives.scala 121:29:@13017.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_io_ins_6; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_io_ins_7; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_io_ins_8; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_io_outs_6; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_io_outs_7; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_1_io_outs_8; // @[MemPrimitives.scala 121:29:@13106.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_io_ins_6; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_io_ins_7; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_io_ins_8; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_io_outs_6; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_io_outs_7; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_2_io_outs_8; // @[MemPrimitives.scala 121:29:@13195.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_io_ins_6; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_io_ins_7; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_io_ins_8; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_io_outs_6; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_io_outs_7; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_3_io_outs_8; // @[MemPrimitives.scala 121:29:@13284.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_io_ins_6; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_io_ins_7; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_io_ins_8; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_io_outs_6; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_io_outs_7; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_4_io_outs_8; // @[MemPrimitives.scala 121:29:@13373.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_io_ins_6; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_io_ins_7; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_io_ins_8; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_io_outs_6; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_io_outs_7; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_5_io_outs_8; // @[MemPrimitives.scala 121:29:@13462.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_io_ins_6; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_io_ins_7; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_io_ins_8; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_io_outs_6; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_io_outs_7; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_6_io_outs_8; // @[MemPrimitives.scala 121:29:@13551.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_io_ins_6; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_io_ins_7; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_io_ins_8; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_io_outs_6; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_io_outs_7; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_7_io_outs_8; // @[MemPrimitives.scala 121:29:@13640.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_io_ins_6; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_io_ins_7; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_io_ins_8; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_io_outs_6; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_io_outs_7; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_8_io_outs_8; // @[MemPrimitives.scala 121:29:@13729.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_io_ins_6; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_io_ins_7; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_io_ins_8; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_io_outs_6; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_io_outs_7; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_9_io_outs_8; // @[MemPrimitives.scala 121:29:@13818.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_io_ins_6; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_io_ins_7; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_io_ins_8; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_io_outs_6; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_io_outs_7; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_10_io_outs_8; // @[MemPrimitives.scala 121:29:@13907.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_io_ins_6; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_io_ins_7; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_io_ins_8; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_io_outs_6; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_io_outs_7; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  StickySelects_11_io_outs_8; // @[MemPrimitives.scala 121:29:@13996.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@14086.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@14086.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@14086.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@14086.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@14086.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@14094.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@14094.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@14094.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@14094.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@14094.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@14102.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@14102.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@14102.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@14102.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@14102.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@14110.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@14110.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@14110.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@14110.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@14110.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@14118.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@14118.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@14118.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@14118.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@14118.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@14126.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@14126.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@14126.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@14126.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@14126.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@14134.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@14134.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@14134.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@14134.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@14134.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@14142.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@14142.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@14142.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@14142.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@14142.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@14150.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@14150.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@14150.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@14150.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@14150.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@14158.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@14158.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@14158.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@14158.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@14158.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@14166.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@14166.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@14166.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@14166.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@14166.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@14174.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@14174.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@14174.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@14174.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@14174.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@14230.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@14230.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@14230.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@14230.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@14230.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@14238.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@14238.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@14238.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@14238.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@14238.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@14246.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@14246.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@14246.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@14246.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@14246.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@14254.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@14254.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@14254.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@14254.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@14254.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@14262.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@14262.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@14262.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@14262.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@14262.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@14270.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@14270.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@14270.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@14270.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@14270.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@14278.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@14278.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@14278.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@14278.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@14278.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@14286.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@14286.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@14286.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@14286.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@14286.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@14294.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@14294.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@14294.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@14294.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@14294.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@14302.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@14302.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@14302.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@14302.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@14302.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@14310.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@14310.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@14310.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@14310.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@14310.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@14318.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@14318.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@14318.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@14318.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@14318.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@14374.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@14374.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@14374.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@14374.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@14374.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@14382.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@14382.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@14382.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@14382.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@14382.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@14390.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@14390.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@14390.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@14390.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@14390.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@14398.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@14398.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@14398.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@14398.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@14398.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@14406.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@14406.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@14406.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@14406.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@14406.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@14414.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@14414.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@14414.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@14414.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@14414.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@14422.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@14422.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@14422.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@14422.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@14422.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@14430.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@14430.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@14430.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@14430.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@14430.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@14438.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@14438.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@14438.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@14438.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@14438.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@14446.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@14446.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@14446.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@14446.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@14446.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@14454.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@14454.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@14454.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@14454.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@14454.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@14462.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@14462.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@14462.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@14462.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@14462.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@14518.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@14518.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@14518.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@14518.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@14518.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@14526.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@14526.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@14526.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@14526.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@14526.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@14534.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@14534.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@14534.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@14534.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@14534.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@14542.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@14542.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@14542.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@14542.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@14542.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@14550.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@14550.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@14550.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@14550.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@14550.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@14558.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@14558.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@14558.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@14558.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@14558.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@14566.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@14566.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@14566.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@14566.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@14566.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@14574.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@14574.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@14574.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@14574.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@14574.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@14582.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@14582.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@14582.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@14582.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@14582.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@14590.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@14590.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@14590.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@14590.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@14590.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@14598.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@14598.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@14598.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@14598.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@14598.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@14606.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@14606.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@14606.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@14606.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@14606.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@14662.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@14662.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@14662.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@14662.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@14662.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@14670.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@14670.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@14670.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@14670.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@14670.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@14678.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@14678.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@14678.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@14678.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@14678.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@14686.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@14686.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@14686.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@14686.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@14686.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@14694.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@14694.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@14694.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@14694.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@14694.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@14702.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@14702.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@14702.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@14702.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@14702.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@14710.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@14710.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@14710.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@14710.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@14710.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@14718.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@14718.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@14718.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@14718.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@14718.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@14726.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@14726.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@14726.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@14726.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@14726.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@14734.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@14734.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@14734.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@14734.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@14734.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@14742.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@14742.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@14742.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@14742.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@14742.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@14750.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@14750.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@14750.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@14750.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@14750.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@14806.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@14806.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@14806.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@14806.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@14806.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@14814.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@14814.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@14814.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@14814.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@14814.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@14822.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@14822.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@14822.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@14822.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@14822.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@14830.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@14830.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@14830.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@14830.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@14830.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@14838.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@14838.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@14838.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@14838.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@14838.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@14846.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@14846.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@14846.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@14846.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@14846.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@14854.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@14854.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@14854.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@14854.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@14854.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@14862.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@14870.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@14870.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@14870.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@14870.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@14870.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@14878.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@14878.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@14878.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@14878.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@14878.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@14886.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@14886.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@14886.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@14886.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@14886.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@14894.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@14894.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@14894.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@14894.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@14894.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@14950.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@14950.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@14950.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@14950.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@14950.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@14958.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@14966.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@14966.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@14966.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@14966.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@14966.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@14974.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@14974.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@14974.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@14974.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@14974.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@14982.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@14990.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@14990.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@14990.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@14990.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@14990.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@14998.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@14998.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@14998.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@14998.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@14998.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@15006.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@15006.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@15006.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@15006.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@15006.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@15014.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@15014.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@15014.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@15014.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@15014.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@15022.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@15022.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@15022.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@15022.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@15022.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@15030.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@15030.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@15030.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@15030.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@15030.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@15038.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@15038.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@15038.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@15038.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@15038.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@15094.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@15094.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@15094.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@15094.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@15094.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@15102.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@15102.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@15102.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@15102.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@15102.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@15110.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@15110.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@15110.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@15110.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@15110.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@15118.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@15118.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@15118.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@15118.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@15118.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@15126.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@15126.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@15126.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@15126.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@15126.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@15134.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@15134.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@15134.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@15134.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@15134.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@15142.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@15142.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@15142.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@15142.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@15142.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@15150.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@15150.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@15150.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@15150.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@15150.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@15158.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@15158.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@15158.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@15158.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@15158.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@15166.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@15166.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@15166.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@15166.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@15166.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@15174.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@15174.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@15174.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@15174.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@15174.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@15182.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@15182.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@15182.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@15182.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@15182.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@15238.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@15238.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@15238.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@15238.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@15238.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@15246.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@15246.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@15246.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@15246.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@15246.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@15254.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@15254.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@15254.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@15254.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@15254.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@15262.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@15262.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@15262.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@15262.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@15262.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@15270.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@15270.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@15270.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@15270.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@15270.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@15278.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@15278.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@15278.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@15278.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@15278.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@15286.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@15286.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@15286.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@15286.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@15286.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@15294.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@15294.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@15294.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@15294.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@15294.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@15302.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@15302.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@15302.4]
  wire  RetimeWrapper_104_io_in; // @[package.scala 93:22:@15302.4]
  wire  RetimeWrapper_104_io_out; // @[package.scala 93:22:@15302.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@15310.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@15310.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@15310.4]
  wire  RetimeWrapper_105_io_in; // @[package.scala 93:22:@15310.4]
  wire  RetimeWrapper_105_io_out; // @[package.scala 93:22:@15310.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@15318.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@15318.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@15318.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@15318.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@15318.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@15326.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@15326.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@15326.4]
  wire  RetimeWrapper_107_io_in; // @[package.scala 93:22:@15326.4]
  wire  RetimeWrapper_107_io_out; // @[package.scala 93:22:@15326.4]
  wire  _T_316; // @[MemPrimitives.scala 82:210:@12837.4]
  wire  _T_318; // @[MemPrimitives.scala 82:210:@12838.4]
  wire  _T_319; // @[MemPrimitives.scala 82:228:@12839.4]
  wire  _T_320; // @[MemPrimitives.scala 83:102:@12840.4]
  wire [18:0] _T_322; // @[Cat.scala 30:58:@12842.4]
  wire  _T_329; // @[MemPrimitives.scala 82:210:@12850.4]
  wire  _T_330; // @[MemPrimitives.scala 82:228:@12851.4]
  wire  _T_331; // @[MemPrimitives.scala 83:102:@12852.4]
  wire [18:0] _T_333; // @[Cat.scala 30:58:@12854.4]
  wire  _T_340; // @[MemPrimitives.scala 82:210:@12862.4]
  wire  _T_341; // @[MemPrimitives.scala 82:228:@12863.4]
  wire  _T_342; // @[MemPrimitives.scala 83:102:@12864.4]
  wire [18:0] _T_344; // @[Cat.scala 30:58:@12866.4]
  wire  _T_349; // @[MemPrimitives.scala 82:210:@12873.4]
  wire  _T_352; // @[MemPrimitives.scala 82:228:@12875.4]
  wire  _T_353; // @[MemPrimitives.scala 83:102:@12876.4]
  wire [18:0] _T_355; // @[Cat.scala 30:58:@12878.4]
  wire  _T_363; // @[MemPrimitives.scala 82:228:@12887.4]
  wire  _T_364; // @[MemPrimitives.scala 83:102:@12888.4]
  wire [18:0] _T_366; // @[Cat.scala 30:58:@12890.4]
  wire  _T_374; // @[MemPrimitives.scala 82:228:@12899.4]
  wire  _T_375; // @[MemPrimitives.scala 83:102:@12900.4]
  wire [18:0] _T_377; // @[Cat.scala 30:58:@12902.4]
  wire  _T_382; // @[MemPrimitives.scala 82:210:@12909.4]
  wire  _T_385; // @[MemPrimitives.scala 82:228:@12911.4]
  wire  _T_386; // @[MemPrimitives.scala 83:102:@12912.4]
  wire [18:0] _T_388; // @[Cat.scala 30:58:@12914.4]
  wire  _T_396; // @[MemPrimitives.scala 82:228:@12923.4]
  wire  _T_397; // @[MemPrimitives.scala 83:102:@12924.4]
  wire [18:0] _T_399; // @[Cat.scala 30:58:@12926.4]
  wire  _T_407; // @[MemPrimitives.scala 82:228:@12935.4]
  wire  _T_408; // @[MemPrimitives.scala 83:102:@12936.4]
  wire [18:0] _T_410; // @[Cat.scala 30:58:@12938.4]
  wire  _T_415; // @[MemPrimitives.scala 82:210:@12945.4]
  wire  _T_418; // @[MemPrimitives.scala 82:228:@12947.4]
  wire  _T_419; // @[MemPrimitives.scala 83:102:@12948.4]
  wire [18:0] _T_421; // @[Cat.scala 30:58:@12950.4]
  wire  _T_429; // @[MemPrimitives.scala 82:228:@12959.4]
  wire  _T_430; // @[MemPrimitives.scala 83:102:@12960.4]
  wire [18:0] _T_432; // @[Cat.scala 30:58:@12962.4]
  wire  _T_440; // @[MemPrimitives.scala 82:228:@12971.4]
  wire  _T_441; // @[MemPrimitives.scala 83:102:@12972.4]
  wire [18:0] _T_443; // @[Cat.scala 30:58:@12974.4]
  wire  _T_448; // @[MemPrimitives.scala 110:210:@12981.4]
  wire  _T_450; // @[MemPrimitives.scala 110:210:@12982.4]
  wire  _T_451; // @[MemPrimitives.scala 110:228:@12983.4]
  wire  _T_454; // @[MemPrimitives.scala 110:210:@12985.4]
  wire  _T_456; // @[MemPrimitives.scala 110:210:@12986.4]
  wire  _T_457; // @[MemPrimitives.scala 110:228:@12987.4]
  wire  _T_460; // @[MemPrimitives.scala 110:210:@12989.4]
  wire  _T_462; // @[MemPrimitives.scala 110:210:@12990.4]
  wire  _T_463; // @[MemPrimitives.scala 110:228:@12991.4]
  wire  _T_466; // @[MemPrimitives.scala 110:210:@12993.4]
  wire  _T_468; // @[MemPrimitives.scala 110:210:@12994.4]
  wire  _T_469; // @[MemPrimitives.scala 110:228:@12995.4]
  wire  _T_472; // @[MemPrimitives.scala 110:210:@12997.4]
  wire  _T_474; // @[MemPrimitives.scala 110:210:@12998.4]
  wire  _T_475; // @[MemPrimitives.scala 110:228:@12999.4]
  wire  _T_478; // @[MemPrimitives.scala 110:210:@13001.4]
  wire  _T_480; // @[MemPrimitives.scala 110:210:@13002.4]
  wire  _T_481; // @[MemPrimitives.scala 110:228:@13003.4]
  wire  _T_484; // @[MemPrimitives.scala 110:210:@13005.4]
  wire  _T_486; // @[MemPrimitives.scala 110:210:@13006.4]
  wire  _T_487; // @[MemPrimitives.scala 110:228:@13007.4]
  wire  _T_490; // @[MemPrimitives.scala 110:210:@13009.4]
  wire  _T_492; // @[MemPrimitives.scala 110:210:@13010.4]
  wire  _T_493; // @[MemPrimitives.scala 110:228:@13011.4]
  wire  _T_496; // @[MemPrimitives.scala 110:210:@13013.4]
  wire  _T_498; // @[MemPrimitives.scala 110:210:@13014.4]
  wire  _T_499; // @[MemPrimitives.scala 110:228:@13015.4]
  wire  _T_501; // @[MemPrimitives.scala 123:41:@13029.4]
  wire  _T_502; // @[MemPrimitives.scala 123:41:@13030.4]
  wire  _T_503; // @[MemPrimitives.scala 123:41:@13031.4]
  wire  _T_504; // @[MemPrimitives.scala 123:41:@13032.4]
  wire  _T_505; // @[MemPrimitives.scala 123:41:@13033.4]
  wire  _T_506; // @[MemPrimitives.scala 123:41:@13034.4]
  wire  _T_507; // @[MemPrimitives.scala 123:41:@13035.4]
  wire  _T_508; // @[MemPrimitives.scala 123:41:@13036.4]
  wire  _T_509; // @[MemPrimitives.scala 123:41:@13037.4]
  wire [11:0] _T_511; // @[Cat.scala 30:58:@13039.4]
  wire [11:0] _T_513; // @[Cat.scala 30:58:@13041.4]
  wire [11:0] _T_515; // @[Cat.scala 30:58:@13043.4]
  wire [11:0] _T_517; // @[Cat.scala 30:58:@13045.4]
  wire [11:0] _T_519; // @[Cat.scala 30:58:@13047.4]
  wire [11:0] _T_521; // @[Cat.scala 30:58:@13049.4]
  wire [11:0] _T_523; // @[Cat.scala 30:58:@13051.4]
  wire [11:0] _T_525; // @[Cat.scala 30:58:@13053.4]
  wire [11:0] _T_527; // @[Cat.scala 30:58:@13055.4]
  wire [11:0] _T_528; // @[Mux.scala 31:69:@13056.4]
  wire [11:0] _T_529; // @[Mux.scala 31:69:@13057.4]
  wire [11:0] _T_530; // @[Mux.scala 31:69:@13058.4]
  wire [11:0] _T_531; // @[Mux.scala 31:69:@13059.4]
  wire [11:0] _T_532; // @[Mux.scala 31:69:@13060.4]
  wire [11:0] _T_533; // @[Mux.scala 31:69:@13061.4]
  wire [11:0] _T_534; // @[Mux.scala 31:69:@13062.4]
  wire [11:0] _T_535; // @[Mux.scala 31:69:@13063.4]
  wire  _T_542; // @[MemPrimitives.scala 110:210:@13071.4]
  wire  _T_543; // @[MemPrimitives.scala 110:228:@13072.4]
  wire  _T_548; // @[MemPrimitives.scala 110:210:@13075.4]
  wire  _T_549; // @[MemPrimitives.scala 110:228:@13076.4]
  wire  _T_554; // @[MemPrimitives.scala 110:210:@13079.4]
  wire  _T_555; // @[MemPrimitives.scala 110:228:@13080.4]
  wire  _T_560; // @[MemPrimitives.scala 110:210:@13083.4]
  wire  _T_561; // @[MemPrimitives.scala 110:228:@13084.4]
  wire  _T_566; // @[MemPrimitives.scala 110:210:@13087.4]
  wire  _T_567; // @[MemPrimitives.scala 110:228:@13088.4]
  wire  _T_572; // @[MemPrimitives.scala 110:210:@13091.4]
  wire  _T_573; // @[MemPrimitives.scala 110:228:@13092.4]
  wire  _T_578; // @[MemPrimitives.scala 110:210:@13095.4]
  wire  _T_579; // @[MemPrimitives.scala 110:228:@13096.4]
  wire  _T_584; // @[MemPrimitives.scala 110:210:@13099.4]
  wire  _T_585; // @[MemPrimitives.scala 110:228:@13100.4]
  wire  _T_590; // @[MemPrimitives.scala 110:210:@13103.4]
  wire  _T_591; // @[MemPrimitives.scala 110:228:@13104.4]
  wire  _T_593; // @[MemPrimitives.scala 123:41:@13118.4]
  wire  _T_594; // @[MemPrimitives.scala 123:41:@13119.4]
  wire  _T_595; // @[MemPrimitives.scala 123:41:@13120.4]
  wire  _T_596; // @[MemPrimitives.scala 123:41:@13121.4]
  wire  _T_597; // @[MemPrimitives.scala 123:41:@13122.4]
  wire  _T_598; // @[MemPrimitives.scala 123:41:@13123.4]
  wire  _T_599; // @[MemPrimitives.scala 123:41:@13124.4]
  wire  _T_600; // @[MemPrimitives.scala 123:41:@13125.4]
  wire  _T_601; // @[MemPrimitives.scala 123:41:@13126.4]
  wire [11:0] _T_603; // @[Cat.scala 30:58:@13128.4]
  wire [11:0] _T_605; // @[Cat.scala 30:58:@13130.4]
  wire [11:0] _T_607; // @[Cat.scala 30:58:@13132.4]
  wire [11:0] _T_609; // @[Cat.scala 30:58:@13134.4]
  wire [11:0] _T_611; // @[Cat.scala 30:58:@13136.4]
  wire [11:0] _T_613; // @[Cat.scala 30:58:@13138.4]
  wire [11:0] _T_615; // @[Cat.scala 30:58:@13140.4]
  wire [11:0] _T_617; // @[Cat.scala 30:58:@13142.4]
  wire [11:0] _T_619; // @[Cat.scala 30:58:@13144.4]
  wire [11:0] _T_620; // @[Mux.scala 31:69:@13145.4]
  wire [11:0] _T_621; // @[Mux.scala 31:69:@13146.4]
  wire [11:0] _T_622; // @[Mux.scala 31:69:@13147.4]
  wire [11:0] _T_623; // @[Mux.scala 31:69:@13148.4]
  wire [11:0] _T_624; // @[Mux.scala 31:69:@13149.4]
  wire [11:0] _T_625; // @[Mux.scala 31:69:@13150.4]
  wire [11:0] _T_626; // @[Mux.scala 31:69:@13151.4]
  wire [11:0] _T_627; // @[Mux.scala 31:69:@13152.4]
  wire  _T_634; // @[MemPrimitives.scala 110:210:@13160.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@13161.4]
  wire  _T_640; // @[MemPrimitives.scala 110:210:@13164.4]
  wire  _T_641; // @[MemPrimitives.scala 110:228:@13165.4]
  wire  _T_646; // @[MemPrimitives.scala 110:210:@13168.4]
  wire  _T_647; // @[MemPrimitives.scala 110:228:@13169.4]
  wire  _T_652; // @[MemPrimitives.scala 110:210:@13172.4]
  wire  _T_653; // @[MemPrimitives.scala 110:228:@13173.4]
  wire  _T_658; // @[MemPrimitives.scala 110:210:@13176.4]
  wire  _T_659; // @[MemPrimitives.scala 110:228:@13177.4]
  wire  _T_664; // @[MemPrimitives.scala 110:210:@13180.4]
  wire  _T_665; // @[MemPrimitives.scala 110:228:@13181.4]
  wire  _T_670; // @[MemPrimitives.scala 110:210:@13184.4]
  wire  _T_671; // @[MemPrimitives.scala 110:228:@13185.4]
  wire  _T_676; // @[MemPrimitives.scala 110:210:@13188.4]
  wire  _T_677; // @[MemPrimitives.scala 110:228:@13189.4]
  wire  _T_682; // @[MemPrimitives.scala 110:210:@13192.4]
  wire  _T_683; // @[MemPrimitives.scala 110:228:@13193.4]
  wire  _T_685; // @[MemPrimitives.scala 123:41:@13207.4]
  wire  _T_686; // @[MemPrimitives.scala 123:41:@13208.4]
  wire  _T_687; // @[MemPrimitives.scala 123:41:@13209.4]
  wire  _T_688; // @[MemPrimitives.scala 123:41:@13210.4]
  wire  _T_689; // @[MemPrimitives.scala 123:41:@13211.4]
  wire  _T_690; // @[MemPrimitives.scala 123:41:@13212.4]
  wire  _T_691; // @[MemPrimitives.scala 123:41:@13213.4]
  wire  _T_692; // @[MemPrimitives.scala 123:41:@13214.4]
  wire  _T_693; // @[MemPrimitives.scala 123:41:@13215.4]
  wire [11:0] _T_695; // @[Cat.scala 30:58:@13217.4]
  wire [11:0] _T_697; // @[Cat.scala 30:58:@13219.4]
  wire [11:0] _T_699; // @[Cat.scala 30:58:@13221.4]
  wire [11:0] _T_701; // @[Cat.scala 30:58:@13223.4]
  wire [11:0] _T_703; // @[Cat.scala 30:58:@13225.4]
  wire [11:0] _T_705; // @[Cat.scala 30:58:@13227.4]
  wire [11:0] _T_707; // @[Cat.scala 30:58:@13229.4]
  wire [11:0] _T_709; // @[Cat.scala 30:58:@13231.4]
  wire [11:0] _T_711; // @[Cat.scala 30:58:@13233.4]
  wire [11:0] _T_712; // @[Mux.scala 31:69:@13234.4]
  wire [11:0] _T_713; // @[Mux.scala 31:69:@13235.4]
  wire [11:0] _T_714; // @[Mux.scala 31:69:@13236.4]
  wire [11:0] _T_715; // @[Mux.scala 31:69:@13237.4]
  wire [11:0] _T_716; // @[Mux.scala 31:69:@13238.4]
  wire [11:0] _T_717; // @[Mux.scala 31:69:@13239.4]
  wire [11:0] _T_718; // @[Mux.scala 31:69:@13240.4]
  wire [11:0] _T_719; // @[Mux.scala 31:69:@13241.4]
  wire  _T_724; // @[MemPrimitives.scala 110:210:@13248.4]
  wire  _T_727; // @[MemPrimitives.scala 110:228:@13250.4]
  wire  _T_730; // @[MemPrimitives.scala 110:210:@13252.4]
  wire  _T_733; // @[MemPrimitives.scala 110:228:@13254.4]
  wire  _T_736; // @[MemPrimitives.scala 110:210:@13256.4]
  wire  _T_739; // @[MemPrimitives.scala 110:228:@13258.4]
  wire  _T_742; // @[MemPrimitives.scala 110:210:@13260.4]
  wire  _T_745; // @[MemPrimitives.scala 110:228:@13262.4]
  wire  _T_748; // @[MemPrimitives.scala 110:210:@13264.4]
  wire  _T_751; // @[MemPrimitives.scala 110:228:@13266.4]
  wire  _T_754; // @[MemPrimitives.scala 110:210:@13268.4]
  wire  _T_757; // @[MemPrimitives.scala 110:228:@13270.4]
  wire  _T_760; // @[MemPrimitives.scala 110:210:@13272.4]
  wire  _T_763; // @[MemPrimitives.scala 110:228:@13274.4]
  wire  _T_766; // @[MemPrimitives.scala 110:210:@13276.4]
  wire  _T_769; // @[MemPrimitives.scala 110:228:@13278.4]
  wire  _T_772; // @[MemPrimitives.scala 110:210:@13280.4]
  wire  _T_775; // @[MemPrimitives.scala 110:228:@13282.4]
  wire  _T_777; // @[MemPrimitives.scala 123:41:@13296.4]
  wire  _T_778; // @[MemPrimitives.scala 123:41:@13297.4]
  wire  _T_779; // @[MemPrimitives.scala 123:41:@13298.4]
  wire  _T_780; // @[MemPrimitives.scala 123:41:@13299.4]
  wire  _T_781; // @[MemPrimitives.scala 123:41:@13300.4]
  wire  _T_782; // @[MemPrimitives.scala 123:41:@13301.4]
  wire  _T_783; // @[MemPrimitives.scala 123:41:@13302.4]
  wire  _T_784; // @[MemPrimitives.scala 123:41:@13303.4]
  wire  _T_785; // @[MemPrimitives.scala 123:41:@13304.4]
  wire [11:0] _T_787; // @[Cat.scala 30:58:@13306.4]
  wire [11:0] _T_789; // @[Cat.scala 30:58:@13308.4]
  wire [11:0] _T_791; // @[Cat.scala 30:58:@13310.4]
  wire [11:0] _T_793; // @[Cat.scala 30:58:@13312.4]
  wire [11:0] _T_795; // @[Cat.scala 30:58:@13314.4]
  wire [11:0] _T_797; // @[Cat.scala 30:58:@13316.4]
  wire [11:0] _T_799; // @[Cat.scala 30:58:@13318.4]
  wire [11:0] _T_801; // @[Cat.scala 30:58:@13320.4]
  wire [11:0] _T_803; // @[Cat.scala 30:58:@13322.4]
  wire [11:0] _T_804; // @[Mux.scala 31:69:@13323.4]
  wire [11:0] _T_805; // @[Mux.scala 31:69:@13324.4]
  wire [11:0] _T_806; // @[Mux.scala 31:69:@13325.4]
  wire [11:0] _T_807; // @[Mux.scala 31:69:@13326.4]
  wire [11:0] _T_808; // @[Mux.scala 31:69:@13327.4]
  wire [11:0] _T_809; // @[Mux.scala 31:69:@13328.4]
  wire [11:0] _T_810; // @[Mux.scala 31:69:@13329.4]
  wire [11:0] _T_811; // @[Mux.scala 31:69:@13330.4]
  wire  _T_819; // @[MemPrimitives.scala 110:228:@13339.4]
  wire  _T_825; // @[MemPrimitives.scala 110:228:@13343.4]
  wire  _T_831; // @[MemPrimitives.scala 110:228:@13347.4]
  wire  _T_837; // @[MemPrimitives.scala 110:228:@13351.4]
  wire  _T_843; // @[MemPrimitives.scala 110:228:@13355.4]
  wire  _T_849; // @[MemPrimitives.scala 110:228:@13359.4]
  wire  _T_855; // @[MemPrimitives.scala 110:228:@13363.4]
  wire  _T_861; // @[MemPrimitives.scala 110:228:@13367.4]
  wire  _T_867; // @[MemPrimitives.scala 110:228:@13371.4]
  wire  _T_869; // @[MemPrimitives.scala 123:41:@13385.4]
  wire  _T_870; // @[MemPrimitives.scala 123:41:@13386.4]
  wire  _T_871; // @[MemPrimitives.scala 123:41:@13387.4]
  wire  _T_872; // @[MemPrimitives.scala 123:41:@13388.4]
  wire  _T_873; // @[MemPrimitives.scala 123:41:@13389.4]
  wire  _T_874; // @[MemPrimitives.scala 123:41:@13390.4]
  wire  _T_875; // @[MemPrimitives.scala 123:41:@13391.4]
  wire  _T_876; // @[MemPrimitives.scala 123:41:@13392.4]
  wire  _T_877; // @[MemPrimitives.scala 123:41:@13393.4]
  wire [11:0] _T_879; // @[Cat.scala 30:58:@13395.4]
  wire [11:0] _T_881; // @[Cat.scala 30:58:@13397.4]
  wire [11:0] _T_883; // @[Cat.scala 30:58:@13399.4]
  wire [11:0] _T_885; // @[Cat.scala 30:58:@13401.4]
  wire [11:0] _T_887; // @[Cat.scala 30:58:@13403.4]
  wire [11:0] _T_889; // @[Cat.scala 30:58:@13405.4]
  wire [11:0] _T_891; // @[Cat.scala 30:58:@13407.4]
  wire [11:0] _T_893; // @[Cat.scala 30:58:@13409.4]
  wire [11:0] _T_895; // @[Cat.scala 30:58:@13411.4]
  wire [11:0] _T_896; // @[Mux.scala 31:69:@13412.4]
  wire [11:0] _T_897; // @[Mux.scala 31:69:@13413.4]
  wire [11:0] _T_898; // @[Mux.scala 31:69:@13414.4]
  wire [11:0] _T_899; // @[Mux.scala 31:69:@13415.4]
  wire [11:0] _T_900; // @[Mux.scala 31:69:@13416.4]
  wire [11:0] _T_901; // @[Mux.scala 31:69:@13417.4]
  wire [11:0] _T_902; // @[Mux.scala 31:69:@13418.4]
  wire [11:0] _T_903; // @[Mux.scala 31:69:@13419.4]
  wire  _T_911; // @[MemPrimitives.scala 110:228:@13428.4]
  wire  _T_917; // @[MemPrimitives.scala 110:228:@13432.4]
  wire  _T_923; // @[MemPrimitives.scala 110:228:@13436.4]
  wire  _T_929; // @[MemPrimitives.scala 110:228:@13440.4]
  wire  _T_935; // @[MemPrimitives.scala 110:228:@13444.4]
  wire  _T_941; // @[MemPrimitives.scala 110:228:@13448.4]
  wire  _T_947; // @[MemPrimitives.scala 110:228:@13452.4]
  wire  _T_953; // @[MemPrimitives.scala 110:228:@13456.4]
  wire  _T_959; // @[MemPrimitives.scala 110:228:@13460.4]
  wire  _T_961; // @[MemPrimitives.scala 123:41:@13474.4]
  wire  _T_962; // @[MemPrimitives.scala 123:41:@13475.4]
  wire  _T_963; // @[MemPrimitives.scala 123:41:@13476.4]
  wire  _T_964; // @[MemPrimitives.scala 123:41:@13477.4]
  wire  _T_965; // @[MemPrimitives.scala 123:41:@13478.4]
  wire  _T_966; // @[MemPrimitives.scala 123:41:@13479.4]
  wire  _T_967; // @[MemPrimitives.scala 123:41:@13480.4]
  wire  _T_968; // @[MemPrimitives.scala 123:41:@13481.4]
  wire  _T_969; // @[MemPrimitives.scala 123:41:@13482.4]
  wire [11:0] _T_971; // @[Cat.scala 30:58:@13484.4]
  wire [11:0] _T_973; // @[Cat.scala 30:58:@13486.4]
  wire [11:0] _T_975; // @[Cat.scala 30:58:@13488.4]
  wire [11:0] _T_977; // @[Cat.scala 30:58:@13490.4]
  wire [11:0] _T_979; // @[Cat.scala 30:58:@13492.4]
  wire [11:0] _T_981; // @[Cat.scala 30:58:@13494.4]
  wire [11:0] _T_983; // @[Cat.scala 30:58:@13496.4]
  wire [11:0] _T_985; // @[Cat.scala 30:58:@13498.4]
  wire [11:0] _T_987; // @[Cat.scala 30:58:@13500.4]
  wire [11:0] _T_988; // @[Mux.scala 31:69:@13501.4]
  wire [11:0] _T_989; // @[Mux.scala 31:69:@13502.4]
  wire [11:0] _T_990; // @[Mux.scala 31:69:@13503.4]
  wire [11:0] _T_991; // @[Mux.scala 31:69:@13504.4]
  wire [11:0] _T_992; // @[Mux.scala 31:69:@13505.4]
  wire [11:0] _T_993; // @[Mux.scala 31:69:@13506.4]
  wire [11:0] _T_994; // @[Mux.scala 31:69:@13507.4]
  wire [11:0] _T_995; // @[Mux.scala 31:69:@13508.4]
  wire  _T_1000; // @[MemPrimitives.scala 110:210:@13515.4]
  wire  _T_1003; // @[MemPrimitives.scala 110:228:@13517.4]
  wire  _T_1006; // @[MemPrimitives.scala 110:210:@13519.4]
  wire  _T_1009; // @[MemPrimitives.scala 110:228:@13521.4]
  wire  _T_1012; // @[MemPrimitives.scala 110:210:@13523.4]
  wire  _T_1015; // @[MemPrimitives.scala 110:228:@13525.4]
  wire  _T_1018; // @[MemPrimitives.scala 110:210:@13527.4]
  wire  _T_1021; // @[MemPrimitives.scala 110:228:@13529.4]
  wire  _T_1024; // @[MemPrimitives.scala 110:210:@13531.4]
  wire  _T_1027; // @[MemPrimitives.scala 110:228:@13533.4]
  wire  _T_1030; // @[MemPrimitives.scala 110:210:@13535.4]
  wire  _T_1033; // @[MemPrimitives.scala 110:228:@13537.4]
  wire  _T_1036; // @[MemPrimitives.scala 110:210:@13539.4]
  wire  _T_1039; // @[MemPrimitives.scala 110:228:@13541.4]
  wire  _T_1042; // @[MemPrimitives.scala 110:210:@13543.4]
  wire  _T_1045; // @[MemPrimitives.scala 110:228:@13545.4]
  wire  _T_1048; // @[MemPrimitives.scala 110:210:@13547.4]
  wire  _T_1051; // @[MemPrimitives.scala 110:228:@13549.4]
  wire  _T_1053; // @[MemPrimitives.scala 123:41:@13563.4]
  wire  _T_1054; // @[MemPrimitives.scala 123:41:@13564.4]
  wire  _T_1055; // @[MemPrimitives.scala 123:41:@13565.4]
  wire  _T_1056; // @[MemPrimitives.scala 123:41:@13566.4]
  wire  _T_1057; // @[MemPrimitives.scala 123:41:@13567.4]
  wire  _T_1058; // @[MemPrimitives.scala 123:41:@13568.4]
  wire  _T_1059; // @[MemPrimitives.scala 123:41:@13569.4]
  wire  _T_1060; // @[MemPrimitives.scala 123:41:@13570.4]
  wire  _T_1061; // @[MemPrimitives.scala 123:41:@13571.4]
  wire [11:0] _T_1063; // @[Cat.scala 30:58:@13573.4]
  wire [11:0] _T_1065; // @[Cat.scala 30:58:@13575.4]
  wire [11:0] _T_1067; // @[Cat.scala 30:58:@13577.4]
  wire [11:0] _T_1069; // @[Cat.scala 30:58:@13579.4]
  wire [11:0] _T_1071; // @[Cat.scala 30:58:@13581.4]
  wire [11:0] _T_1073; // @[Cat.scala 30:58:@13583.4]
  wire [11:0] _T_1075; // @[Cat.scala 30:58:@13585.4]
  wire [11:0] _T_1077; // @[Cat.scala 30:58:@13587.4]
  wire [11:0] _T_1079; // @[Cat.scala 30:58:@13589.4]
  wire [11:0] _T_1080; // @[Mux.scala 31:69:@13590.4]
  wire [11:0] _T_1081; // @[Mux.scala 31:69:@13591.4]
  wire [11:0] _T_1082; // @[Mux.scala 31:69:@13592.4]
  wire [11:0] _T_1083; // @[Mux.scala 31:69:@13593.4]
  wire [11:0] _T_1084; // @[Mux.scala 31:69:@13594.4]
  wire [11:0] _T_1085; // @[Mux.scala 31:69:@13595.4]
  wire [11:0] _T_1086; // @[Mux.scala 31:69:@13596.4]
  wire [11:0] _T_1087; // @[Mux.scala 31:69:@13597.4]
  wire  _T_1095; // @[MemPrimitives.scala 110:228:@13606.4]
  wire  _T_1101; // @[MemPrimitives.scala 110:228:@13610.4]
  wire  _T_1107; // @[MemPrimitives.scala 110:228:@13614.4]
  wire  _T_1113; // @[MemPrimitives.scala 110:228:@13618.4]
  wire  _T_1119; // @[MemPrimitives.scala 110:228:@13622.4]
  wire  _T_1125; // @[MemPrimitives.scala 110:228:@13626.4]
  wire  _T_1131; // @[MemPrimitives.scala 110:228:@13630.4]
  wire  _T_1137; // @[MemPrimitives.scala 110:228:@13634.4]
  wire  _T_1143; // @[MemPrimitives.scala 110:228:@13638.4]
  wire  _T_1145; // @[MemPrimitives.scala 123:41:@13652.4]
  wire  _T_1146; // @[MemPrimitives.scala 123:41:@13653.4]
  wire  _T_1147; // @[MemPrimitives.scala 123:41:@13654.4]
  wire  _T_1148; // @[MemPrimitives.scala 123:41:@13655.4]
  wire  _T_1149; // @[MemPrimitives.scala 123:41:@13656.4]
  wire  _T_1150; // @[MemPrimitives.scala 123:41:@13657.4]
  wire  _T_1151; // @[MemPrimitives.scala 123:41:@13658.4]
  wire  _T_1152; // @[MemPrimitives.scala 123:41:@13659.4]
  wire  _T_1153; // @[MemPrimitives.scala 123:41:@13660.4]
  wire [11:0] _T_1155; // @[Cat.scala 30:58:@13662.4]
  wire [11:0] _T_1157; // @[Cat.scala 30:58:@13664.4]
  wire [11:0] _T_1159; // @[Cat.scala 30:58:@13666.4]
  wire [11:0] _T_1161; // @[Cat.scala 30:58:@13668.4]
  wire [11:0] _T_1163; // @[Cat.scala 30:58:@13670.4]
  wire [11:0] _T_1165; // @[Cat.scala 30:58:@13672.4]
  wire [11:0] _T_1167; // @[Cat.scala 30:58:@13674.4]
  wire [11:0] _T_1169; // @[Cat.scala 30:58:@13676.4]
  wire [11:0] _T_1171; // @[Cat.scala 30:58:@13678.4]
  wire [11:0] _T_1172; // @[Mux.scala 31:69:@13679.4]
  wire [11:0] _T_1173; // @[Mux.scala 31:69:@13680.4]
  wire [11:0] _T_1174; // @[Mux.scala 31:69:@13681.4]
  wire [11:0] _T_1175; // @[Mux.scala 31:69:@13682.4]
  wire [11:0] _T_1176; // @[Mux.scala 31:69:@13683.4]
  wire [11:0] _T_1177; // @[Mux.scala 31:69:@13684.4]
  wire [11:0] _T_1178; // @[Mux.scala 31:69:@13685.4]
  wire [11:0] _T_1179; // @[Mux.scala 31:69:@13686.4]
  wire  _T_1187; // @[MemPrimitives.scala 110:228:@13695.4]
  wire  _T_1193; // @[MemPrimitives.scala 110:228:@13699.4]
  wire  _T_1199; // @[MemPrimitives.scala 110:228:@13703.4]
  wire  _T_1205; // @[MemPrimitives.scala 110:228:@13707.4]
  wire  _T_1211; // @[MemPrimitives.scala 110:228:@13711.4]
  wire  _T_1217; // @[MemPrimitives.scala 110:228:@13715.4]
  wire  _T_1223; // @[MemPrimitives.scala 110:228:@13719.4]
  wire  _T_1229; // @[MemPrimitives.scala 110:228:@13723.4]
  wire  _T_1235; // @[MemPrimitives.scala 110:228:@13727.4]
  wire  _T_1237; // @[MemPrimitives.scala 123:41:@13741.4]
  wire  _T_1238; // @[MemPrimitives.scala 123:41:@13742.4]
  wire  _T_1239; // @[MemPrimitives.scala 123:41:@13743.4]
  wire  _T_1240; // @[MemPrimitives.scala 123:41:@13744.4]
  wire  _T_1241; // @[MemPrimitives.scala 123:41:@13745.4]
  wire  _T_1242; // @[MemPrimitives.scala 123:41:@13746.4]
  wire  _T_1243; // @[MemPrimitives.scala 123:41:@13747.4]
  wire  _T_1244; // @[MemPrimitives.scala 123:41:@13748.4]
  wire  _T_1245; // @[MemPrimitives.scala 123:41:@13749.4]
  wire [11:0] _T_1247; // @[Cat.scala 30:58:@13751.4]
  wire [11:0] _T_1249; // @[Cat.scala 30:58:@13753.4]
  wire [11:0] _T_1251; // @[Cat.scala 30:58:@13755.4]
  wire [11:0] _T_1253; // @[Cat.scala 30:58:@13757.4]
  wire [11:0] _T_1255; // @[Cat.scala 30:58:@13759.4]
  wire [11:0] _T_1257; // @[Cat.scala 30:58:@13761.4]
  wire [11:0] _T_1259; // @[Cat.scala 30:58:@13763.4]
  wire [11:0] _T_1261; // @[Cat.scala 30:58:@13765.4]
  wire [11:0] _T_1263; // @[Cat.scala 30:58:@13767.4]
  wire [11:0] _T_1264; // @[Mux.scala 31:69:@13768.4]
  wire [11:0] _T_1265; // @[Mux.scala 31:69:@13769.4]
  wire [11:0] _T_1266; // @[Mux.scala 31:69:@13770.4]
  wire [11:0] _T_1267; // @[Mux.scala 31:69:@13771.4]
  wire [11:0] _T_1268; // @[Mux.scala 31:69:@13772.4]
  wire [11:0] _T_1269; // @[Mux.scala 31:69:@13773.4]
  wire [11:0] _T_1270; // @[Mux.scala 31:69:@13774.4]
  wire [11:0] _T_1271; // @[Mux.scala 31:69:@13775.4]
  wire  _T_1276; // @[MemPrimitives.scala 110:210:@13782.4]
  wire  _T_1279; // @[MemPrimitives.scala 110:228:@13784.4]
  wire  _T_1282; // @[MemPrimitives.scala 110:210:@13786.4]
  wire  _T_1285; // @[MemPrimitives.scala 110:228:@13788.4]
  wire  _T_1288; // @[MemPrimitives.scala 110:210:@13790.4]
  wire  _T_1291; // @[MemPrimitives.scala 110:228:@13792.4]
  wire  _T_1294; // @[MemPrimitives.scala 110:210:@13794.4]
  wire  _T_1297; // @[MemPrimitives.scala 110:228:@13796.4]
  wire  _T_1300; // @[MemPrimitives.scala 110:210:@13798.4]
  wire  _T_1303; // @[MemPrimitives.scala 110:228:@13800.4]
  wire  _T_1306; // @[MemPrimitives.scala 110:210:@13802.4]
  wire  _T_1309; // @[MemPrimitives.scala 110:228:@13804.4]
  wire  _T_1312; // @[MemPrimitives.scala 110:210:@13806.4]
  wire  _T_1315; // @[MemPrimitives.scala 110:228:@13808.4]
  wire  _T_1318; // @[MemPrimitives.scala 110:210:@13810.4]
  wire  _T_1321; // @[MemPrimitives.scala 110:228:@13812.4]
  wire  _T_1324; // @[MemPrimitives.scala 110:210:@13814.4]
  wire  _T_1327; // @[MemPrimitives.scala 110:228:@13816.4]
  wire  _T_1329; // @[MemPrimitives.scala 123:41:@13830.4]
  wire  _T_1330; // @[MemPrimitives.scala 123:41:@13831.4]
  wire  _T_1331; // @[MemPrimitives.scala 123:41:@13832.4]
  wire  _T_1332; // @[MemPrimitives.scala 123:41:@13833.4]
  wire  _T_1333; // @[MemPrimitives.scala 123:41:@13834.4]
  wire  _T_1334; // @[MemPrimitives.scala 123:41:@13835.4]
  wire  _T_1335; // @[MemPrimitives.scala 123:41:@13836.4]
  wire  _T_1336; // @[MemPrimitives.scala 123:41:@13837.4]
  wire  _T_1337; // @[MemPrimitives.scala 123:41:@13838.4]
  wire [11:0] _T_1339; // @[Cat.scala 30:58:@13840.4]
  wire [11:0] _T_1341; // @[Cat.scala 30:58:@13842.4]
  wire [11:0] _T_1343; // @[Cat.scala 30:58:@13844.4]
  wire [11:0] _T_1345; // @[Cat.scala 30:58:@13846.4]
  wire [11:0] _T_1347; // @[Cat.scala 30:58:@13848.4]
  wire [11:0] _T_1349; // @[Cat.scala 30:58:@13850.4]
  wire [11:0] _T_1351; // @[Cat.scala 30:58:@13852.4]
  wire [11:0] _T_1353; // @[Cat.scala 30:58:@13854.4]
  wire [11:0] _T_1355; // @[Cat.scala 30:58:@13856.4]
  wire [11:0] _T_1356; // @[Mux.scala 31:69:@13857.4]
  wire [11:0] _T_1357; // @[Mux.scala 31:69:@13858.4]
  wire [11:0] _T_1358; // @[Mux.scala 31:69:@13859.4]
  wire [11:0] _T_1359; // @[Mux.scala 31:69:@13860.4]
  wire [11:0] _T_1360; // @[Mux.scala 31:69:@13861.4]
  wire [11:0] _T_1361; // @[Mux.scala 31:69:@13862.4]
  wire [11:0] _T_1362; // @[Mux.scala 31:69:@13863.4]
  wire [11:0] _T_1363; // @[Mux.scala 31:69:@13864.4]
  wire  _T_1371; // @[MemPrimitives.scala 110:228:@13873.4]
  wire  _T_1377; // @[MemPrimitives.scala 110:228:@13877.4]
  wire  _T_1383; // @[MemPrimitives.scala 110:228:@13881.4]
  wire  _T_1389; // @[MemPrimitives.scala 110:228:@13885.4]
  wire  _T_1395; // @[MemPrimitives.scala 110:228:@13889.4]
  wire  _T_1401; // @[MemPrimitives.scala 110:228:@13893.4]
  wire  _T_1407; // @[MemPrimitives.scala 110:228:@13897.4]
  wire  _T_1413; // @[MemPrimitives.scala 110:228:@13901.4]
  wire  _T_1419; // @[MemPrimitives.scala 110:228:@13905.4]
  wire  _T_1421; // @[MemPrimitives.scala 123:41:@13919.4]
  wire  _T_1422; // @[MemPrimitives.scala 123:41:@13920.4]
  wire  _T_1423; // @[MemPrimitives.scala 123:41:@13921.4]
  wire  _T_1424; // @[MemPrimitives.scala 123:41:@13922.4]
  wire  _T_1425; // @[MemPrimitives.scala 123:41:@13923.4]
  wire  _T_1426; // @[MemPrimitives.scala 123:41:@13924.4]
  wire  _T_1427; // @[MemPrimitives.scala 123:41:@13925.4]
  wire  _T_1428; // @[MemPrimitives.scala 123:41:@13926.4]
  wire  _T_1429; // @[MemPrimitives.scala 123:41:@13927.4]
  wire [11:0] _T_1431; // @[Cat.scala 30:58:@13929.4]
  wire [11:0] _T_1433; // @[Cat.scala 30:58:@13931.4]
  wire [11:0] _T_1435; // @[Cat.scala 30:58:@13933.4]
  wire [11:0] _T_1437; // @[Cat.scala 30:58:@13935.4]
  wire [11:0] _T_1439; // @[Cat.scala 30:58:@13937.4]
  wire [11:0] _T_1441; // @[Cat.scala 30:58:@13939.4]
  wire [11:0] _T_1443; // @[Cat.scala 30:58:@13941.4]
  wire [11:0] _T_1445; // @[Cat.scala 30:58:@13943.4]
  wire [11:0] _T_1447; // @[Cat.scala 30:58:@13945.4]
  wire [11:0] _T_1448; // @[Mux.scala 31:69:@13946.4]
  wire [11:0] _T_1449; // @[Mux.scala 31:69:@13947.4]
  wire [11:0] _T_1450; // @[Mux.scala 31:69:@13948.4]
  wire [11:0] _T_1451; // @[Mux.scala 31:69:@13949.4]
  wire [11:0] _T_1452; // @[Mux.scala 31:69:@13950.4]
  wire [11:0] _T_1453; // @[Mux.scala 31:69:@13951.4]
  wire [11:0] _T_1454; // @[Mux.scala 31:69:@13952.4]
  wire [11:0] _T_1455; // @[Mux.scala 31:69:@13953.4]
  wire  _T_1463; // @[MemPrimitives.scala 110:228:@13962.4]
  wire  _T_1469; // @[MemPrimitives.scala 110:228:@13966.4]
  wire  _T_1475; // @[MemPrimitives.scala 110:228:@13970.4]
  wire  _T_1481; // @[MemPrimitives.scala 110:228:@13974.4]
  wire  _T_1487; // @[MemPrimitives.scala 110:228:@13978.4]
  wire  _T_1493; // @[MemPrimitives.scala 110:228:@13982.4]
  wire  _T_1499; // @[MemPrimitives.scala 110:228:@13986.4]
  wire  _T_1505; // @[MemPrimitives.scala 110:228:@13990.4]
  wire  _T_1511; // @[MemPrimitives.scala 110:228:@13994.4]
  wire  _T_1513; // @[MemPrimitives.scala 123:41:@14008.4]
  wire  _T_1514; // @[MemPrimitives.scala 123:41:@14009.4]
  wire  _T_1515; // @[MemPrimitives.scala 123:41:@14010.4]
  wire  _T_1516; // @[MemPrimitives.scala 123:41:@14011.4]
  wire  _T_1517; // @[MemPrimitives.scala 123:41:@14012.4]
  wire  _T_1518; // @[MemPrimitives.scala 123:41:@14013.4]
  wire  _T_1519; // @[MemPrimitives.scala 123:41:@14014.4]
  wire  _T_1520; // @[MemPrimitives.scala 123:41:@14015.4]
  wire  _T_1521; // @[MemPrimitives.scala 123:41:@14016.4]
  wire [11:0] _T_1523; // @[Cat.scala 30:58:@14018.4]
  wire [11:0] _T_1525; // @[Cat.scala 30:58:@14020.4]
  wire [11:0] _T_1527; // @[Cat.scala 30:58:@14022.4]
  wire [11:0] _T_1529; // @[Cat.scala 30:58:@14024.4]
  wire [11:0] _T_1531; // @[Cat.scala 30:58:@14026.4]
  wire [11:0] _T_1533; // @[Cat.scala 30:58:@14028.4]
  wire [11:0] _T_1535; // @[Cat.scala 30:58:@14030.4]
  wire [11:0] _T_1537; // @[Cat.scala 30:58:@14032.4]
  wire [11:0] _T_1539; // @[Cat.scala 30:58:@14034.4]
  wire [11:0] _T_1540; // @[Mux.scala 31:69:@14035.4]
  wire [11:0] _T_1541; // @[Mux.scala 31:69:@14036.4]
  wire [11:0] _T_1542; // @[Mux.scala 31:69:@14037.4]
  wire [11:0] _T_1543; // @[Mux.scala 31:69:@14038.4]
  wire [11:0] _T_1544; // @[Mux.scala 31:69:@14039.4]
  wire [11:0] _T_1545; // @[Mux.scala 31:69:@14040.4]
  wire [11:0] _T_1546; // @[Mux.scala 31:69:@14041.4]
  wire [11:0] _T_1547; // @[Mux.scala 31:69:@14042.4]
  wire  _T_1643; // @[package.scala 96:25:@14171.4 package.scala 96:25:@14172.4]
  wire [7:0] _T_1647; // @[Mux.scala 31:69:@14181.4]
  wire  _T_1640; // @[package.scala 96:25:@14163.4 package.scala 96:25:@14164.4]
  wire [7:0] _T_1648; // @[Mux.scala 31:69:@14182.4]
  wire  _T_1637; // @[package.scala 96:25:@14155.4 package.scala 96:25:@14156.4]
  wire [7:0] _T_1649; // @[Mux.scala 31:69:@14183.4]
  wire  _T_1634; // @[package.scala 96:25:@14147.4 package.scala 96:25:@14148.4]
  wire [7:0] _T_1650; // @[Mux.scala 31:69:@14184.4]
  wire  _T_1631; // @[package.scala 96:25:@14139.4 package.scala 96:25:@14140.4]
  wire [7:0] _T_1651; // @[Mux.scala 31:69:@14185.4]
  wire  _T_1628; // @[package.scala 96:25:@14131.4 package.scala 96:25:@14132.4]
  wire [7:0] _T_1652; // @[Mux.scala 31:69:@14186.4]
  wire  _T_1625; // @[package.scala 96:25:@14123.4 package.scala 96:25:@14124.4]
  wire [7:0] _T_1653; // @[Mux.scala 31:69:@14187.4]
  wire  _T_1622; // @[package.scala 96:25:@14115.4 package.scala 96:25:@14116.4]
  wire [7:0] _T_1654; // @[Mux.scala 31:69:@14188.4]
  wire  _T_1619; // @[package.scala 96:25:@14107.4 package.scala 96:25:@14108.4]
  wire [7:0] _T_1655; // @[Mux.scala 31:69:@14189.4]
  wire  _T_1616; // @[package.scala 96:25:@14099.4 package.scala 96:25:@14100.4]
  wire [7:0] _T_1656; // @[Mux.scala 31:69:@14190.4]
  wire  _T_1613; // @[package.scala 96:25:@14091.4 package.scala 96:25:@14092.4]
  wire  _T_1750; // @[package.scala 96:25:@14315.4 package.scala 96:25:@14316.4]
  wire [7:0] _T_1754; // @[Mux.scala 31:69:@14325.4]
  wire  _T_1747; // @[package.scala 96:25:@14307.4 package.scala 96:25:@14308.4]
  wire [7:0] _T_1755; // @[Mux.scala 31:69:@14326.4]
  wire  _T_1744; // @[package.scala 96:25:@14299.4 package.scala 96:25:@14300.4]
  wire [7:0] _T_1756; // @[Mux.scala 31:69:@14327.4]
  wire  _T_1741; // @[package.scala 96:25:@14291.4 package.scala 96:25:@14292.4]
  wire [7:0] _T_1757; // @[Mux.scala 31:69:@14328.4]
  wire  _T_1738; // @[package.scala 96:25:@14283.4 package.scala 96:25:@14284.4]
  wire [7:0] _T_1758; // @[Mux.scala 31:69:@14329.4]
  wire  _T_1735; // @[package.scala 96:25:@14275.4 package.scala 96:25:@14276.4]
  wire [7:0] _T_1759; // @[Mux.scala 31:69:@14330.4]
  wire  _T_1732; // @[package.scala 96:25:@14267.4 package.scala 96:25:@14268.4]
  wire [7:0] _T_1760; // @[Mux.scala 31:69:@14331.4]
  wire  _T_1729; // @[package.scala 96:25:@14259.4 package.scala 96:25:@14260.4]
  wire [7:0] _T_1761; // @[Mux.scala 31:69:@14332.4]
  wire  _T_1726; // @[package.scala 96:25:@14251.4 package.scala 96:25:@14252.4]
  wire [7:0] _T_1762; // @[Mux.scala 31:69:@14333.4]
  wire  _T_1723; // @[package.scala 96:25:@14243.4 package.scala 96:25:@14244.4]
  wire [7:0] _T_1763; // @[Mux.scala 31:69:@14334.4]
  wire  _T_1720; // @[package.scala 96:25:@14235.4 package.scala 96:25:@14236.4]
  wire  _T_1857; // @[package.scala 96:25:@14459.4 package.scala 96:25:@14460.4]
  wire [7:0] _T_1861; // @[Mux.scala 31:69:@14469.4]
  wire  _T_1854; // @[package.scala 96:25:@14451.4 package.scala 96:25:@14452.4]
  wire [7:0] _T_1862; // @[Mux.scala 31:69:@14470.4]
  wire  _T_1851; // @[package.scala 96:25:@14443.4 package.scala 96:25:@14444.4]
  wire [7:0] _T_1863; // @[Mux.scala 31:69:@14471.4]
  wire  _T_1848; // @[package.scala 96:25:@14435.4 package.scala 96:25:@14436.4]
  wire [7:0] _T_1864; // @[Mux.scala 31:69:@14472.4]
  wire  _T_1845; // @[package.scala 96:25:@14427.4 package.scala 96:25:@14428.4]
  wire [7:0] _T_1865; // @[Mux.scala 31:69:@14473.4]
  wire  _T_1842; // @[package.scala 96:25:@14419.4 package.scala 96:25:@14420.4]
  wire [7:0] _T_1866; // @[Mux.scala 31:69:@14474.4]
  wire  _T_1839; // @[package.scala 96:25:@14411.4 package.scala 96:25:@14412.4]
  wire [7:0] _T_1867; // @[Mux.scala 31:69:@14475.4]
  wire  _T_1836; // @[package.scala 96:25:@14403.4 package.scala 96:25:@14404.4]
  wire [7:0] _T_1868; // @[Mux.scala 31:69:@14476.4]
  wire  _T_1833; // @[package.scala 96:25:@14395.4 package.scala 96:25:@14396.4]
  wire [7:0] _T_1869; // @[Mux.scala 31:69:@14477.4]
  wire  _T_1830; // @[package.scala 96:25:@14387.4 package.scala 96:25:@14388.4]
  wire [7:0] _T_1870; // @[Mux.scala 31:69:@14478.4]
  wire  _T_1827; // @[package.scala 96:25:@14379.4 package.scala 96:25:@14380.4]
  wire  _T_1964; // @[package.scala 96:25:@14603.4 package.scala 96:25:@14604.4]
  wire [7:0] _T_1968; // @[Mux.scala 31:69:@14613.4]
  wire  _T_1961; // @[package.scala 96:25:@14595.4 package.scala 96:25:@14596.4]
  wire [7:0] _T_1969; // @[Mux.scala 31:69:@14614.4]
  wire  _T_1958; // @[package.scala 96:25:@14587.4 package.scala 96:25:@14588.4]
  wire [7:0] _T_1970; // @[Mux.scala 31:69:@14615.4]
  wire  _T_1955; // @[package.scala 96:25:@14579.4 package.scala 96:25:@14580.4]
  wire [7:0] _T_1971; // @[Mux.scala 31:69:@14616.4]
  wire  _T_1952; // @[package.scala 96:25:@14571.4 package.scala 96:25:@14572.4]
  wire [7:0] _T_1972; // @[Mux.scala 31:69:@14617.4]
  wire  _T_1949; // @[package.scala 96:25:@14563.4 package.scala 96:25:@14564.4]
  wire [7:0] _T_1973; // @[Mux.scala 31:69:@14618.4]
  wire  _T_1946; // @[package.scala 96:25:@14555.4 package.scala 96:25:@14556.4]
  wire [7:0] _T_1974; // @[Mux.scala 31:69:@14619.4]
  wire  _T_1943; // @[package.scala 96:25:@14547.4 package.scala 96:25:@14548.4]
  wire [7:0] _T_1975; // @[Mux.scala 31:69:@14620.4]
  wire  _T_1940; // @[package.scala 96:25:@14539.4 package.scala 96:25:@14540.4]
  wire [7:0] _T_1976; // @[Mux.scala 31:69:@14621.4]
  wire  _T_1937; // @[package.scala 96:25:@14531.4 package.scala 96:25:@14532.4]
  wire [7:0] _T_1977; // @[Mux.scala 31:69:@14622.4]
  wire  _T_1934; // @[package.scala 96:25:@14523.4 package.scala 96:25:@14524.4]
  wire  _T_2071; // @[package.scala 96:25:@14747.4 package.scala 96:25:@14748.4]
  wire [7:0] _T_2075; // @[Mux.scala 31:69:@14757.4]
  wire  _T_2068; // @[package.scala 96:25:@14739.4 package.scala 96:25:@14740.4]
  wire [7:0] _T_2076; // @[Mux.scala 31:69:@14758.4]
  wire  _T_2065; // @[package.scala 96:25:@14731.4 package.scala 96:25:@14732.4]
  wire [7:0] _T_2077; // @[Mux.scala 31:69:@14759.4]
  wire  _T_2062; // @[package.scala 96:25:@14723.4 package.scala 96:25:@14724.4]
  wire [7:0] _T_2078; // @[Mux.scala 31:69:@14760.4]
  wire  _T_2059; // @[package.scala 96:25:@14715.4 package.scala 96:25:@14716.4]
  wire [7:0] _T_2079; // @[Mux.scala 31:69:@14761.4]
  wire  _T_2056; // @[package.scala 96:25:@14707.4 package.scala 96:25:@14708.4]
  wire [7:0] _T_2080; // @[Mux.scala 31:69:@14762.4]
  wire  _T_2053; // @[package.scala 96:25:@14699.4 package.scala 96:25:@14700.4]
  wire [7:0] _T_2081; // @[Mux.scala 31:69:@14763.4]
  wire  _T_2050; // @[package.scala 96:25:@14691.4 package.scala 96:25:@14692.4]
  wire [7:0] _T_2082; // @[Mux.scala 31:69:@14764.4]
  wire  _T_2047; // @[package.scala 96:25:@14683.4 package.scala 96:25:@14684.4]
  wire [7:0] _T_2083; // @[Mux.scala 31:69:@14765.4]
  wire  _T_2044; // @[package.scala 96:25:@14675.4 package.scala 96:25:@14676.4]
  wire [7:0] _T_2084; // @[Mux.scala 31:69:@14766.4]
  wire  _T_2041; // @[package.scala 96:25:@14667.4 package.scala 96:25:@14668.4]
  wire  _T_2178; // @[package.scala 96:25:@14891.4 package.scala 96:25:@14892.4]
  wire [7:0] _T_2182; // @[Mux.scala 31:69:@14901.4]
  wire  _T_2175; // @[package.scala 96:25:@14883.4 package.scala 96:25:@14884.4]
  wire [7:0] _T_2183; // @[Mux.scala 31:69:@14902.4]
  wire  _T_2172; // @[package.scala 96:25:@14875.4 package.scala 96:25:@14876.4]
  wire [7:0] _T_2184; // @[Mux.scala 31:69:@14903.4]
  wire  _T_2169; // @[package.scala 96:25:@14867.4 package.scala 96:25:@14868.4]
  wire [7:0] _T_2185; // @[Mux.scala 31:69:@14904.4]
  wire  _T_2166; // @[package.scala 96:25:@14859.4 package.scala 96:25:@14860.4]
  wire [7:0] _T_2186; // @[Mux.scala 31:69:@14905.4]
  wire  _T_2163; // @[package.scala 96:25:@14851.4 package.scala 96:25:@14852.4]
  wire [7:0] _T_2187; // @[Mux.scala 31:69:@14906.4]
  wire  _T_2160; // @[package.scala 96:25:@14843.4 package.scala 96:25:@14844.4]
  wire [7:0] _T_2188; // @[Mux.scala 31:69:@14907.4]
  wire  _T_2157; // @[package.scala 96:25:@14835.4 package.scala 96:25:@14836.4]
  wire [7:0] _T_2189; // @[Mux.scala 31:69:@14908.4]
  wire  _T_2154; // @[package.scala 96:25:@14827.4 package.scala 96:25:@14828.4]
  wire [7:0] _T_2190; // @[Mux.scala 31:69:@14909.4]
  wire  _T_2151; // @[package.scala 96:25:@14819.4 package.scala 96:25:@14820.4]
  wire [7:0] _T_2191; // @[Mux.scala 31:69:@14910.4]
  wire  _T_2148; // @[package.scala 96:25:@14811.4 package.scala 96:25:@14812.4]
  wire  _T_2285; // @[package.scala 96:25:@15035.4 package.scala 96:25:@15036.4]
  wire [7:0] _T_2289; // @[Mux.scala 31:69:@15045.4]
  wire  _T_2282; // @[package.scala 96:25:@15027.4 package.scala 96:25:@15028.4]
  wire [7:0] _T_2290; // @[Mux.scala 31:69:@15046.4]
  wire  _T_2279; // @[package.scala 96:25:@15019.4 package.scala 96:25:@15020.4]
  wire [7:0] _T_2291; // @[Mux.scala 31:69:@15047.4]
  wire  _T_2276; // @[package.scala 96:25:@15011.4 package.scala 96:25:@15012.4]
  wire [7:0] _T_2292; // @[Mux.scala 31:69:@15048.4]
  wire  _T_2273; // @[package.scala 96:25:@15003.4 package.scala 96:25:@15004.4]
  wire [7:0] _T_2293; // @[Mux.scala 31:69:@15049.4]
  wire  _T_2270; // @[package.scala 96:25:@14995.4 package.scala 96:25:@14996.4]
  wire [7:0] _T_2294; // @[Mux.scala 31:69:@15050.4]
  wire  _T_2267; // @[package.scala 96:25:@14987.4 package.scala 96:25:@14988.4]
  wire [7:0] _T_2295; // @[Mux.scala 31:69:@15051.4]
  wire  _T_2264; // @[package.scala 96:25:@14979.4 package.scala 96:25:@14980.4]
  wire [7:0] _T_2296; // @[Mux.scala 31:69:@15052.4]
  wire  _T_2261; // @[package.scala 96:25:@14971.4 package.scala 96:25:@14972.4]
  wire [7:0] _T_2297; // @[Mux.scala 31:69:@15053.4]
  wire  _T_2258; // @[package.scala 96:25:@14963.4 package.scala 96:25:@14964.4]
  wire [7:0] _T_2298; // @[Mux.scala 31:69:@15054.4]
  wire  _T_2255; // @[package.scala 96:25:@14955.4 package.scala 96:25:@14956.4]
  wire  _T_2392; // @[package.scala 96:25:@15179.4 package.scala 96:25:@15180.4]
  wire [7:0] _T_2396; // @[Mux.scala 31:69:@15189.4]
  wire  _T_2389; // @[package.scala 96:25:@15171.4 package.scala 96:25:@15172.4]
  wire [7:0] _T_2397; // @[Mux.scala 31:69:@15190.4]
  wire  _T_2386; // @[package.scala 96:25:@15163.4 package.scala 96:25:@15164.4]
  wire [7:0] _T_2398; // @[Mux.scala 31:69:@15191.4]
  wire  _T_2383; // @[package.scala 96:25:@15155.4 package.scala 96:25:@15156.4]
  wire [7:0] _T_2399; // @[Mux.scala 31:69:@15192.4]
  wire  _T_2380; // @[package.scala 96:25:@15147.4 package.scala 96:25:@15148.4]
  wire [7:0] _T_2400; // @[Mux.scala 31:69:@15193.4]
  wire  _T_2377; // @[package.scala 96:25:@15139.4 package.scala 96:25:@15140.4]
  wire [7:0] _T_2401; // @[Mux.scala 31:69:@15194.4]
  wire  _T_2374; // @[package.scala 96:25:@15131.4 package.scala 96:25:@15132.4]
  wire [7:0] _T_2402; // @[Mux.scala 31:69:@15195.4]
  wire  _T_2371; // @[package.scala 96:25:@15123.4 package.scala 96:25:@15124.4]
  wire [7:0] _T_2403; // @[Mux.scala 31:69:@15196.4]
  wire  _T_2368; // @[package.scala 96:25:@15115.4 package.scala 96:25:@15116.4]
  wire [7:0] _T_2404; // @[Mux.scala 31:69:@15197.4]
  wire  _T_2365; // @[package.scala 96:25:@15107.4 package.scala 96:25:@15108.4]
  wire [7:0] _T_2405; // @[Mux.scala 31:69:@15198.4]
  wire  _T_2362; // @[package.scala 96:25:@15099.4 package.scala 96:25:@15100.4]
  wire  _T_2499; // @[package.scala 96:25:@15323.4 package.scala 96:25:@15324.4]
  wire [7:0] _T_2503; // @[Mux.scala 31:69:@15333.4]
  wire  _T_2496; // @[package.scala 96:25:@15315.4 package.scala 96:25:@15316.4]
  wire [7:0] _T_2504; // @[Mux.scala 31:69:@15334.4]
  wire  _T_2493; // @[package.scala 96:25:@15307.4 package.scala 96:25:@15308.4]
  wire [7:0] _T_2505; // @[Mux.scala 31:69:@15335.4]
  wire  _T_2490; // @[package.scala 96:25:@15299.4 package.scala 96:25:@15300.4]
  wire [7:0] _T_2506; // @[Mux.scala 31:69:@15336.4]
  wire  _T_2487; // @[package.scala 96:25:@15291.4 package.scala 96:25:@15292.4]
  wire [7:0] _T_2507; // @[Mux.scala 31:69:@15337.4]
  wire  _T_2484; // @[package.scala 96:25:@15283.4 package.scala 96:25:@15284.4]
  wire [7:0] _T_2508; // @[Mux.scala 31:69:@15338.4]
  wire  _T_2481; // @[package.scala 96:25:@15275.4 package.scala 96:25:@15276.4]
  wire [7:0] _T_2509; // @[Mux.scala 31:69:@15339.4]
  wire  _T_2478; // @[package.scala 96:25:@15267.4 package.scala 96:25:@15268.4]
  wire [7:0] _T_2510; // @[Mux.scala 31:69:@15340.4]
  wire  _T_2475; // @[package.scala 96:25:@15259.4 package.scala 96:25:@15260.4]
  wire [7:0] _T_2511; // @[Mux.scala 31:69:@15341.4]
  wire  _T_2472; // @[package.scala 96:25:@15251.4 package.scala 96:25:@15252.4]
  wire [7:0] _T_2512; // @[Mux.scala 31:69:@15342.4]
  wire  _T_2469; // @[package.scala 96:25:@15243.4 package.scala 96:25:@15244.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@12645.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@12661.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@12677.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@12693.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@12709.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@12725.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@12741.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@12757.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@12773.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@12789.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@12805.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@12821.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  StickySelects_1 StickySelects ( // @[MemPrimitives.scala 121:29:@13017.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_ins_6(StickySelects_io_ins_6),
    .io_ins_7(StickySelects_io_ins_7),
    .io_ins_8(StickySelects_io_ins_8),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5),
    .io_outs_6(StickySelects_io_outs_6),
    .io_outs_7(StickySelects_io_outs_7),
    .io_outs_8(StickySelects_io_outs_8)
  );
  StickySelects_1 StickySelects_1 ( // @[MemPrimitives.scala 121:29:@13106.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_ins_6(StickySelects_1_io_ins_6),
    .io_ins_7(StickySelects_1_io_ins_7),
    .io_ins_8(StickySelects_1_io_ins_8),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5),
    .io_outs_6(StickySelects_1_io_outs_6),
    .io_outs_7(StickySelects_1_io_outs_7),
    .io_outs_8(StickySelects_1_io_outs_8)
  );
  StickySelects_1 StickySelects_2 ( // @[MemPrimitives.scala 121:29:@13195.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_ins_6(StickySelects_2_io_ins_6),
    .io_ins_7(StickySelects_2_io_ins_7),
    .io_ins_8(StickySelects_2_io_ins_8),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5),
    .io_outs_6(StickySelects_2_io_outs_6),
    .io_outs_7(StickySelects_2_io_outs_7),
    .io_outs_8(StickySelects_2_io_outs_8)
  );
  StickySelects_1 StickySelects_3 ( // @[MemPrimitives.scala 121:29:@13284.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_ins_6(StickySelects_3_io_ins_6),
    .io_ins_7(StickySelects_3_io_ins_7),
    .io_ins_8(StickySelects_3_io_ins_8),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5),
    .io_outs_6(StickySelects_3_io_outs_6),
    .io_outs_7(StickySelects_3_io_outs_7),
    .io_outs_8(StickySelects_3_io_outs_8)
  );
  StickySelects_1 StickySelects_4 ( // @[MemPrimitives.scala 121:29:@13373.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_ins_6(StickySelects_4_io_ins_6),
    .io_ins_7(StickySelects_4_io_ins_7),
    .io_ins_8(StickySelects_4_io_ins_8),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5),
    .io_outs_6(StickySelects_4_io_outs_6),
    .io_outs_7(StickySelects_4_io_outs_7),
    .io_outs_8(StickySelects_4_io_outs_8)
  );
  StickySelects_1 StickySelects_5 ( // @[MemPrimitives.scala 121:29:@13462.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_ins_6(StickySelects_5_io_ins_6),
    .io_ins_7(StickySelects_5_io_ins_7),
    .io_ins_8(StickySelects_5_io_ins_8),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5),
    .io_outs_6(StickySelects_5_io_outs_6),
    .io_outs_7(StickySelects_5_io_outs_7),
    .io_outs_8(StickySelects_5_io_outs_8)
  );
  StickySelects_1 StickySelects_6 ( // @[MemPrimitives.scala 121:29:@13551.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_ins_6(StickySelects_6_io_ins_6),
    .io_ins_7(StickySelects_6_io_ins_7),
    .io_ins_8(StickySelects_6_io_ins_8),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5),
    .io_outs_6(StickySelects_6_io_outs_6),
    .io_outs_7(StickySelects_6_io_outs_7),
    .io_outs_8(StickySelects_6_io_outs_8)
  );
  StickySelects_1 StickySelects_7 ( // @[MemPrimitives.scala 121:29:@13640.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_ins_6(StickySelects_7_io_ins_6),
    .io_ins_7(StickySelects_7_io_ins_7),
    .io_ins_8(StickySelects_7_io_ins_8),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5),
    .io_outs_6(StickySelects_7_io_outs_6),
    .io_outs_7(StickySelects_7_io_outs_7),
    .io_outs_8(StickySelects_7_io_outs_8)
  );
  StickySelects_1 StickySelects_8 ( // @[MemPrimitives.scala 121:29:@13729.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_ins_6(StickySelects_8_io_ins_6),
    .io_ins_7(StickySelects_8_io_ins_7),
    .io_ins_8(StickySelects_8_io_ins_8),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5),
    .io_outs_6(StickySelects_8_io_outs_6),
    .io_outs_7(StickySelects_8_io_outs_7),
    .io_outs_8(StickySelects_8_io_outs_8)
  );
  StickySelects_1 StickySelects_9 ( // @[MemPrimitives.scala 121:29:@13818.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_ins_6(StickySelects_9_io_ins_6),
    .io_ins_7(StickySelects_9_io_ins_7),
    .io_ins_8(StickySelects_9_io_ins_8),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5),
    .io_outs_6(StickySelects_9_io_outs_6),
    .io_outs_7(StickySelects_9_io_outs_7),
    .io_outs_8(StickySelects_9_io_outs_8)
  );
  StickySelects_1 StickySelects_10 ( // @[MemPrimitives.scala 121:29:@13907.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_ins_6(StickySelects_10_io_ins_6),
    .io_ins_7(StickySelects_10_io_ins_7),
    .io_ins_8(StickySelects_10_io_ins_8),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5),
    .io_outs_6(StickySelects_10_io_outs_6),
    .io_outs_7(StickySelects_10_io_outs_7),
    .io_outs_8(StickySelects_10_io_outs_8)
  );
  StickySelects_1 StickySelects_11 ( // @[MemPrimitives.scala 121:29:@13996.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_ins_6(StickySelects_11_io_ins_6),
    .io_ins_7(StickySelects_11_io_ins_7),
    .io_ins_8(StickySelects_11_io_ins_8),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5),
    .io_outs_6(StickySelects_11_io_outs_6),
    .io_outs_7(StickySelects_11_io_outs_7),
    .io_outs_8(StickySelects_11_io_outs_8)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@14086.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@14094.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@14102.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@14110.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@14118.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@14126.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@14134.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@14142.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@14150.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@14158.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@14166.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@14174.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@14230.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@14238.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@14246.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@14254.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@14262.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@14270.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@14278.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@14286.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@14294.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@14302.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@14310.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@14318.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@14374.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@14382.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@14390.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@14398.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@14406.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@14414.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@14422.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@14430.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@14438.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@14446.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@14454.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@14462.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@14518.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@14526.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@14534.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@14542.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@14550.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@14558.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@14566.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@14574.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@14582.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@14590.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@14598.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@14606.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_48 ( // @[package.scala 93:22:@14662.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@14670.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_50 ( // @[package.scala 93:22:@14678.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@14686.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@14694.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_53 ( // @[package.scala 93:22:@14702.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@14710.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_55 ( // @[package.scala 93:22:@14718.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@14726.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_57 ( // @[package.scala 93:22:@14734.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@14742.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_59 ( // @[package.scala 93:22:@14750.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_60 ( // @[package.scala 93:22:@14806.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_61 ( // @[package.scala 93:22:@14814.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_62 ( // @[package.scala 93:22:@14822.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_63 ( // @[package.scala 93:22:@14830.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_64 ( // @[package.scala 93:22:@14838.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_65 ( // @[package.scala 93:22:@14846.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_66 ( // @[package.scala 93:22:@14854.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_67 ( // @[package.scala 93:22:@14862.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_68 ( // @[package.scala 93:22:@14870.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_69 ( // @[package.scala 93:22:@14878.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_70 ( // @[package.scala 93:22:@14886.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_71 ( // @[package.scala 93:22:@14894.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_72 ( // @[package.scala 93:22:@14950.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_73 ( // @[package.scala 93:22:@14958.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_74 ( // @[package.scala 93:22:@14966.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_75 ( // @[package.scala 93:22:@14974.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_76 ( // @[package.scala 93:22:@14982.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_77 ( // @[package.scala 93:22:@14990.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_78 ( // @[package.scala 93:22:@14998.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_79 ( // @[package.scala 93:22:@15006.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_80 ( // @[package.scala 93:22:@15014.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_81 ( // @[package.scala 93:22:@15022.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_82 ( // @[package.scala 93:22:@15030.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_83 ( // @[package.scala 93:22:@15038.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_84 ( // @[package.scala 93:22:@15094.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_85 ( // @[package.scala 93:22:@15102.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_86 ( // @[package.scala 93:22:@15110.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_87 ( // @[package.scala 93:22:@15118.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_88 ( // @[package.scala 93:22:@15126.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_89 ( // @[package.scala 93:22:@15134.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_90 ( // @[package.scala 93:22:@15142.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_91 ( // @[package.scala 93:22:@15150.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_92 ( // @[package.scala 93:22:@15158.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_93 ( // @[package.scala 93:22:@15166.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_94 ( // @[package.scala 93:22:@15174.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_95 ( // @[package.scala 93:22:@15182.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_96 ( // @[package.scala 93:22:@15238.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_97 ( // @[package.scala 93:22:@15246.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_98 ( // @[package.scala 93:22:@15254.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_99 ( // @[package.scala 93:22:@15262.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_100 ( // @[package.scala 93:22:@15270.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_101 ( // @[package.scala 93:22:@15278.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_102 ( // @[package.scala 93:22:@15286.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_103 ( // @[package.scala 93:22:@15294.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_104 ( // @[package.scala 93:22:@15302.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_105 ( // @[package.scala 93:22:@15310.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_106 ( // @[package.scala 93:22:@15318.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_107 ( // @[package.scala 93:22:@15326.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  assign _T_316 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@12837.4]
  assign _T_318 = io_wPort_0_banks_1 == 2'h0; // @[MemPrimitives.scala 82:210:@12838.4]
  assign _T_319 = _T_316 & _T_318; // @[MemPrimitives.scala 82:228:@12839.4]
  assign _T_320 = io_wPort_0_en_0 & _T_319; // @[MemPrimitives.scala 83:102:@12840.4]
  assign _T_322 = {_T_320,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12842.4]
  assign _T_329 = io_wPort_0_banks_1 == 2'h1; // @[MemPrimitives.scala 82:210:@12850.4]
  assign _T_330 = _T_316 & _T_329; // @[MemPrimitives.scala 82:228:@12851.4]
  assign _T_331 = io_wPort_0_en_0 & _T_330; // @[MemPrimitives.scala 83:102:@12852.4]
  assign _T_333 = {_T_331,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12854.4]
  assign _T_340 = io_wPort_0_banks_1 == 2'h2; // @[MemPrimitives.scala 82:210:@12862.4]
  assign _T_341 = _T_316 & _T_340; // @[MemPrimitives.scala 82:228:@12863.4]
  assign _T_342 = io_wPort_0_en_0 & _T_341; // @[MemPrimitives.scala 83:102:@12864.4]
  assign _T_344 = {_T_342,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12866.4]
  assign _T_349 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@12873.4]
  assign _T_352 = _T_349 & _T_318; // @[MemPrimitives.scala 82:228:@12875.4]
  assign _T_353 = io_wPort_0_en_0 & _T_352; // @[MemPrimitives.scala 83:102:@12876.4]
  assign _T_355 = {_T_353,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12878.4]
  assign _T_363 = _T_349 & _T_329; // @[MemPrimitives.scala 82:228:@12887.4]
  assign _T_364 = io_wPort_0_en_0 & _T_363; // @[MemPrimitives.scala 83:102:@12888.4]
  assign _T_366 = {_T_364,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12890.4]
  assign _T_374 = _T_349 & _T_340; // @[MemPrimitives.scala 82:228:@12899.4]
  assign _T_375 = io_wPort_0_en_0 & _T_374; // @[MemPrimitives.scala 83:102:@12900.4]
  assign _T_377 = {_T_375,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12902.4]
  assign _T_382 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@12909.4]
  assign _T_385 = _T_382 & _T_318; // @[MemPrimitives.scala 82:228:@12911.4]
  assign _T_386 = io_wPort_0_en_0 & _T_385; // @[MemPrimitives.scala 83:102:@12912.4]
  assign _T_388 = {_T_386,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12914.4]
  assign _T_396 = _T_382 & _T_329; // @[MemPrimitives.scala 82:228:@12923.4]
  assign _T_397 = io_wPort_0_en_0 & _T_396; // @[MemPrimitives.scala 83:102:@12924.4]
  assign _T_399 = {_T_397,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12926.4]
  assign _T_407 = _T_382 & _T_340; // @[MemPrimitives.scala 82:228:@12935.4]
  assign _T_408 = io_wPort_0_en_0 & _T_407; // @[MemPrimitives.scala 83:102:@12936.4]
  assign _T_410 = {_T_408,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12938.4]
  assign _T_415 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@12945.4]
  assign _T_418 = _T_415 & _T_318; // @[MemPrimitives.scala 82:228:@12947.4]
  assign _T_419 = io_wPort_0_en_0 & _T_418; // @[MemPrimitives.scala 83:102:@12948.4]
  assign _T_421 = {_T_419,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12950.4]
  assign _T_429 = _T_415 & _T_329; // @[MemPrimitives.scala 82:228:@12959.4]
  assign _T_430 = io_wPort_0_en_0 & _T_429; // @[MemPrimitives.scala 83:102:@12960.4]
  assign _T_432 = {_T_430,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12962.4]
  assign _T_440 = _T_415 & _T_340; // @[MemPrimitives.scala 82:228:@12971.4]
  assign _T_441 = io_wPort_0_en_0 & _T_440; // @[MemPrimitives.scala 83:102:@12972.4]
  assign _T_443 = {_T_441,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12974.4]
  assign _T_448 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12981.4]
  assign _T_450 = io_rPort_0_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12982.4]
  assign _T_451 = _T_448 & _T_450; // @[MemPrimitives.scala 110:228:@12983.4]
  assign _T_454 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12985.4]
  assign _T_456 = io_rPort_1_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12986.4]
  assign _T_457 = _T_454 & _T_456; // @[MemPrimitives.scala 110:228:@12987.4]
  assign _T_460 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12989.4]
  assign _T_462 = io_rPort_2_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12990.4]
  assign _T_463 = _T_460 & _T_462; // @[MemPrimitives.scala 110:228:@12991.4]
  assign _T_466 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12993.4]
  assign _T_468 = io_rPort_3_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12994.4]
  assign _T_469 = _T_466 & _T_468; // @[MemPrimitives.scala 110:228:@12995.4]
  assign _T_472 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12997.4]
  assign _T_474 = io_rPort_4_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@12998.4]
  assign _T_475 = _T_472 & _T_474; // @[MemPrimitives.scala 110:228:@12999.4]
  assign _T_478 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13001.4]
  assign _T_480 = io_rPort_5_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13002.4]
  assign _T_481 = _T_478 & _T_480; // @[MemPrimitives.scala 110:228:@13003.4]
  assign _T_484 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13005.4]
  assign _T_486 = io_rPort_6_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13006.4]
  assign _T_487 = _T_484 & _T_486; // @[MemPrimitives.scala 110:228:@13007.4]
  assign _T_490 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13009.4]
  assign _T_492 = io_rPort_7_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13010.4]
  assign _T_493 = _T_490 & _T_492; // @[MemPrimitives.scala 110:228:@13011.4]
  assign _T_496 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13013.4]
  assign _T_498 = io_rPort_8_banks_1 == 2'h0; // @[MemPrimitives.scala 110:210:@13014.4]
  assign _T_499 = _T_496 & _T_498; // @[MemPrimitives.scala 110:228:@13015.4]
  assign _T_501 = StickySelects_io_outs_0; // @[MemPrimitives.scala 123:41:@13029.4]
  assign _T_502 = StickySelects_io_outs_1; // @[MemPrimitives.scala 123:41:@13030.4]
  assign _T_503 = StickySelects_io_outs_2; // @[MemPrimitives.scala 123:41:@13031.4]
  assign _T_504 = StickySelects_io_outs_3; // @[MemPrimitives.scala 123:41:@13032.4]
  assign _T_505 = StickySelects_io_outs_4; // @[MemPrimitives.scala 123:41:@13033.4]
  assign _T_506 = StickySelects_io_outs_5; // @[MemPrimitives.scala 123:41:@13034.4]
  assign _T_507 = StickySelects_io_outs_6; // @[MemPrimitives.scala 123:41:@13035.4]
  assign _T_508 = StickySelects_io_outs_7; // @[MemPrimitives.scala 123:41:@13036.4]
  assign _T_509 = StickySelects_io_outs_8; // @[MemPrimitives.scala 123:41:@13037.4]
  assign _T_511 = {_T_501,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13039.4]
  assign _T_513 = {_T_502,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13041.4]
  assign _T_515 = {_T_503,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13043.4]
  assign _T_517 = {_T_504,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13045.4]
  assign _T_519 = {_T_505,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13047.4]
  assign _T_521 = {_T_506,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13049.4]
  assign _T_523 = {_T_507,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13051.4]
  assign _T_525 = {_T_508,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13053.4]
  assign _T_527 = {_T_509,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13055.4]
  assign _T_528 = _T_508 ? _T_525 : _T_527; // @[Mux.scala 31:69:@13056.4]
  assign _T_529 = _T_507 ? _T_523 : _T_528; // @[Mux.scala 31:69:@13057.4]
  assign _T_530 = _T_506 ? _T_521 : _T_529; // @[Mux.scala 31:69:@13058.4]
  assign _T_531 = _T_505 ? _T_519 : _T_530; // @[Mux.scala 31:69:@13059.4]
  assign _T_532 = _T_504 ? _T_517 : _T_531; // @[Mux.scala 31:69:@13060.4]
  assign _T_533 = _T_503 ? _T_515 : _T_532; // @[Mux.scala 31:69:@13061.4]
  assign _T_534 = _T_502 ? _T_513 : _T_533; // @[Mux.scala 31:69:@13062.4]
  assign _T_535 = _T_501 ? _T_511 : _T_534; // @[Mux.scala 31:69:@13063.4]
  assign _T_542 = io_rPort_0_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13071.4]
  assign _T_543 = _T_448 & _T_542; // @[MemPrimitives.scala 110:228:@13072.4]
  assign _T_548 = io_rPort_1_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13075.4]
  assign _T_549 = _T_454 & _T_548; // @[MemPrimitives.scala 110:228:@13076.4]
  assign _T_554 = io_rPort_2_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13079.4]
  assign _T_555 = _T_460 & _T_554; // @[MemPrimitives.scala 110:228:@13080.4]
  assign _T_560 = io_rPort_3_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13083.4]
  assign _T_561 = _T_466 & _T_560; // @[MemPrimitives.scala 110:228:@13084.4]
  assign _T_566 = io_rPort_4_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13087.4]
  assign _T_567 = _T_472 & _T_566; // @[MemPrimitives.scala 110:228:@13088.4]
  assign _T_572 = io_rPort_5_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13091.4]
  assign _T_573 = _T_478 & _T_572; // @[MemPrimitives.scala 110:228:@13092.4]
  assign _T_578 = io_rPort_6_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13095.4]
  assign _T_579 = _T_484 & _T_578; // @[MemPrimitives.scala 110:228:@13096.4]
  assign _T_584 = io_rPort_7_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13099.4]
  assign _T_585 = _T_490 & _T_584; // @[MemPrimitives.scala 110:228:@13100.4]
  assign _T_590 = io_rPort_8_banks_1 == 2'h1; // @[MemPrimitives.scala 110:210:@13103.4]
  assign _T_591 = _T_496 & _T_590; // @[MemPrimitives.scala 110:228:@13104.4]
  assign _T_593 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 123:41:@13118.4]
  assign _T_594 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 123:41:@13119.4]
  assign _T_595 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 123:41:@13120.4]
  assign _T_596 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 123:41:@13121.4]
  assign _T_597 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 123:41:@13122.4]
  assign _T_598 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 123:41:@13123.4]
  assign _T_599 = StickySelects_1_io_outs_6; // @[MemPrimitives.scala 123:41:@13124.4]
  assign _T_600 = StickySelects_1_io_outs_7; // @[MemPrimitives.scala 123:41:@13125.4]
  assign _T_601 = StickySelects_1_io_outs_8; // @[MemPrimitives.scala 123:41:@13126.4]
  assign _T_603 = {_T_593,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13128.4]
  assign _T_605 = {_T_594,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13130.4]
  assign _T_607 = {_T_595,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13132.4]
  assign _T_609 = {_T_596,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13134.4]
  assign _T_611 = {_T_597,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13136.4]
  assign _T_613 = {_T_598,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13138.4]
  assign _T_615 = {_T_599,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13140.4]
  assign _T_617 = {_T_600,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13142.4]
  assign _T_619 = {_T_601,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13144.4]
  assign _T_620 = _T_600 ? _T_617 : _T_619; // @[Mux.scala 31:69:@13145.4]
  assign _T_621 = _T_599 ? _T_615 : _T_620; // @[Mux.scala 31:69:@13146.4]
  assign _T_622 = _T_598 ? _T_613 : _T_621; // @[Mux.scala 31:69:@13147.4]
  assign _T_623 = _T_597 ? _T_611 : _T_622; // @[Mux.scala 31:69:@13148.4]
  assign _T_624 = _T_596 ? _T_609 : _T_623; // @[Mux.scala 31:69:@13149.4]
  assign _T_625 = _T_595 ? _T_607 : _T_624; // @[Mux.scala 31:69:@13150.4]
  assign _T_626 = _T_594 ? _T_605 : _T_625; // @[Mux.scala 31:69:@13151.4]
  assign _T_627 = _T_593 ? _T_603 : _T_626; // @[Mux.scala 31:69:@13152.4]
  assign _T_634 = io_rPort_0_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13160.4]
  assign _T_635 = _T_448 & _T_634; // @[MemPrimitives.scala 110:228:@13161.4]
  assign _T_640 = io_rPort_1_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13164.4]
  assign _T_641 = _T_454 & _T_640; // @[MemPrimitives.scala 110:228:@13165.4]
  assign _T_646 = io_rPort_2_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13168.4]
  assign _T_647 = _T_460 & _T_646; // @[MemPrimitives.scala 110:228:@13169.4]
  assign _T_652 = io_rPort_3_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13172.4]
  assign _T_653 = _T_466 & _T_652; // @[MemPrimitives.scala 110:228:@13173.4]
  assign _T_658 = io_rPort_4_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13176.4]
  assign _T_659 = _T_472 & _T_658; // @[MemPrimitives.scala 110:228:@13177.4]
  assign _T_664 = io_rPort_5_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13180.4]
  assign _T_665 = _T_478 & _T_664; // @[MemPrimitives.scala 110:228:@13181.4]
  assign _T_670 = io_rPort_6_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13184.4]
  assign _T_671 = _T_484 & _T_670; // @[MemPrimitives.scala 110:228:@13185.4]
  assign _T_676 = io_rPort_7_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13188.4]
  assign _T_677 = _T_490 & _T_676; // @[MemPrimitives.scala 110:228:@13189.4]
  assign _T_682 = io_rPort_8_banks_1 == 2'h2; // @[MemPrimitives.scala 110:210:@13192.4]
  assign _T_683 = _T_496 & _T_682; // @[MemPrimitives.scala 110:228:@13193.4]
  assign _T_685 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 123:41:@13207.4]
  assign _T_686 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 123:41:@13208.4]
  assign _T_687 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 123:41:@13209.4]
  assign _T_688 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 123:41:@13210.4]
  assign _T_689 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 123:41:@13211.4]
  assign _T_690 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 123:41:@13212.4]
  assign _T_691 = StickySelects_2_io_outs_6; // @[MemPrimitives.scala 123:41:@13213.4]
  assign _T_692 = StickySelects_2_io_outs_7; // @[MemPrimitives.scala 123:41:@13214.4]
  assign _T_693 = StickySelects_2_io_outs_8; // @[MemPrimitives.scala 123:41:@13215.4]
  assign _T_695 = {_T_685,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13217.4]
  assign _T_697 = {_T_686,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13219.4]
  assign _T_699 = {_T_687,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13221.4]
  assign _T_701 = {_T_688,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13223.4]
  assign _T_703 = {_T_689,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13225.4]
  assign _T_705 = {_T_690,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13227.4]
  assign _T_707 = {_T_691,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13229.4]
  assign _T_709 = {_T_692,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13231.4]
  assign _T_711 = {_T_693,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13233.4]
  assign _T_712 = _T_692 ? _T_709 : _T_711; // @[Mux.scala 31:69:@13234.4]
  assign _T_713 = _T_691 ? _T_707 : _T_712; // @[Mux.scala 31:69:@13235.4]
  assign _T_714 = _T_690 ? _T_705 : _T_713; // @[Mux.scala 31:69:@13236.4]
  assign _T_715 = _T_689 ? _T_703 : _T_714; // @[Mux.scala 31:69:@13237.4]
  assign _T_716 = _T_688 ? _T_701 : _T_715; // @[Mux.scala 31:69:@13238.4]
  assign _T_717 = _T_687 ? _T_699 : _T_716; // @[Mux.scala 31:69:@13239.4]
  assign _T_718 = _T_686 ? _T_697 : _T_717; // @[Mux.scala 31:69:@13240.4]
  assign _T_719 = _T_685 ? _T_695 : _T_718; // @[Mux.scala 31:69:@13241.4]
  assign _T_724 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13248.4]
  assign _T_727 = _T_724 & _T_450; // @[MemPrimitives.scala 110:228:@13250.4]
  assign _T_730 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13252.4]
  assign _T_733 = _T_730 & _T_456; // @[MemPrimitives.scala 110:228:@13254.4]
  assign _T_736 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13256.4]
  assign _T_739 = _T_736 & _T_462; // @[MemPrimitives.scala 110:228:@13258.4]
  assign _T_742 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13260.4]
  assign _T_745 = _T_742 & _T_468; // @[MemPrimitives.scala 110:228:@13262.4]
  assign _T_748 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13264.4]
  assign _T_751 = _T_748 & _T_474; // @[MemPrimitives.scala 110:228:@13266.4]
  assign _T_754 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13268.4]
  assign _T_757 = _T_754 & _T_480; // @[MemPrimitives.scala 110:228:@13270.4]
  assign _T_760 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13272.4]
  assign _T_763 = _T_760 & _T_486; // @[MemPrimitives.scala 110:228:@13274.4]
  assign _T_766 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13276.4]
  assign _T_769 = _T_766 & _T_492; // @[MemPrimitives.scala 110:228:@13278.4]
  assign _T_772 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13280.4]
  assign _T_775 = _T_772 & _T_498; // @[MemPrimitives.scala 110:228:@13282.4]
  assign _T_777 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 123:41:@13296.4]
  assign _T_778 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 123:41:@13297.4]
  assign _T_779 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 123:41:@13298.4]
  assign _T_780 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 123:41:@13299.4]
  assign _T_781 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 123:41:@13300.4]
  assign _T_782 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 123:41:@13301.4]
  assign _T_783 = StickySelects_3_io_outs_6; // @[MemPrimitives.scala 123:41:@13302.4]
  assign _T_784 = StickySelects_3_io_outs_7; // @[MemPrimitives.scala 123:41:@13303.4]
  assign _T_785 = StickySelects_3_io_outs_8; // @[MemPrimitives.scala 123:41:@13304.4]
  assign _T_787 = {_T_777,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13306.4]
  assign _T_789 = {_T_778,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13308.4]
  assign _T_791 = {_T_779,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13310.4]
  assign _T_793 = {_T_780,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13312.4]
  assign _T_795 = {_T_781,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13314.4]
  assign _T_797 = {_T_782,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13316.4]
  assign _T_799 = {_T_783,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13318.4]
  assign _T_801 = {_T_784,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13320.4]
  assign _T_803 = {_T_785,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13322.4]
  assign _T_804 = _T_784 ? _T_801 : _T_803; // @[Mux.scala 31:69:@13323.4]
  assign _T_805 = _T_783 ? _T_799 : _T_804; // @[Mux.scala 31:69:@13324.4]
  assign _T_806 = _T_782 ? _T_797 : _T_805; // @[Mux.scala 31:69:@13325.4]
  assign _T_807 = _T_781 ? _T_795 : _T_806; // @[Mux.scala 31:69:@13326.4]
  assign _T_808 = _T_780 ? _T_793 : _T_807; // @[Mux.scala 31:69:@13327.4]
  assign _T_809 = _T_779 ? _T_791 : _T_808; // @[Mux.scala 31:69:@13328.4]
  assign _T_810 = _T_778 ? _T_789 : _T_809; // @[Mux.scala 31:69:@13329.4]
  assign _T_811 = _T_777 ? _T_787 : _T_810; // @[Mux.scala 31:69:@13330.4]
  assign _T_819 = _T_724 & _T_542; // @[MemPrimitives.scala 110:228:@13339.4]
  assign _T_825 = _T_730 & _T_548; // @[MemPrimitives.scala 110:228:@13343.4]
  assign _T_831 = _T_736 & _T_554; // @[MemPrimitives.scala 110:228:@13347.4]
  assign _T_837 = _T_742 & _T_560; // @[MemPrimitives.scala 110:228:@13351.4]
  assign _T_843 = _T_748 & _T_566; // @[MemPrimitives.scala 110:228:@13355.4]
  assign _T_849 = _T_754 & _T_572; // @[MemPrimitives.scala 110:228:@13359.4]
  assign _T_855 = _T_760 & _T_578; // @[MemPrimitives.scala 110:228:@13363.4]
  assign _T_861 = _T_766 & _T_584; // @[MemPrimitives.scala 110:228:@13367.4]
  assign _T_867 = _T_772 & _T_590; // @[MemPrimitives.scala 110:228:@13371.4]
  assign _T_869 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 123:41:@13385.4]
  assign _T_870 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 123:41:@13386.4]
  assign _T_871 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 123:41:@13387.4]
  assign _T_872 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 123:41:@13388.4]
  assign _T_873 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 123:41:@13389.4]
  assign _T_874 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 123:41:@13390.4]
  assign _T_875 = StickySelects_4_io_outs_6; // @[MemPrimitives.scala 123:41:@13391.4]
  assign _T_876 = StickySelects_4_io_outs_7; // @[MemPrimitives.scala 123:41:@13392.4]
  assign _T_877 = StickySelects_4_io_outs_8; // @[MemPrimitives.scala 123:41:@13393.4]
  assign _T_879 = {_T_869,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13395.4]
  assign _T_881 = {_T_870,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13397.4]
  assign _T_883 = {_T_871,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13399.4]
  assign _T_885 = {_T_872,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13401.4]
  assign _T_887 = {_T_873,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13403.4]
  assign _T_889 = {_T_874,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13405.4]
  assign _T_891 = {_T_875,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13407.4]
  assign _T_893 = {_T_876,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13409.4]
  assign _T_895 = {_T_877,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13411.4]
  assign _T_896 = _T_876 ? _T_893 : _T_895; // @[Mux.scala 31:69:@13412.4]
  assign _T_897 = _T_875 ? _T_891 : _T_896; // @[Mux.scala 31:69:@13413.4]
  assign _T_898 = _T_874 ? _T_889 : _T_897; // @[Mux.scala 31:69:@13414.4]
  assign _T_899 = _T_873 ? _T_887 : _T_898; // @[Mux.scala 31:69:@13415.4]
  assign _T_900 = _T_872 ? _T_885 : _T_899; // @[Mux.scala 31:69:@13416.4]
  assign _T_901 = _T_871 ? _T_883 : _T_900; // @[Mux.scala 31:69:@13417.4]
  assign _T_902 = _T_870 ? _T_881 : _T_901; // @[Mux.scala 31:69:@13418.4]
  assign _T_903 = _T_869 ? _T_879 : _T_902; // @[Mux.scala 31:69:@13419.4]
  assign _T_911 = _T_724 & _T_634; // @[MemPrimitives.scala 110:228:@13428.4]
  assign _T_917 = _T_730 & _T_640; // @[MemPrimitives.scala 110:228:@13432.4]
  assign _T_923 = _T_736 & _T_646; // @[MemPrimitives.scala 110:228:@13436.4]
  assign _T_929 = _T_742 & _T_652; // @[MemPrimitives.scala 110:228:@13440.4]
  assign _T_935 = _T_748 & _T_658; // @[MemPrimitives.scala 110:228:@13444.4]
  assign _T_941 = _T_754 & _T_664; // @[MemPrimitives.scala 110:228:@13448.4]
  assign _T_947 = _T_760 & _T_670; // @[MemPrimitives.scala 110:228:@13452.4]
  assign _T_953 = _T_766 & _T_676; // @[MemPrimitives.scala 110:228:@13456.4]
  assign _T_959 = _T_772 & _T_682; // @[MemPrimitives.scala 110:228:@13460.4]
  assign _T_961 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 123:41:@13474.4]
  assign _T_962 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 123:41:@13475.4]
  assign _T_963 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 123:41:@13476.4]
  assign _T_964 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 123:41:@13477.4]
  assign _T_965 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 123:41:@13478.4]
  assign _T_966 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 123:41:@13479.4]
  assign _T_967 = StickySelects_5_io_outs_6; // @[MemPrimitives.scala 123:41:@13480.4]
  assign _T_968 = StickySelects_5_io_outs_7; // @[MemPrimitives.scala 123:41:@13481.4]
  assign _T_969 = StickySelects_5_io_outs_8; // @[MemPrimitives.scala 123:41:@13482.4]
  assign _T_971 = {_T_961,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13484.4]
  assign _T_973 = {_T_962,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13486.4]
  assign _T_975 = {_T_963,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13488.4]
  assign _T_977 = {_T_964,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13490.4]
  assign _T_979 = {_T_965,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13492.4]
  assign _T_981 = {_T_966,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13494.4]
  assign _T_983 = {_T_967,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13496.4]
  assign _T_985 = {_T_968,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13498.4]
  assign _T_987 = {_T_969,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13500.4]
  assign _T_988 = _T_968 ? _T_985 : _T_987; // @[Mux.scala 31:69:@13501.4]
  assign _T_989 = _T_967 ? _T_983 : _T_988; // @[Mux.scala 31:69:@13502.4]
  assign _T_990 = _T_966 ? _T_981 : _T_989; // @[Mux.scala 31:69:@13503.4]
  assign _T_991 = _T_965 ? _T_979 : _T_990; // @[Mux.scala 31:69:@13504.4]
  assign _T_992 = _T_964 ? _T_977 : _T_991; // @[Mux.scala 31:69:@13505.4]
  assign _T_993 = _T_963 ? _T_975 : _T_992; // @[Mux.scala 31:69:@13506.4]
  assign _T_994 = _T_962 ? _T_973 : _T_993; // @[Mux.scala 31:69:@13507.4]
  assign _T_995 = _T_961 ? _T_971 : _T_994; // @[Mux.scala 31:69:@13508.4]
  assign _T_1000 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13515.4]
  assign _T_1003 = _T_1000 & _T_450; // @[MemPrimitives.scala 110:228:@13517.4]
  assign _T_1006 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13519.4]
  assign _T_1009 = _T_1006 & _T_456; // @[MemPrimitives.scala 110:228:@13521.4]
  assign _T_1012 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13523.4]
  assign _T_1015 = _T_1012 & _T_462; // @[MemPrimitives.scala 110:228:@13525.4]
  assign _T_1018 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13527.4]
  assign _T_1021 = _T_1018 & _T_468; // @[MemPrimitives.scala 110:228:@13529.4]
  assign _T_1024 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13531.4]
  assign _T_1027 = _T_1024 & _T_474; // @[MemPrimitives.scala 110:228:@13533.4]
  assign _T_1030 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13535.4]
  assign _T_1033 = _T_1030 & _T_480; // @[MemPrimitives.scala 110:228:@13537.4]
  assign _T_1036 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13539.4]
  assign _T_1039 = _T_1036 & _T_486; // @[MemPrimitives.scala 110:228:@13541.4]
  assign _T_1042 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13543.4]
  assign _T_1045 = _T_1042 & _T_492; // @[MemPrimitives.scala 110:228:@13545.4]
  assign _T_1048 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13547.4]
  assign _T_1051 = _T_1048 & _T_498; // @[MemPrimitives.scala 110:228:@13549.4]
  assign _T_1053 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 123:41:@13563.4]
  assign _T_1054 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 123:41:@13564.4]
  assign _T_1055 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 123:41:@13565.4]
  assign _T_1056 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 123:41:@13566.4]
  assign _T_1057 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 123:41:@13567.4]
  assign _T_1058 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 123:41:@13568.4]
  assign _T_1059 = StickySelects_6_io_outs_6; // @[MemPrimitives.scala 123:41:@13569.4]
  assign _T_1060 = StickySelects_6_io_outs_7; // @[MemPrimitives.scala 123:41:@13570.4]
  assign _T_1061 = StickySelects_6_io_outs_8; // @[MemPrimitives.scala 123:41:@13571.4]
  assign _T_1063 = {_T_1053,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13573.4]
  assign _T_1065 = {_T_1054,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13575.4]
  assign _T_1067 = {_T_1055,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13577.4]
  assign _T_1069 = {_T_1056,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13579.4]
  assign _T_1071 = {_T_1057,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13581.4]
  assign _T_1073 = {_T_1058,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13583.4]
  assign _T_1075 = {_T_1059,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13585.4]
  assign _T_1077 = {_T_1060,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13587.4]
  assign _T_1079 = {_T_1061,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13589.4]
  assign _T_1080 = _T_1060 ? _T_1077 : _T_1079; // @[Mux.scala 31:69:@13590.4]
  assign _T_1081 = _T_1059 ? _T_1075 : _T_1080; // @[Mux.scala 31:69:@13591.4]
  assign _T_1082 = _T_1058 ? _T_1073 : _T_1081; // @[Mux.scala 31:69:@13592.4]
  assign _T_1083 = _T_1057 ? _T_1071 : _T_1082; // @[Mux.scala 31:69:@13593.4]
  assign _T_1084 = _T_1056 ? _T_1069 : _T_1083; // @[Mux.scala 31:69:@13594.4]
  assign _T_1085 = _T_1055 ? _T_1067 : _T_1084; // @[Mux.scala 31:69:@13595.4]
  assign _T_1086 = _T_1054 ? _T_1065 : _T_1085; // @[Mux.scala 31:69:@13596.4]
  assign _T_1087 = _T_1053 ? _T_1063 : _T_1086; // @[Mux.scala 31:69:@13597.4]
  assign _T_1095 = _T_1000 & _T_542; // @[MemPrimitives.scala 110:228:@13606.4]
  assign _T_1101 = _T_1006 & _T_548; // @[MemPrimitives.scala 110:228:@13610.4]
  assign _T_1107 = _T_1012 & _T_554; // @[MemPrimitives.scala 110:228:@13614.4]
  assign _T_1113 = _T_1018 & _T_560; // @[MemPrimitives.scala 110:228:@13618.4]
  assign _T_1119 = _T_1024 & _T_566; // @[MemPrimitives.scala 110:228:@13622.4]
  assign _T_1125 = _T_1030 & _T_572; // @[MemPrimitives.scala 110:228:@13626.4]
  assign _T_1131 = _T_1036 & _T_578; // @[MemPrimitives.scala 110:228:@13630.4]
  assign _T_1137 = _T_1042 & _T_584; // @[MemPrimitives.scala 110:228:@13634.4]
  assign _T_1143 = _T_1048 & _T_590; // @[MemPrimitives.scala 110:228:@13638.4]
  assign _T_1145 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 123:41:@13652.4]
  assign _T_1146 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 123:41:@13653.4]
  assign _T_1147 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 123:41:@13654.4]
  assign _T_1148 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 123:41:@13655.4]
  assign _T_1149 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 123:41:@13656.4]
  assign _T_1150 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 123:41:@13657.4]
  assign _T_1151 = StickySelects_7_io_outs_6; // @[MemPrimitives.scala 123:41:@13658.4]
  assign _T_1152 = StickySelects_7_io_outs_7; // @[MemPrimitives.scala 123:41:@13659.4]
  assign _T_1153 = StickySelects_7_io_outs_8; // @[MemPrimitives.scala 123:41:@13660.4]
  assign _T_1155 = {_T_1145,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13662.4]
  assign _T_1157 = {_T_1146,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13664.4]
  assign _T_1159 = {_T_1147,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13666.4]
  assign _T_1161 = {_T_1148,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13668.4]
  assign _T_1163 = {_T_1149,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13670.4]
  assign _T_1165 = {_T_1150,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13672.4]
  assign _T_1167 = {_T_1151,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13674.4]
  assign _T_1169 = {_T_1152,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13676.4]
  assign _T_1171 = {_T_1153,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13678.4]
  assign _T_1172 = _T_1152 ? _T_1169 : _T_1171; // @[Mux.scala 31:69:@13679.4]
  assign _T_1173 = _T_1151 ? _T_1167 : _T_1172; // @[Mux.scala 31:69:@13680.4]
  assign _T_1174 = _T_1150 ? _T_1165 : _T_1173; // @[Mux.scala 31:69:@13681.4]
  assign _T_1175 = _T_1149 ? _T_1163 : _T_1174; // @[Mux.scala 31:69:@13682.4]
  assign _T_1176 = _T_1148 ? _T_1161 : _T_1175; // @[Mux.scala 31:69:@13683.4]
  assign _T_1177 = _T_1147 ? _T_1159 : _T_1176; // @[Mux.scala 31:69:@13684.4]
  assign _T_1178 = _T_1146 ? _T_1157 : _T_1177; // @[Mux.scala 31:69:@13685.4]
  assign _T_1179 = _T_1145 ? _T_1155 : _T_1178; // @[Mux.scala 31:69:@13686.4]
  assign _T_1187 = _T_1000 & _T_634; // @[MemPrimitives.scala 110:228:@13695.4]
  assign _T_1193 = _T_1006 & _T_640; // @[MemPrimitives.scala 110:228:@13699.4]
  assign _T_1199 = _T_1012 & _T_646; // @[MemPrimitives.scala 110:228:@13703.4]
  assign _T_1205 = _T_1018 & _T_652; // @[MemPrimitives.scala 110:228:@13707.4]
  assign _T_1211 = _T_1024 & _T_658; // @[MemPrimitives.scala 110:228:@13711.4]
  assign _T_1217 = _T_1030 & _T_664; // @[MemPrimitives.scala 110:228:@13715.4]
  assign _T_1223 = _T_1036 & _T_670; // @[MemPrimitives.scala 110:228:@13719.4]
  assign _T_1229 = _T_1042 & _T_676; // @[MemPrimitives.scala 110:228:@13723.4]
  assign _T_1235 = _T_1048 & _T_682; // @[MemPrimitives.scala 110:228:@13727.4]
  assign _T_1237 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 123:41:@13741.4]
  assign _T_1238 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 123:41:@13742.4]
  assign _T_1239 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 123:41:@13743.4]
  assign _T_1240 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 123:41:@13744.4]
  assign _T_1241 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 123:41:@13745.4]
  assign _T_1242 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 123:41:@13746.4]
  assign _T_1243 = StickySelects_8_io_outs_6; // @[MemPrimitives.scala 123:41:@13747.4]
  assign _T_1244 = StickySelects_8_io_outs_7; // @[MemPrimitives.scala 123:41:@13748.4]
  assign _T_1245 = StickySelects_8_io_outs_8; // @[MemPrimitives.scala 123:41:@13749.4]
  assign _T_1247 = {_T_1237,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13751.4]
  assign _T_1249 = {_T_1238,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13753.4]
  assign _T_1251 = {_T_1239,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13755.4]
  assign _T_1253 = {_T_1240,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13757.4]
  assign _T_1255 = {_T_1241,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13759.4]
  assign _T_1257 = {_T_1242,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13761.4]
  assign _T_1259 = {_T_1243,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13763.4]
  assign _T_1261 = {_T_1244,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13765.4]
  assign _T_1263 = {_T_1245,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13767.4]
  assign _T_1264 = _T_1244 ? _T_1261 : _T_1263; // @[Mux.scala 31:69:@13768.4]
  assign _T_1265 = _T_1243 ? _T_1259 : _T_1264; // @[Mux.scala 31:69:@13769.4]
  assign _T_1266 = _T_1242 ? _T_1257 : _T_1265; // @[Mux.scala 31:69:@13770.4]
  assign _T_1267 = _T_1241 ? _T_1255 : _T_1266; // @[Mux.scala 31:69:@13771.4]
  assign _T_1268 = _T_1240 ? _T_1253 : _T_1267; // @[Mux.scala 31:69:@13772.4]
  assign _T_1269 = _T_1239 ? _T_1251 : _T_1268; // @[Mux.scala 31:69:@13773.4]
  assign _T_1270 = _T_1238 ? _T_1249 : _T_1269; // @[Mux.scala 31:69:@13774.4]
  assign _T_1271 = _T_1237 ? _T_1247 : _T_1270; // @[Mux.scala 31:69:@13775.4]
  assign _T_1276 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13782.4]
  assign _T_1279 = _T_1276 & _T_450; // @[MemPrimitives.scala 110:228:@13784.4]
  assign _T_1282 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13786.4]
  assign _T_1285 = _T_1282 & _T_456; // @[MemPrimitives.scala 110:228:@13788.4]
  assign _T_1288 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13790.4]
  assign _T_1291 = _T_1288 & _T_462; // @[MemPrimitives.scala 110:228:@13792.4]
  assign _T_1294 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13794.4]
  assign _T_1297 = _T_1294 & _T_468; // @[MemPrimitives.scala 110:228:@13796.4]
  assign _T_1300 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13798.4]
  assign _T_1303 = _T_1300 & _T_474; // @[MemPrimitives.scala 110:228:@13800.4]
  assign _T_1306 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13802.4]
  assign _T_1309 = _T_1306 & _T_480; // @[MemPrimitives.scala 110:228:@13804.4]
  assign _T_1312 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13806.4]
  assign _T_1315 = _T_1312 & _T_486; // @[MemPrimitives.scala 110:228:@13808.4]
  assign _T_1318 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13810.4]
  assign _T_1321 = _T_1318 & _T_492; // @[MemPrimitives.scala 110:228:@13812.4]
  assign _T_1324 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13814.4]
  assign _T_1327 = _T_1324 & _T_498; // @[MemPrimitives.scala 110:228:@13816.4]
  assign _T_1329 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 123:41:@13830.4]
  assign _T_1330 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 123:41:@13831.4]
  assign _T_1331 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 123:41:@13832.4]
  assign _T_1332 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 123:41:@13833.4]
  assign _T_1333 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 123:41:@13834.4]
  assign _T_1334 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 123:41:@13835.4]
  assign _T_1335 = StickySelects_9_io_outs_6; // @[MemPrimitives.scala 123:41:@13836.4]
  assign _T_1336 = StickySelects_9_io_outs_7; // @[MemPrimitives.scala 123:41:@13837.4]
  assign _T_1337 = StickySelects_9_io_outs_8; // @[MemPrimitives.scala 123:41:@13838.4]
  assign _T_1339 = {_T_1329,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13840.4]
  assign _T_1341 = {_T_1330,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13842.4]
  assign _T_1343 = {_T_1331,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13844.4]
  assign _T_1345 = {_T_1332,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13846.4]
  assign _T_1347 = {_T_1333,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13848.4]
  assign _T_1349 = {_T_1334,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13850.4]
  assign _T_1351 = {_T_1335,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13852.4]
  assign _T_1353 = {_T_1336,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13854.4]
  assign _T_1355 = {_T_1337,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13856.4]
  assign _T_1356 = _T_1336 ? _T_1353 : _T_1355; // @[Mux.scala 31:69:@13857.4]
  assign _T_1357 = _T_1335 ? _T_1351 : _T_1356; // @[Mux.scala 31:69:@13858.4]
  assign _T_1358 = _T_1334 ? _T_1349 : _T_1357; // @[Mux.scala 31:69:@13859.4]
  assign _T_1359 = _T_1333 ? _T_1347 : _T_1358; // @[Mux.scala 31:69:@13860.4]
  assign _T_1360 = _T_1332 ? _T_1345 : _T_1359; // @[Mux.scala 31:69:@13861.4]
  assign _T_1361 = _T_1331 ? _T_1343 : _T_1360; // @[Mux.scala 31:69:@13862.4]
  assign _T_1362 = _T_1330 ? _T_1341 : _T_1361; // @[Mux.scala 31:69:@13863.4]
  assign _T_1363 = _T_1329 ? _T_1339 : _T_1362; // @[Mux.scala 31:69:@13864.4]
  assign _T_1371 = _T_1276 & _T_542; // @[MemPrimitives.scala 110:228:@13873.4]
  assign _T_1377 = _T_1282 & _T_548; // @[MemPrimitives.scala 110:228:@13877.4]
  assign _T_1383 = _T_1288 & _T_554; // @[MemPrimitives.scala 110:228:@13881.4]
  assign _T_1389 = _T_1294 & _T_560; // @[MemPrimitives.scala 110:228:@13885.4]
  assign _T_1395 = _T_1300 & _T_566; // @[MemPrimitives.scala 110:228:@13889.4]
  assign _T_1401 = _T_1306 & _T_572; // @[MemPrimitives.scala 110:228:@13893.4]
  assign _T_1407 = _T_1312 & _T_578; // @[MemPrimitives.scala 110:228:@13897.4]
  assign _T_1413 = _T_1318 & _T_584; // @[MemPrimitives.scala 110:228:@13901.4]
  assign _T_1419 = _T_1324 & _T_590; // @[MemPrimitives.scala 110:228:@13905.4]
  assign _T_1421 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 123:41:@13919.4]
  assign _T_1422 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 123:41:@13920.4]
  assign _T_1423 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 123:41:@13921.4]
  assign _T_1424 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 123:41:@13922.4]
  assign _T_1425 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 123:41:@13923.4]
  assign _T_1426 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 123:41:@13924.4]
  assign _T_1427 = StickySelects_10_io_outs_6; // @[MemPrimitives.scala 123:41:@13925.4]
  assign _T_1428 = StickySelects_10_io_outs_7; // @[MemPrimitives.scala 123:41:@13926.4]
  assign _T_1429 = StickySelects_10_io_outs_8; // @[MemPrimitives.scala 123:41:@13927.4]
  assign _T_1431 = {_T_1421,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13929.4]
  assign _T_1433 = {_T_1422,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13931.4]
  assign _T_1435 = {_T_1423,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13933.4]
  assign _T_1437 = {_T_1424,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13935.4]
  assign _T_1439 = {_T_1425,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13937.4]
  assign _T_1441 = {_T_1426,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13939.4]
  assign _T_1443 = {_T_1427,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13941.4]
  assign _T_1445 = {_T_1428,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13943.4]
  assign _T_1447 = {_T_1429,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13945.4]
  assign _T_1448 = _T_1428 ? _T_1445 : _T_1447; // @[Mux.scala 31:69:@13946.4]
  assign _T_1449 = _T_1427 ? _T_1443 : _T_1448; // @[Mux.scala 31:69:@13947.4]
  assign _T_1450 = _T_1426 ? _T_1441 : _T_1449; // @[Mux.scala 31:69:@13948.4]
  assign _T_1451 = _T_1425 ? _T_1439 : _T_1450; // @[Mux.scala 31:69:@13949.4]
  assign _T_1452 = _T_1424 ? _T_1437 : _T_1451; // @[Mux.scala 31:69:@13950.4]
  assign _T_1453 = _T_1423 ? _T_1435 : _T_1452; // @[Mux.scala 31:69:@13951.4]
  assign _T_1454 = _T_1422 ? _T_1433 : _T_1453; // @[Mux.scala 31:69:@13952.4]
  assign _T_1455 = _T_1421 ? _T_1431 : _T_1454; // @[Mux.scala 31:69:@13953.4]
  assign _T_1463 = _T_1276 & _T_634; // @[MemPrimitives.scala 110:228:@13962.4]
  assign _T_1469 = _T_1282 & _T_640; // @[MemPrimitives.scala 110:228:@13966.4]
  assign _T_1475 = _T_1288 & _T_646; // @[MemPrimitives.scala 110:228:@13970.4]
  assign _T_1481 = _T_1294 & _T_652; // @[MemPrimitives.scala 110:228:@13974.4]
  assign _T_1487 = _T_1300 & _T_658; // @[MemPrimitives.scala 110:228:@13978.4]
  assign _T_1493 = _T_1306 & _T_664; // @[MemPrimitives.scala 110:228:@13982.4]
  assign _T_1499 = _T_1312 & _T_670; // @[MemPrimitives.scala 110:228:@13986.4]
  assign _T_1505 = _T_1318 & _T_676; // @[MemPrimitives.scala 110:228:@13990.4]
  assign _T_1511 = _T_1324 & _T_682; // @[MemPrimitives.scala 110:228:@13994.4]
  assign _T_1513 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 123:41:@14008.4]
  assign _T_1514 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 123:41:@14009.4]
  assign _T_1515 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 123:41:@14010.4]
  assign _T_1516 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 123:41:@14011.4]
  assign _T_1517 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 123:41:@14012.4]
  assign _T_1518 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 123:41:@14013.4]
  assign _T_1519 = StickySelects_11_io_outs_6; // @[MemPrimitives.scala 123:41:@14014.4]
  assign _T_1520 = StickySelects_11_io_outs_7; // @[MemPrimitives.scala 123:41:@14015.4]
  assign _T_1521 = StickySelects_11_io_outs_8; // @[MemPrimitives.scala 123:41:@14016.4]
  assign _T_1523 = {_T_1513,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@14018.4]
  assign _T_1525 = {_T_1514,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@14020.4]
  assign _T_1527 = {_T_1515,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@14022.4]
  assign _T_1529 = {_T_1516,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@14024.4]
  assign _T_1531 = {_T_1517,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@14026.4]
  assign _T_1533 = {_T_1518,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@14028.4]
  assign _T_1535 = {_T_1519,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@14030.4]
  assign _T_1537 = {_T_1520,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@14032.4]
  assign _T_1539 = {_T_1521,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@14034.4]
  assign _T_1540 = _T_1520 ? _T_1537 : _T_1539; // @[Mux.scala 31:69:@14035.4]
  assign _T_1541 = _T_1519 ? _T_1535 : _T_1540; // @[Mux.scala 31:69:@14036.4]
  assign _T_1542 = _T_1518 ? _T_1533 : _T_1541; // @[Mux.scala 31:69:@14037.4]
  assign _T_1543 = _T_1517 ? _T_1531 : _T_1542; // @[Mux.scala 31:69:@14038.4]
  assign _T_1544 = _T_1516 ? _T_1529 : _T_1543; // @[Mux.scala 31:69:@14039.4]
  assign _T_1545 = _T_1515 ? _T_1527 : _T_1544; // @[Mux.scala 31:69:@14040.4]
  assign _T_1546 = _T_1514 ? _T_1525 : _T_1545; // @[Mux.scala 31:69:@14041.4]
  assign _T_1547 = _T_1513 ? _T_1523 : _T_1546; // @[Mux.scala 31:69:@14042.4]
  assign _T_1643 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@14171.4 package.scala 96:25:@14172.4]
  assign _T_1647 = _T_1643 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14181.4]
  assign _T_1640 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@14163.4 package.scala 96:25:@14164.4]
  assign _T_1648 = _T_1640 ? Mem1D_9_io_output : _T_1647; // @[Mux.scala 31:69:@14182.4]
  assign _T_1637 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@14155.4 package.scala 96:25:@14156.4]
  assign _T_1649 = _T_1637 ? Mem1D_8_io_output : _T_1648; // @[Mux.scala 31:69:@14183.4]
  assign _T_1634 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@14147.4 package.scala 96:25:@14148.4]
  assign _T_1650 = _T_1634 ? Mem1D_7_io_output : _T_1649; // @[Mux.scala 31:69:@14184.4]
  assign _T_1631 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@14139.4 package.scala 96:25:@14140.4]
  assign _T_1651 = _T_1631 ? Mem1D_6_io_output : _T_1650; // @[Mux.scala 31:69:@14185.4]
  assign _T_1628 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@14131.4 package.scala 96:25:@14132.4]
  assign _T_1652 = _T_1628 ? Mem1D_5_io_output : _T_1651; // @[Mux.scala 31:69:@14186.4]
  assign _T_1625 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@14123.4 package.scala 96:25:@14124.4]
  assign _T_1653 = _T_1625 ? Mem1D_4_io_output : _T_1652; // @[Mux.scala 31:69:@14187.4]
  assign _T_1622 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@14115.4 package.scala 96:25:@14116.4]
  assign _T_1654 = _T_1622 ? Mem1D_3_io_output : _T_1653; // @[Mux.scala 31:69:@14188.4]
  assign _T_1619 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@14107.4 package.scala 96:25:@14108.4]
  assign _T_1655 = _T_1619 ? Mem1D_2_io_output : _T_1654; // @[Mux.scala 31:69:@14189.4]
  assign _T_1616 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@14099.4 package.scala 96:25:@14100.4]
  assign _T_1656 = _T_1616 ? Mem1D_1_io_output : _T_1655; // @[Mux.scala 31:69:@14190.4]
  assign _T_1613 = RetimeWrapper_io_out; // @[package.scala 96:25:@14091.4 package.scala 96:25:@14092.4]
  assign _T_1750 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@14315.4 package.scala 96:25:@14316.4]
  assign _T_1754 = _T_1750 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14325.4]
  assign _T_1747 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@14307.4 package.scala 96:25:@14308.4]
  assign _T_1755 = _T_1747 ? Mem1D_9_io_output : _T_1754; // @[Mux.scala 31:69:@14326.4]
  assign _T_1744 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@14299.4 package.scala 96:25:@14300.4]
  assign _T_1756 = _T_1744 ? Mem1D_8_io_output : _T_1755; // @[Mux.scala 31:69:@14327.4]
  assign _T_1741 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@14291.4 package.scala 96:25:@14292.4]
  assign _T_1757 = _T_1741 ? Mem1D_7_io_output : _T_1756; // @[Mux.scala 31:69:@14328.4]
  assign _T_1738 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@14283.4 package.scala 96:25:@14284.4]
  assign _T_1758 = _T_1738 ? Mem1D_6_io_output : _T_1757; // @[Mux.scala 31:69:@14329.4]
  assign _T_1735 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@14275.4 package.scala 96:25:@14276.4]
  assign _T_1759 = _T_1735 ? Mem1D_5_io_output : _T_1758; // @[Mux.scala 31:69:@14330.4]
  assign _T_1732 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@14267.4 package.scala 96:25:@14268.4]
  assign _T_1760 = _T_1732 ? Mem1D_4_io_output : _T_1759; // @[Mux.scala 31:69:@14331.4]
  assign _T_1729 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@14259.4 package.scala 96:25:@14260.4]
  assign _T_1761 = _T_1729 ? Mem1D_3_io_output : _T_1760; // @[Mux.scala 31:69:@14332.4]
  assign _T_1726 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@14251.4 package.scala 96:25:@14252.4]
  assign _T_1762 = _T_1726 ? Mem1D_2_io_output : _T_1761; // @[Mux.scala 31:69:@14333.4]
  assign _T_1723 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@14243.4 package.scala 96:25:@14244.4]
  assign _T_1763 = _T_1723 ? Mem1D_1_io_output : _T_1762; // @[Mux.scala 31:69:@14334.4]
  assign _T_1720 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@14235.4 package.scala 96:25:@14236.4]
  assign _T_1857 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@14459.4 package.scala 96:25:@14460.4]
  assign _T_1861 = _T_1857 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14469.4]
  assign _T_1854 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@14451.4 package.scala 96:25:@14452.4]
  assign _T_1862 = _T_1854 ? Mem1D_9_io_output : _T_1861; // @[Mux.scala 31:69:@14470.4]
  assign _T_1851 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@14443.4 package.scala 96:25:@14444.4]
  assign _T_1863 = _T_1851 ? Mem1D_8_io_output : _T_1862; // @[Mux.scala 31:69:@14471.4]
  assign _T_1848 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@14435.4 package.scala 96:25:@14436.4]
  assign _T_1864 = _T_1848 ? Mem1D_7_io_output : _T_1863; // @[Mux.scala 31:69:@14472.4]
  assign _T_1845 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@14427.4 package.scala 96:25:@14428.4]
  assign _T_1865 = _T_1845 ? Mem1D_6_io_output : _T_1864; // @[Mux.scala 31:69:@14473.4]
  assign _T_1842 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@14419.4 package.scala 96:25:@14420.4]
  assign _T_1866 = _T_1842 ? Mem1D_5_io_output : _T_1865; // @[Mux.scala 31:69:@14474.4]
  assign _T_1839 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@14411.4 package.scala 96:25:@14412.4]
  assign _T_1867 = _T_1839 ? Mem1D_4_io_output : _T_1866; // @[Mux.scala 31:69:@14475.4]
  assign _T_1836 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@14403.4 package.scala 96:25:@14404.4]
  assign _T_1868 = _T_1836 ? Mem1D_3_io_output : _T_1867; // @[Mux.scala 31:69:@14476.4]
  assign _T_1833 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@14395.4 package.scala 96:25:@14396.4]
  assign _T_1869 = _T_1833 ? Mem1D_2_io_output : _T_1868; // @[Mux.scala 31:69:@14477.4]
  assign _T_1830 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@14387.4 package.scala 96:25:@14388.4]
  assign _T_1870 = _T_1830 ? Mem1D_1_io_output : _T_1869; // @[Mux.scala 31:69:@14478.4]
  assign _T_1827 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@14379.4 package.scala 96:25:@14380.4]
  assign _T_1964 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@14603.4 package.scala 96:25:@14604.4]
  assign _T_1968 = _T_1964 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14613.4]
  assign _T_1961 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@14595.4 package.scala 96:25:@14596.4]
  assign _T_1969 = _T_1961 ? Mem1D_9_io_output : _T_1968; // @[Mux.scala 31:69:@14614.4]
  assign _T_1958 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@14587.4 package.scala 96:25:@14588.4]
  assign _T_1970 = _T_1958 ? Mem1D_8_io_output : _T_1969; // @[Mux.scala 31:69:@14615.4]
  assign _T_1955 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@14579.4 package.scala 96:25:@14580.4]
  assign _T_1971 = _T_1955 ? Mem1D_7_io_output : _T_1970; // @[Mux.scala 31:69:@14616.4]
  assign _T_1952 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@14571.4 package.scala 96:25:@14572.4]
  assign _T_1972 = _T_1952 ? Mem1D_6_io_output : _T_1971; // @[Mux.scala 31:69:@14617.4]
  assign _T_1949 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@14563.4 package.scala 96:25:@14564.4]
  assign _T_1973 = _T_1949 ? Mem1D_5_io_output : _T_1972; // @[Mux.scala 31:69:@14618.4]
  assign _T_1946 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@14555.4 package.scala 96:25:@14556.4]
  assign _T_1974 = _T_1946 ? Mem1D_4_io_output : _T_1973; // @[Mux.scala 31:69:@14619.4]
  assign _T_1943 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@14547.4 package.scala 96:25:@14548.4]
  assign _T_1975 = _T_1943 ? Mem1D_3_io_output : _T_1974; // @[Mux.scala 31:69:@14620.4]
  assign _T_1940 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@14539.4 package.scala 96:25:@14540.4]
  assign _T_1976 = _T_1940 ? Mem1D_2_io_output : _T_1975; // @[Mux.scala 31:69:@14621.4]
  assign _T_1937 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@14531.4 package.scala 96:25:@14532.4]
  assign _T_1977 = _T_1937 ? Mem1D_1_io_output : _T_1976; // @[Mux.scala 31:69:@14622.4]
  assign _T_1934 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@14523.4 package.scala 96:25:@14524.4]
  assign _T_2071 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@14747.4 package.scala 96:25:@14748.4]
  assign _T_2075 = _T_2071 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14757.4]
  assign _T_2068 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@14739.4 package.scala 96:25:@14740.4]
  assign _T_2076 = _T_2068 ? Mem1D_9_io_output : _T_2075; // @[Mux.scala 31:69:@14758.4]
  assign _T_2065 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@14731.4 package.scala 96:25:@14732.4]
  assign _T_2077 = _T_2065 ? Mem1D_8_io_output : _T_2076; // @[Mux.scala 31:69:@14759.4]
  assign _T_2062 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@14723.4 package.scala 96:25:@14724.4]
  assign _T_2078 = _T_2062 ? Mem1D_7_io_output : _T_2077; // @[Mux.scala 31:69:@14760.4]
  assign _T_2059 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@14715.4 package.scala 96:25:@14716.4]
  assign _T_2079 = _T_2059 ? Mem1D_6_io_output : _T_2078; // @[Mux.scala 31:69:@14761.4]
  assign _T_2056 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@14707.4 package.scala 96:25:@14708.4]
  assign _T_2080 = _T_2056 ? Mem1D_5_io_output : _T_2079; // @[Mux.scala 31:69:@14762.4]
  assign _T_2053 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@14699.4 package.scala 96:25:@14700.4]
  assign _T_2081 = _T_2053 ? Mem1D_4_io_output : _T_2080; // @[Mux.scala 31:69:@14763.4]
  assign _T_2050 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@14691.4 package.scala 96:25:@14692.4]
  assign _T_2082 = _T_2050 ? Mem1D_3_io_output : _T_2081; // @[Mux.scala 31:69:@14764.4]
  assign _T_2047 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@14683.4 package.scala 96:25:@14684.4]
  assign _T_2083 = _T_2047 ? Mem1D_2_io_output : _T_2082; // @[Mux.scala 31:69:@14765.4]
  assign _T_2044 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@14675.4 package.scala 96:25:@14676.4]
  assign _T_2084 = _T_2044 ? Mem1D_1_io_output : _T_2083; // @[Mux.scala 31:69:@14766.4]
  assign _T_2041 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@14667.4 package.scala 96:25:@14668.4]
  assign _T_2178 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@14891.4 package.scala 96:25:@14892.4]
  assign _T_2182 = _T_2178 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@14901.4]
  assign _T_2175 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@14883.4 package.scala 96:25:@14884.4]
  assign _T_2183 = _T_2175 ? Mem1D_9_io_output : _T_2182; // @[Mux.scala 31:69:@14902.4]
  assign _T_2172 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@14875.4 package.scala 96:25:@14876.4]
  assign _T_2184 = _T_2172 ? Mem1D_8_io_output : _T_2183; // @[Mux.scala 31:69:@14903.4]
  assign _T_2169 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@14867.4 package.scala 96:25:@14868.4]
  assign _T_2185 = _T_2169 ? Mem1D_7_io_output : _T_2184; // @[Mux.scala 31:69:@14904.4]
  assign _T_2166 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@14859.4 package.scala 96:25:@14860.4]
  assign _T_2186 = _T_2166 ? Mem1D_6_io_output : _T_2185; // @[Mux.scala 31:69:@14905.4]
  assign _T_2163 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@14851.4 package.scala 96:25:@14852.4]
  assign _T_2187 = _T_2163 ? Mem1D_5_io_output : _T_2186; // @[Mux.scala 31:69:@14906.4]
  assign _T_2160 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@14843.4 package.scala 96:25:@14844.4]
  assign _T_2188 = _T_2160 ? Mem1D_4_io_output : _T_2187; // @[Mux.scala 31:69:@14907.4]
  assign _T_2157 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@14835.4 package.scala 96:25:@14836.4]
  assign _T_2189 = _T_2157 ? Mem1D_3_io_output : _T_2188; // @[Mux.scala 31:69:@14908.4]
  assign _T_2154 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@14827.4 package.scala 96:25:@14828.4]
  assign _T_2190 = _T_2154 ? Mem1D_2_io_output : _T_2189; // @[Mux.scala 31:69:@14909.4]
  assign _T_2151 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@14819.4 package.scala 96:25:@14820.4]
  assign _T_2191 = _T_2151 ? Mem1D_1_io_output : _T_2190; // @[Mux.scala 31:69:@14910.4]
  assign _T_2148 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@14811.4 package.scala 96:25:@14812.4]
  assign _T_2285 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@15035.4 package.scala 96:25:@15036.4]
  assign _T_2289 = _T_2285 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@15045.4]
  assign _T_2282 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@15027.4 package.scala 96:25:@15028.4]
  assign _T_2290 = _T_2282 ? Mem1D_9_io_output : _T_2289; // @[Mux.scala 31:69:@15046.4]
  assign _T_2279 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@15019.4 package.scala 96:25:@15020.4]
  assign _T_2291 = _T_2279 ? Mem1D_8_io_output : _T_2290; // @[Mux.scala 31:69:@15047.4]
  assign _T_2276 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@15011.4 package.scala 96:25:@15012.4]
  assign _T_2292 = _T_2276 ? Mem1D_7_io_output : _T_2291; // @[Mux.scala 31:69:@15048.4]
  assign _T_2273 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@15003.4 package.scala 96:25:@15004.4]
  assign _T_2293 = _T_2273 ? Mem1D_6_io_output : _T_2292; // @[Mux.scala 31:69:@15049.4]
  assign _T_2270 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@14995.4 package.scala 96:25:@14996.4]
  assign _T_2294 = _T_2270 ? Mem1D_5_io_output : _T_2293; // @[Mux.scala 31:69:@15050.4]
  assign _T_2267 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@14987.4 package.scala 96:25:@14988.4]
  assign _T_2295 = _T_2267 ? Mem1D_4_io_output : _T_2294; // @[Mux.scala 31:69:@15051.4]
  assign _T_2264 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@14979.4 package.scala 96:25:@14980.4]
  assign _T_2296 = _T_2264 ? Mem1D_3_io_output : _T_2295; // @[Mux.scala 31:69:@15052.4]
  assign _T_2261 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@14971.4 package.scala 96:25:@14972.4]
  assign _T_2297 = _T_2261 ? Mem1D_2_io_output : _T_2296; // @[Mux.scala 31:69:@15053.4]
  assign _T_2258 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@14963.4 package.scala 96:25:@14964.4]
  assign _T_2298 = _T_2258 ? Mem1D_1_io_output : _T_2297; // @[Mux.scala 31:69:@15054.4]
  assign _T_2255 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@14955.4 package.scala 96:25:@14956.4]
  assign _T_2392 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@15179.4 package.scala 96:25:@15180.4]
  assign _T_2396 = _T_2392 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@15189.4]
  assign _T_2389 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@15171.4 package.scala 96:25:@15172.4]
  assign _T_2397 = _T_2389 ? Mem1D_9_io_output : _T_2396; // @[Mux.scala 31:69:@15190.4]
  assign _T_2386 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@15163.4 package.scala 96:25:@15164.4]
  assign _T_2398 = _T_2386 ? Mem1D_8_io_output : _T_2397; // @[Mux.scala 31:69:@15191.4]
  assign _T_2383 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@15155.4 package.scala 96:25:@15156.4]
  assign _T_2399 = _T_2383 ? Mem1D_7_io_output : _T_2398; // @[Mux.scala 31:69:@15192.4]
  assign _T_2380 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@15147.4 package.scala 96:25:@15148.4]
  assign _T_2400 = _T_2380 ? Mem1D_6_io_output : _T_2399; // @[Mux.scala 31:69:@15193.4]
  assign _T_2377 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@15139.4 package.scala 96:25:@15140.4]
  assign _T_2401 = _T_2377 ? Mem1D_5_io_output : _T_2400; // @[Mux.scala 31:69:@15194.4]
  assign _T_2374 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@15131.4 package.scala 96:25:@15132.4]
  assign _T_2402 = _T_2374 ? Mem1D_4_io_output : _T_2401; // @[Mux.scala 31:69:@15195.4]
  assign _T_2371 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@15123.4 package.scala 96:25:@15124.4]
  assign _T_2403 = _T_2371 ? Mem1D_3_io_output : _T_2402; // @[Mux.scala 31:69:@15196.4]
  assign _T_2368 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@15115.4 package.scala 96:25:@15116.4]
  assign _T_2404 = _T_2368 ? Mem1D_2_io_output : _T_2403; // @[Mux.scala 31:69:@15197.4]
  assign _T_2365 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@15107.4 package.scala 96:25:@15108.4]
  assign _T_2405 = _T_2365 ? Mem1D_1_io_output : _T_2404; // @[Mux.scala 31:69:@15198.4]
  assign _T_2362 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@15099.4 package.scala 96:25:@15100.4]
  assign _T_2499 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@15323.4 package.scala 96:25:@15324.4]
  assign _T_2503 = _T_2499 ? Mem1D_10_io_output : Mem1D_11_io_output; // @[Mux.scala 31:69:@15333.4]
  assign _T_2496 = RetimeWrapper_105_io_out; // @[package.scala 96:25:@15315.4 package.scala 96:25:@15316.4]
  assign _T_2504 = _T_2496 ? Mem1D_9_io_output : _T_2503; // @[Mux.scala 31:69:@15334.4]
  assign _T_2493 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@15307.4 package.scala 96:25:@15308.4]
  assign _T_2505 = _T_2493 ? Mem1D_8_io_output : _T_2504; // @[Mux.scala 31:69:@15335.4]
  assign _T_2490 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@15299.4 package.scala 96:25:@15300.4]
  assign _T_2506 = _T_2490 ? Mem1D_7_io_output : _T_2505; // @[Mux.scala 31:69:@15336.4]
  assign _T_2487 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@15291.4 package.scala 96:25:@15292.4]
  assign _T_2507 = _T_2487 ? Mem1D_6_io_output : _T_2506; // @[Mux.scala 31:69:@15337.4]
  assign _T_2484 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@15283.4 package.scala 96:25:@15284.4]
  assign _T_2508 = _T_2484 ? Mem1D_5_io_output : _T_2507; // @[Mux.scala 31:69:@15338.4]
  assign _T_2481 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@15275.4 package.scala 96:25:@15276.4]
  assign _T_2509 = _T_2481 ? Mem1D_4_io_output : _T_2508; // @[Mux.scala 31:69:@15339.4]
  assign _T_2478 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@15267.4 package.scala 96:25:@15268.4]
  assign _T_2510 = _T_2478 ? Mem1D_3_io_output : _T_2509; // @[Mux.scala 31:69:@15340.4]
  assign _T_2475 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@15259.4 package.scala 96:25:@15260.4]
  assign _T_2511 = _T_2475 ? Mem1D_2_io_output : _T_2510; // @[Mux.scala 31:69:@15341.4]
  assign _T_2472 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@15251.4 package.scala 96:25:@15252.4]
  assign _T_2512 = _T_2472 ? Mem1D_1_io_output : _T_2511; // @[Mux.scala 31:69:@15342.4]
  assign _T_2469 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@15243.4 package.scala 96:25:@15244.4]
  assign io_rPort_8_output_0 = _T_2469 ? Mem1D_io_output : _T_2512; // @[MemPrimitives.scala 148:13:@15344.4]
  assign io_rPort_7_output_0 = _T_2362 ? Mem1D_io_output : _T_2405; // @[MemPrimitives.scala 148:13:@15200.4]
  assign io_rPort_6_output_0 = _T_2255 ? Mem1D_io_output : _T_2298; // @[MemPrimitives.scala 148:13:@15056.4]
  assign io_rPort_5_output_0 = _T_2148 ? Mem1D_io_output : _T_2191; // @[MemPrimitives.scala 148:13:@14912.4]
  assign io_rPort_4_output_0 = _T_2041 ? Mem1D_io_output : _T_2084; // @[MemPrimitives.scala 148:13:@14768.4]
  assign io_rPort_3_output_0 = _T_1934 ? Mem1D_io_output : _T_1977; // @[MemPrimitives.scala 148:13:@14624.4]
  assign io_rPort_2_output_0 = _T_1827 ? Mem1D_io_output : _T_1870; // @[MemPrimitives.scala 148:13:@14480.4]
  assign io_rPort_1_output_0 = _T_1720 ? Mem1D_io_output : _T_1763; // @[MemPrimitives.scala 148:13:@14336.4]
  assign io_rPort_0_output_0 = _T_1613 ? Mem1D_io_output : _T_1656; // @[MemPrimitives.scala 148:13:@14192.4]
  assign Mem1D_clock = clock; // @[:@12646.4]
  assign Mem1D_reset = reset; // @[:@12647.4]
  assign Mem1D_io_r_ofs_0 = _T_535[9:0]; // @[MemPrimitives.scala 127:28:@13067.4]
  assign Mem1D_io_r_backpressure = _T_535[10]; // @[MemPrimitives.scala 128:32:@13068.4]
  assign Mem1D_io_w_ofs_0 = _T_322[9:0]; // @[MemPrimitives.scala 94:28:@12846.4]
  assign Mem1D_io_w_data_0 = _T_322[17:10]; // @[MemPrimitives.scala 95:29:@12847.4]
  assign Mem1D_io_w_en_0 = _T_322[18]; // @[MemPrimitives.scala 96:27:@12848.4]
  assign Mem1D_1_clock = clock; // @[:@12662.4]
  assign Mem1D_1_reset = reset; // @[:@12663.4]
  assign Mem1D_1_io_r_ofs_0 = _T_627[9:0]; // @[MemPrimitives.scala 127:28:@13156.4]
  assign Mem1D_1_io_r_backpressure = _T_627[10]; // @[MemPrimitives.scala 128:32:@13157.4]
  assign Mem1D_1_io_w_ofs_0 = _T_333[9:0]; // @[MemPrimitives.scala 94:28:@12858.4]
  assign Mem1D_1_io_w_data_0 = _T_333[17:10]; // @[MemPrimitives.scala 95:29:@12859.4]
  assign Mem1D_1_io_w_en_0 = _T_333[18]; // @[MemPrimitives.scala 96:27:@12860.4]
  assign Mem1D_2_clock = clock; // @[:@12678.4]
  assign Mem1D_2_reset = reset; // @[:@12679.4]
  assign Mem1D_2_io_r_ofs_0 = _T_719[9:0]; // @[MemPrimitives.scala 127:28:@13245.4]
  assign Mem1D_2_io_r_backpressure = _T_719[10]; // @[MemPrimitives.scala 128:32:@13246.4]
  assign Mem1D_2_io_w_ofs_0 = _T_344[9:0]; // @[MemPrimitives.scala 94:28:@12870.4]
  assign Mem1D_2_io_w_data_0 = _T_344[17:10]; // @[MemPrimitives.scala 95:29:@12871.4]
  assign Mem1D_2_io_w_en_0 = _T_344[18]; // @[MemPrimitives.scala 96:27:@12872.4]
  assign Mem1D_3_clock = clock; // @[:@12694.4]
  assign Mem1D_3_reset = reset; // @[:@12695.4]
  assign Mem1D_3_io_r_ofs_0 = _T_811[9:0]; // @[MemPrimitives.scala 127:28:@13334.4]
  assign Mem1D_3_io_r_backpressure = _T_811[10]; // @[MemPrimitives.scala 128:32:@13335.4]
  assign Mem1D_3_io_w_ofs_0 = _T_355[9:0]; // @[MemPrimitives.scala 94:28:@12882.4]
  assign Mem1D_3_io_w_data_0 = _T_355[17:10]; // @[MemPrimitives.scala 95:29:@12883.4]
  assign Mem1D_3_io_w_en_0 = _T_355[18]; // @[MemPrimitives.scala 96:27:@12884.4]
  assign Mem1D_4_clock = clock; // @[:@12710.4]
  assign Mem1D_4_reset = reset; // @[:@12711.4]
  assign Mem1D_4_io_r_ofs_0 = _T_903[9:0]; // @[MemPrimitives.scala 127:28:@13423.4]
  assign Mem1D_4_io_r_backpressure = _T_903[10]; // @[MemPrimitives.scala 128:32:@13424.4]
  assign Mem1D_4_io_w_ofs_0 = _T_366[9:0]; // @[MemPrimitives.scala 94:28:@12894.4]
  assign Mem1D_4_io_w_data_0 = _T_366[17:10]; // @[MemPrimitives.scala 95:29:@12895.4]
  assign Mem1D_4_io_w_en_0 = _T_366[18]; // @[MemPrimitives.scala 96:27:@12896.4]
  assign Mem1D_5_clock = clock; // @[:@12726.4]
  assign Mem1D_5_reset = reset; // @[:@12727.4]
  assign Mem1D_5_io_r_ofs_0 = _T_995[9:0]; // @[MemPrimitives.scala 127:28:@13512.4]
  assign Mem1D_5_io_r_backpressure = _T_995[10]; // @[MemPrimitives.scala 128:32:@13513.4]
  assign Mem1D_5_io_w_ofs_0 = _T_377[9:0]; // @[MemPrimitives.scala 94:28:@12906.4]
  assign Mem1D_5_io_w_data_0 = _T_377[17:10]; // @[MemPrimitives.scala 95:29:@12907.4]
  assign Mem1D_5_io_w_en_0 = _T_377[18]; // @[MemPrimitives.scala 96:27:@12908.4]
  assign Mem1D_6_clock = clock; // @[:@12742.4]
  assign Mem1D_6_reset = reset; // @[:@12743.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1087[9:0]; // @[MemPrimitives.scala 127:28:@13601.4]
  assign Mem1D_6_io_r_backpressure = _T_1087[10]; // @[MemPrimitives.scala 128:32:@13602.4]
  assign Mem1D_6_io_w_ofs_0 = _T_388[9:0]; // @[MemPrimitives.scala 94:28:@12918.4]
  assign Mem1D_6_io_w_data_0 = _T_388[17:10]; // @[MemPrimitives.scala 95:29:@12919.4]
  assign Mem1D_6_io_w_en_0 = _T_388[18]; // @[MemPrimitives.scala 96:27:@12920.4]
  assign Mem1D_7_clock = clock; // @[:@12758.4]
  assign Mem1D_7_reset = reset; // @[:@12759.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1179[9:0]; // @[MemPrimitives.scala 127:28:@13690.4]
  assign Mem1D_7_io_r_backpressure = _T_1179[10]; // @[MemPrimitives.scala 128:32:@13691.4]
  assign Mem1D_7_io_w_ofs_0 = _T_399[9:0]; // @[MemPrimitives.scala 94:28:@12930.4]
  assign Mem1D_7_io_w_data_0 = _T_399[17:10]; // @[MemPrimitives.scala 95:29:@12931.4]
  assign Mem1D_7_io_w_en_0 = _T_399[18]; // @[MemPrimitives.scala 96:27:@12932.4]
  assign Mem1D_8_clock = clock; // @[:@12774.4]
  assign Mem1D_8_reset = reset; // @[:@12775.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1271[9:0]; // @[MemPrimitives.scala 127:28:@13779.4]
  assign Mem1D_8_io_r_backpressure = _T_1271[10]; // @[MemPrimitives.scala 128:32:@13780.4]
  assign Mem1D_8_io_w_ofs_0 = _T_410[9:0]; // @[MemPrimitives.scala 94:28:@12942.4]
  assign Mem1D_8_io_w_data_0 = _T_410[17:10]; // @[MemPrimitives.scala 95:29:@12943.4]
  assign Mem1D_8_io_w_en_0 = _T_410[18]; // @[MemPrimitives.scala 96:27:@12944.4]
  assign Mem1D_9_clock = clock; // @[:@12790.4]
  assign Mem1D_9_reset = reset; // @[:@12791.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1363[9:0]; // @[MemPrimitives.scala 127:28:@13868.4]
  assign Mem1D_9_io_r_backpressure = _T_1363[10]; // @[MemPrimitives.scala 128:32:@13869.4]
  assign Mem1D_9_io_w_ofs_0 = _T_421[9:0]; // @[MemPrimitives.scala 94:28:@12954.4]
  assign Mem1D_9_io_w_data_0 = _T_421[17:10]; // @[MemPrimitives.scala 95:29:@12955.4]
  assign Mem1D_9_io_w_en_0 = _T_421[18]; // @[MemPrimitives.scala 96:27:@12956.4]
  assign Mem1D_10_clock = clock; // @[:@12806.4]
  assign Mem1D_10_reset = reset; // @[:@12807.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1455[9:0]; // @[MemPrimitives.scala 127:28:@13957.4]
  assign Mem1D_10_io_r_backpressure = _T_1455[10]; // @[MemPrimitives.scala 128:32:@13958.4]
  assign Mem1D_10_io_w_ofs_0 = _T_432[9:0]; // @[MemPrimitives.scala 94:28:@12966.4]
  assign Mem1D_10_io_w_data_0 = _T_432[17:10]; // @[MemPrimitives.scala 95:29:@12967.4]
  assign Mem1D_10_io_w_en_0 = _T_432[18]; // @[MemPrimitives.scala 96:27:@12968.4]
  assign Mem1D_11_clock = clock; // @[:@12822.4]
  assign Mem1D_11_reset = reset; // @[:@12823.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1547[9:0]; // @[MemPrimitives.scala 127:28:@14046.4]
  assign Mem1D_11_io_r_backpressure = _T_1547[10]; // @[MemPrimitives.scala 128:32:@14047.4]
  assign Mem1D_11_io_w_ofs_0 = _T_443[9:0]; // @[MemPrimitives.scala 94:28:@12978.4]
  assign Mem1D_11_io_w_data_0 = _T_443[17:10]; // @[MemPrimitives.scala 95:29:@12979.4]
  assign Mem1D_11_io_w_en_0 = _T_443[18]; // @[MemPrimitives.scala 96:27:@12980.4]
  assign StickySelects_clock = clock; // @[:@13018.4]
  assign StickySelects_reset = reset; // @[:@13019.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_451; // @[MemPrimitives.scala 122:60:@13020.4]
  assign StickySelects_io_ins_1 = io_rPort_1_en_0 & _T_457; // @[MemPrimitives.scala 122:60:@13021.4]
  assign StickySelects_io_ins_2 = io_rPort_2_en_0 & _T_463; // @[MemPrimitives.scala 122:60:@13022.4]
  assign StickySelects_io_ins_3 = io_rPort_3_en_0 & _T_469; // @[MemPrimitives.scala 122:60:@13023.4]
  assign StickySelects_io_ins_4 = io_rPort_4_en_0 & _T_475; // @[MemPrimitives.scala 122:60:@13024.4]
  assign StickySelects_io_ins_5 = io_rPort_5_en_0 & _T_481; // @[MemPrimitives.scala 122:60:@13025.4]
  assign StickySelects_io_ins_6 = io_rPort_6_en_0 & _T_487; // @[MemPrimitives.scala 122:60:@13026.4]
  assign StickySelects_io_ins_7 = io_rPort_7_en_0 & _T_493; // @[MemPrimitives.scala 122:60:@13027.4]
  assign StickySelects_io_ins_8 = io_rPort_8_en_0 & _T_499; // @[MemPrimitives.scala 122:60:@13028.4]
  assign StickySelects_1_clock = clock; // @[:@13107.4]
  assign StickySelects_1_reset = reset; // @[:@13108.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_543; // @[MemPrimitives.scala 122:60:@13109.4]
  assign StickySelects_1_io_ins_1 = io_rPort_1_en_0 & _T_549; // @[MemPrimitives.scala 122:60:@13110.4]
  assign StickySelects_1_io_ins_2 = io_rPort_2_en_0 & _T_555; // @[MemPrimitives.scala 122:60:@13111.4]
  assign StickySelects_1_io_ins_3 = io_rPort_3_en_0 & _T_561; // @[MemPrimitives.scala 122:60:@13112.4]
  assign StickySelects_1_io_ins_4 = io_rPort_4_en_0 & _T_567; // @[MemPrimitives.scala 122:60:@13113.4]
  assign StickySelects_1_io_ins_5 = io_rPort_5_en_0 & _T_573; // @[MemPrimitives.scala 122:60:@13114.4]
  assign StickySelects_1_io_ins_6 = io_rPort_6_en_0 & _T_579; // @[MemPrimitives.scala 122:60:@13115.4]
  assign StickySelects_1_io_ins_7 = io_rPort_7_en_0 & _T_585; // @[MemPrimitives.scala 122:60:@13116.4]
  assign StickySelects_1_io_ins_8 = io_rPort_8_en_0 & _T_591; // @[MemPrimitives.scala 122:60:@13117.4]
  assign StickySelects_2_clock = clock; // @[:@13196.4]
  assign StickySelects_2_reset = reset; // @[:@13197.4]
  assign StickySelects_2_io_ins_0 = io_rPort_0_en_0 & _T_635; // @[MemPrimitives.scala 122:60:@13198.4]
  assign StickySelects_2_io_ins_1 = io_rPort_1_en_0 & _T_641; // @[MemPrimitives.scala 122:60:@13199.4]
  assign StickySelects_2_io_ins_2 = io_rPort_2_en_0 & _T_647; // @[MemPrimitives.scala 122:60:@13200.4]
  assign StickySelects_2_io_ins_3 = io_rPort_3_en_0 & _T_653; // @[MemPrimitives.scala 122:60:@13201.4]
  assign StickySelects_2_io_ins_4 = io_rPort_4_en_0 & _T_659; // @[MemPrimitives.scala 122:60:@13202.4]
  assign StickySelects_2_io_ins_5 = io_rPort_5_en_0 & _T_665; // @[MemPrimitives.scala 122:60:@13203.4]
  assign StickySelects_2_io_ins_6 = io_rPort_6_en_0 & _T_671; // @[MemPrimitives.scala 122:60:@13204.4]
  assign StickySelects_2_io_ins_7 = io_rPort_7_en_0 & _T_677; // @[MemPrimitives.scala 122:60:@13205.4]
  assign StickySelects_2_io_ins_8 = io_rPort_8_en_0 & _T_683; // @[MemPrimitives.scala 122:60:@13206.4]
  assign StickySelects_3_clock = clock; // @[:@13285.4]
  assign StickySelects_3_reset = reset; // @[:@13286.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_727; // @[MemPrimitives.scala 122:60:@13287.4]
  assign StickySelects_3_io_ins_1 = io_rPort_1_en_0 & _T_733; // @[MemPrimitives.scala 122:60:@13288.4]
  assign StickySelects_3_io_ins_2 = io_rPort_2_en_0 & _T_739; // @[MemPrimitives.scala 122:60:@13289.4]
  assign StickySelects_3_io_ins_3 = io_rPort_3_en_0 & _T_745; // @[MemPrimitives.scala 122:60:@13290.4]
  assign StickySelects_3_io_ins_4 = io_rPort_4_en_0 & _T_751; // @[MemPrimitives.scala 122:60:@13291.4]
  assign StickySelects_3_io_ins_5 = io_rPort_5_en_0 & _T_757; // @[MemPrimitives.scala 122:60:@13292.4]
  assign StickySelects_3_io_ins_6 = io_rPort_6_en_0 & _T_763; // @[MemPrimitives.scala 122:60:@13293.4]
  assign StickySelects_3_io_ins_7 = io_rPort_7_en_0 & _T_769; // @[MemPrimitives.scala 122:60:@13294.4]
  assign StickySelects_3_io_ins_8 = io_rPort_8_en_0 & _T_775; // @[MemPrimitives.scala 122:60:@13295.4]
  assign StickySelects_4_clock = clock; // @[:@13374.4]
  assign StickySelects_4_reset = reset; // @[:@13375.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_819; // @[MemPrimitives.scala 122:60:@13376.4]
  assign StickySelects_4_io_ins_1 = io_rPort_1_en_0 & _T_825; // @[MemPrimitives.scala 122:60:@13377.4]
  assign StickySelects_4_io_ins_2 = io_rPort_2_en_0 & _T_831; // @[MemPrimitives.scala 122:60:@13378.4]
  assign StickySelects_4_io_ins_3 = io_rPort_3_en_0 & _T_837; // @[MemPrimitives.scala 122:60:@13379.4]
  assign StickySelects_4_io_ins_4 = io_rPort_4_en_0 & _T_843; // @[MemPrimitives.scala 122:60:@13380.4]
  assign StickySelects_4_io_ins_5 = io_rPort_5_en_0 & _T_849; // @[MemPrimitives.scala 122:60:@13381.4]
  assign StickySelects_4_io_ins_6 = io_rPort_6_en_0 & _T_855; // @[MemPrimitives.scala 122:60:@13382.4]
  assign StickySelects_4_io_ins_7 = io_rPort_7_en_0 & _T_861; // @[MemPrimitives.scala 122:60:@13383.4]
  assign StickySelects_4_io_ins_8 = io_rPort_8_en_0 & _T_867; // @[MemPrimitives.scala 122:60:@13384.4]
  assign StickySelects_5_clock = clock; // @[:@13463.4]
  assign StickySelects_5_reset = reset; // @[:@13464.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_911; // @[MemPrimitives.scala 122:60:@13465.4]
  assign StickySelects_5_io_ins_1 = io_rPort_1_en_0 & _T_917; // @[MemPrimitives.scala 122:60:@13466.4]
  assign StickySelects_5_io_ins_2 = io_rPort_2_en_0 & _T_923; // @[MemPrimitives.scala 122:60:@13467.4]
  assign StickySelects_5_io_ins_3 = io_rPort_3_en_0 & _T_929; // @[MemPrimitives.scala 122:60:@13468.4]
  assign StickySelects_5_io_ins_4 = io_rPort_4_en_0 & _T_935; // @[MemPrimitives.scala 122:60:@13469.4]
  assign StickySelects_5_io_ins_5 = io_rPort_5_en_0 & _T_941; // @[MemPrimitives.scala 122:60:@13470.4]
  assign StickySelects_5_io_ins_6 = io_rPort_6_en_0 & _T_947; // @[MemPrimitives.scala 122:60:@13471.4]
  assign StickySelects_5_io_ins_7 = io_rPort_7_en_0 & _T_953; // @[MemPrimitives.scala 122:60:@13472.4]
  assign StickySelects_5_io_ins_8 = io_rPort_8_en_0 & _T_959; // @[MemPrimitives.scala 122:60:@13473.4]
  assign StickySelects_6_clock = clock; // @[:@13552.4]
  assign StickySelects_6_reset = reset; // @[:@13553.4]
  assign StickySelects_6_io_ins_0 = io_rPort_0_en_0 & _T_1003; // @[MemPrimitives.scala 122:60:@13554.4]
  assign StickySelects_6_io_ins_1 = io_rPort_1_en_0 & _T_1009; // @[MemPrimitives.scala 122:60:@13555.4]
  assign StickySelects_6_io_ins_2 = io_rPort_2_en_0 & _T_1015; // @[MemPrimitives.scala 122:60:@13556.4]
  assign StickySelects_6_io_ins_3 = io_rPort_3_en_0 & _T_1021; // @[MemPrimitives.scala 122:60:@13557.4]
  assign StickySelects_6_io_ins_4 = io_rPort_4_en_0 & _T_1027; // @[MemPrimitives.scala 122:60:@13558.4]
  assign StickySelects_6_io_ins_5 = io_rPort_5_en_0 & _T_1033; // @[MemPrimitives.scala 122:60:@13559.4]
  assign StickySelects_6_io_ins_6 = io_rPort_6_en_0 & _T_1039; // @[MemPrimitives.scala 122:60:@13560.4]
  assign StickySelects_6_io_ins_7 = io_rPort_7_en_0 & _T_1045; // @[MemPrimitives.scala 122:60:@13561.4]
  assign StickySelects_6_io_ins_8 = io_rPort_8_en_0 & _T_1051; // @[MemPrimitives.scala 122:60:@13562.4]
  assign StickySelects_7_clock = clock; // @[:@13641.4]
  assign StickySelects_7_reset = reset; // @[:@13642.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_1095; // @[MemPrimitives.scala 122:60:@13643.4]
  assign StickySelects_7_io_ins_1 = io_rPort_1_en_0 & _T_1101; // @[MemPrimitives.scala 122:60:@13644.4]
  assign StickySelects_7_io_ins_2 = io_rPort_2_en_0 & _T_1107; // @[MemPrimitives.scala 122:60:@13645.4]
  assign StickySelects_7_io_ins_3 = io_rPort_3_en_0 & _T_1113; // @[MemPrimitives.scala 122:60:@13646.4]
  assign StickySelects_7_io_ins_4 = io_rPort_4_en_0 & _T_1119; // @[MemPrimitives.scala 122:60:@13647.4]
  assign StickySelects_7_io_ins_5 = io_rPort_5_en_0 & _T_1125; // @[MemPrimitives.scala 122:60:@13648.4]
  assign StickySelects_7_io_ins_6 = io_rPort_6_en_0 & _T_1131; // @[MemPrimitives.scala 122:60:@13649.4]
  assign StickySelects_7_io_ins_7 = io_rPort_7_en_0 & _T_1137; // @[MemPrimitives.scala 122:60:@13650.4]
  assign StickySelects_7_io_ins_8 = io_rPort_8_en_0 & _T_1143; // @[MemPrimitives.scala 122:60:@13651.4]
  assign StickySelects_8_clock = clock; // @[:@13730.4]
  assign StickySelects_8_reset = reset; // @[:@13731.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_1187; // @[MemPrimitives.scala 122:60:@13732.4]
  assign StickySelects_8_io_ins_1 = io_rPort_1_en_0 & _T_1193; // @[MemPrimitives.scala 122:60:@13733.4]
  assign StickySelects_8_io_ins_2 = io_rPort_2_en_0 & _T_1199; // @[MemPrimitives.scala 122:60:@13734.4]
  assign StickySelects_8_io_ins_3 = io_rPort_3_en_0 & _T_1205; // @[MemPrimitives.scala 122:60:@13735.4]
  assign StickySelects_8_io_ins_4 = io_rPort_4_en_0 & _T_1211; // @[MemPrimitives.scala 122:60:@13736.4]
  assign StickySelects_8_io_ins_5 = io_rPort_5_en_0 & _T_1217; // @[MemPrimitives.scala 122:60:@13737.4]
  assign StickySelects_8_io_ins_6 = io_rPort_6_en_0 & _T_1223; // @[MemPrimitives.scala 122:60:@13738.4]
  assign StickySelects_8_io_ins_7 = io_rPort_7_en_0 & _T_1229; // @[MemPrimitives.scala 122:60:@13739.4]
  assign StickySelects_8_io_ins_8 = io_rPort_8_en_0 & _T_1235; // @[MemPrimitives.scala 122:60:@13740.4]
  assign StickySelects_9_clock = clock; // @[:@13819.4]
  assign StickySelects_9_reset = reset; // @[:@13820.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_1279; // @[MemPrimitives.scala 122:60:@13821.4]
  assign StickySelects_9_io_ins_1 = io_rPort_1_en_0 & _T_1285; // @[MemPrimitives.scala 122:60:@13822.4]
  assign StickySelects_9_io_ins_2 = io_rPort_2_en_0 & _T_1291; // @[MemPrimitives.scala 122:60:@13823.4]
  assign StickySelects_9_io_ins_3 = io_rPort_3_en_0 & _T_1297; // @[MemPrimitives.scala 122:60:@13824.4]
  assign StickySelects_9_io_ins_4 = io_rPort_4_en_0 & _T_1303; // @[MemPrimitives.scala 122:60:@13825.4]
  assign StickySelects_9_io_ins_5 = io_rPort_5_en_0 & _T_1309; // @[MemPrimitives.scala 122:60:@13826.4]
  assign StickySelects_9_io_ins_6 = io_rPort_6_en_0 & _T_1315; // @[MemPrimitives.scala 122:60:@13827.4]
  assign StickySelects_9_io_ins_7 = io_rPort_7_en_0 & _T_1321; // @[MemPrimitives.scala 122:60:@13828.4]
  assign StickySelects_9_io_ins_8 = io_rPort_8_en_0 & _T_1327; // @[MemPrimitives.scala 122:60:@13829.4]
  assign StickySelects_10_clock = clock; // @[:@13908.4]
  assign StickySelects_10_reset = reset; // @[:@13909.4]
  assign StickySelects_10_io_ins_0 = io_rPort_0_en_0 & _T_1371; // @[MemPrimitives.scala 122:60:@13910.4]
  assign StickySelects_10_io_ins_1 = io_rPort_1_en_0 & _T_1377; // @[MemPrimitives.scala 122:60:@13911.4]
  assign StickySelects_10_io_ins_2 = io_rPort_2_en_0 & _T_1383; // @[MemPrimitives.scala 122:60:@13912.4]
  assign StickySelects_10_io_ins_3 = io_rPort_3_en_0 & _T_1389; // @[MemPrimitives.scala 122:60:@13913.4]
  assign StickySelects_10_io_ins_4 = io_rPort_4_en_0 & _T_1395; // @[MemPrimitives.scala 122:60:@13914.4]
  assign StickySelects_10_io_ins_5 = io_rPort_5_en_0 & _T_1401; // @[MemPrimitives.scala 122:60:@13915.4]
  assign StickySelects_10_io_ins_6 = io_rPort_6_en_0 & _T_1407; // @[MemPrimitives.scala 122:60:@13916.4]
  assign StickySelects_10_io_ins_7 = io_rPort_7_en_0 & _T_1413; // @[MemPrimitives.scala 122:60:@13917.4]
  assign StickySelects_10_io_ins_8 = io_rPort_8_en_0 & _T_1419; // @[MemPrimitives.scala 122:60:@13918.4]
  assign StickySelects_11_clock = clock; // @[:@13997.4]
  assign StickySelects_11_reset = reset; // @[:@13998.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_1463; // @[MemPrimitives.scala 122:60:@13999.4]
  assign StickySelects_11_io_ins_1 = io_rPort_1_en_0 & _T_1469; // @[MemPrimitives.scala 122:60:@14000.4]
  assign StickySelects_11_io_ins_2 = io_rPort_2_en_0 & _T_1475; // @[MemPrimitives.scala 122:60:@14001.4]
  assign StickySelects_11_io_ins_3 = io_rPort_3_en_0 & _T_1481; // @[MemPrimitives.scala 122:60:@14002.4]
  assign StickySelects_11_io_ins_4 = io_rPort_4_en_0 & _T_1487; // @[MemPrimitives.scala 122:60:@14003.4]
  assign StickySelects_11_io_ins_5 = io_rPort_5_en_0 & _T_1493; // @[MemPrimitives.scala 122:60:@14004.4]
  assign StickySelects_11_io_ins_6 = io_rPort_6_en_0 & _T_1499; // @[MemPrimitives.scala 122:60:@14005.4]
  assign StickySelects_11_io_ins_7 = io_rPort_7_en_0 & _T_1505; // @[MemPrimitives.scala 122:60:@14006.4]
  assign StickySelects_11_io_ins_8 = io_rPort_8_en_0 & _T_1511; // @[MemPrimitives.scala 122:60:@14007.4]
  assign RetimeWrapper_clock = clock; // @[:@14087.4]
  assign RetimeWrapper_reset = reset; // @[:@14088.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14090.4]
  assign RetimeWrapper_io_in = _T_451 & io_rPort_0_en_0; // @[package.scala 94:16:@14089.4]
  assign RetimeWrapper_1_clock = clock; // @[:@14095.4]
  assign RetimeWrapper_1_reset = reset; // @[:@14096.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14098.4]
  assign RetimeWrapper_1_io_in = _T_543 & io_rPort_0_en_0; // @[package.scala 94:16:@14097.4]
  assign RetimeWrapper_2_clock = clock; // @[:@14103.4]
  assign RetimeWrapper_2_reset = reset; // @[:@14104.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14106.4]
  assign RetimeWrapper_2_io_in = _T_635 & io_rPort_0_en_0; // @[package.scala 94:16:@14105.4]
  assign RetimeWrapper_3_clock = clock; // @[:@14111.4]
  assign RetimeWrapper_3_reset = reset; // @[:@14112.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14114.4]
  assign RetimeWrapper_3_io_in = _T_727 & io_rPort_0_en_0; // @[package.scala 94:16:@14113.4]
  assign RetimeWrapper_4_clock = clock; // @[:@14119.4]
  assign RetimeWrapper_4_reset = reset; // @[:@14120.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14122.4]
  assign RetimeWrapper_4_io_in = _T_819 & io_rPort_0_en_0; // @[package.scala 94:16:@14121.4]
  assign RetimeWrapper_5_clock = clock; // @[:@14127.4]
  assign RetimeWrapper_5_reset = reset; // @[:@14128.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14130.4]
  assign RetimeWrapper_5_io_in = _T_911 & io_rPort_0_en_0; // @[package.scala 94:16:@14129.4]
  assign RetimeWrapper_6_clock = clock; // @[:@14135.4]
  assign RetimeWrapper_6_reset = reset; // @[:@14136.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14138.4]
  assign RetimeWrapper_6_io_in = _T_1003 & io_rPort_0_en_0; // @[package.scala 94:16:@14137.4]
  assign RetimeWrapper_7_clock = clock; // @[:@14143.4]
  assign RetimeWrapper_7_reset = reset; // @[:@14144.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14146.4]
  assign RetimeWrapper_7_io_in = _T_1095 & io_rPort_0_en_0; // @[package.scala 94:16:@14145.4]
  assign RetimeWrapper_8_clock = clock; // @[:@14151.4]
  assign RetimeWrapper_8_reset = reset; // @[:@14152.4]
  assign RetimeWrapper_8_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14154.4]
  assign RetimeWrapper_8_io_in = _T_1187 & io_rPort_0_en_0; // @[package.scala 94:16:@14153.4]
  assign RetimeWrapper_9_clock = clock; // @[:@14159.4]
  assign RetimeWrapper_9_reset = reset; // @[:@14160.4]
  assign RetimeWrapper_9_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14162.4]
  assign RetimeWrapper_9_io_in = _T_1279 & io_rPort_0_en_0; // @[package.scala 94:16:@14161.4]
  assign RetimeWrapper_10_clock = clock; // @[:@14167.4]
  assign RetimeWrapper_10_reset = reset; // @[:@14168.4]
  assign RetimeWrapper_10_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14170.4]
  assign RetimeWrapper_10_io_in = _T_1371 & io_rPort_0_en_0; // @[package.scala 94:16:@14169.4]
  assign RetimeWrapper_11_clock = clock; // @[:@14175.4]
  assign RetimeWrapper_11_reset = reset; // @[:@14176.4]
  assign RetimeWrapper_11_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14178.4]
  assign RetimeWrapper_11_io_in = _T_1463 & io_rPort_0_en_0; // @[package.scala 94:16:@14177.4]
  assign RetimeWrapper_12_clock = clock; // @[:@14231.4]
  assign RetimeWrapper_12_reset = reset; // @[:@14232.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14234.4]
  assign RetimeWrapper_12_io_in = _T_457 & io_rPort_1_en_0; // @[package.scala 94:16:@14233.4]
  assign RetimeWrapper_13_clock = clock; // @[:@14239.4]
  assign RetimeWrapper_13_reset = reset; // @[:@14240.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14242.4]
  assign RetimeWrapper_13_io_in = _T_549 & io_rPort_1_en_0; // @[package.scala 94:16:@14241.4]
  assign RetimeWrapper_14_clock = clock; // @[:@14247.4]
  assign RetimeWrapper_14_reset = reset; // @[:@14248.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14250.4]
  assign RetimeWrapper_14_io_in = _T_641 & io_rPort_1_en_0; // @[package.scala 94:16:@14249.4]
  assign RetimeWrapper_15_clock = clock; // @[:@14255.4]
  assign RetimeWrapper_15_reset = reset; // @[:@14256.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14258.4]
  assign RetimeWrapper_15_io_in = _T_733 & io_rPort_1_en_0; // @[package.scala 94:16:@14257.4]
  assign RetimeWrapper_16_clock = clock; // @[:@14263.4]
  assign RetimeWrapper_16_reset = reset; // @[:@14264.4]
  assign RetimeWrapper_16_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14266.4]
  assign RetimeWrapper_16_io_in = _T_825 & io_rPort_1_en_0; // @[package.scala 94:16:@14265.4]
  assign RetimeWrapper_17_clock = clock; // @[:@14271.4]
  assign RetimeWrapper_17_reset = reset; // @[:@14272.4]
  assign RetimeWrapper_17_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14274.4]
  assign RetimeWrapper_17_io_in = _T_917 & io_rPort_1_en_0; // @[package.scala 94:16:@14273.4]
  assign RetimeWrapper_18_clock = clock; // @[:@14279.4]
  assign RetimeWrapper_18_reset = reset; // @[:@14280.4]
  assign RetimeWrapper_18_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14282.4]
  assign RetimeWrapper_18_io_in = _T_1009 & io_rPort_1_en_0; // @[package.scala 94:16:@14281.4]
  assign RetimeWrapper_19_clock = clock; // @[:@14287.4]
  assign RetimeWrapper_19_reset = reset; // @[:@14288.4]
  assign RetimeWrapper_19_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14290.4]
  assign RetimeWrapper_19_io_in = _T_1101 & io_rPort_1_en_0; // @[package.scala 94:16:@14289.4]
  assign RetimeWrapper_20_clock = clock; // @[:@14295.4]
  assign RetimeWrapper_20_reset = reset; // @[:@14296.4]
  assign RetimeWrapper_20_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14298.4]
  assign RetimeWrapper_20_io_in = _T_1193 & io_rPort_1_en_0; // @[package.scala 94:16:@14297.4]
  assign RetimeWrapper_21_clock = clock; // @[:@14303.4]
  assign RetimeWrapper_21_reset = reset; // @[:@14304.4]
  assign RetimeWrapper_21_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14306.4]
  assign RetimeWrapper_21_io_in = _T_1285 & io_rPort_1_en_0; // @[package.scala 94:16:@14305.4]
  assign RetimeWrapper_22_clock = clock; // @[:@14311.4]
  assign RetimeWrapper_22_reset = reset; // @[:@14312.4]
  assign RetimeWrapper_22_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14314.4]
  assign RetimeWrapper_22_io_in = _T_1377 & io_rPort_1_en_0; // @[package.scala 94:16:@14313.4]
  assign RetimeWrapper_23_clock = clock; // @[:@14319.4]
  assign RetimeWrapper_23_reset = reset; // @[:@14320.4]
  assign RetimeWrapper_23_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14322.4]
  assign RetimeWrapper_23_io_in = _T_1469 & io_rPort_1_en_0; // @[package.scala 94:16:@14321.4]
  assign RetimeWrapper_24_clock = clock; // @[:@14375.4]
  assign RetimeWrapper_24_reset = reset; // @[:@14376.4]
  assign RetimeWrapper_24_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14378.4]
  assign RetimeWrapper_24_io_in = _T_463 & io_rPort_2_en_0; // @[package.scala 94:16:@14377.4]
  assign RetimeWrapper_25_clock = clock; // @[:@14383.4]
  assign RetimeWrapper_25_reset = reset; // @[:@14384.4]
  assign RetimeWrapper_25_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14386.4]
  assign RetimeWrapper_25_io_in = _T_555 & io_rPort_2_en_0; // @[package.scala 94:16:@14385.4]
  assign RetimeWrapper_26_clock = clock; // @[:@14391.4]
  assign RetimeWrapper_26_reset = reset; // @[:@14392.4]
  assign RetimeWrapper_26_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14394.4]
  assign RetimeWrapper_26_io_in = _T_647 & io_rPort_2_en_0; // @[package.scala 94:16:@14393.4]
  assign RetimeWrapper_27_clock = clock; // @[:@14399.4]
  assign RetimeWrapper_27_reset = reset; // @[:@14400.4]
  assign RetimeWrapper_27_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14402.4]
  assign RetimeWrapper_27_io_in = _T_739 & io_rPort_2_en_0; // @[package.scala 94:16:@14401.4]
  assign RetimeWrapper_28_clock = clock; // @[:@14407.4]
  assign RetimeWrapper_28_reset = reset; // @[:@14408.4]
  assign RetimeWrapper_28_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14410.4]
  assign RetimeWrapper_28_io_in = _T_831 & io_rPort_2_en_0; // @[package.scala 94:16:@14409.4]
  assign RetimeWrapper_29_clock = clock; // @[:@14415.4]
  assign RetimeWrapper_29_reset = reset; // @[:@14416.4]
  assign RetimeWrapper_29_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14418.4]
  assign RetimeWrapper_29_io_in = _T_923 & io_rPort_2_en_0; // @[package.scala 94:16:@14417.4]
  assign RetimeWrapper_30_clock = clock; // @[:@14423.4]
  assign RetimeWrapper_30_reset = reset; // @[:@14424.4]
  assign RetimeWrapper_30_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14426.4]
  assign RetimeWrapper_30_io_in = _T_1015 & io_rPort_2_en_0; // @[package.scala 94:16:@14425.4]
  assign RetimeWrapper_31_clock = clock; // @[:@14431.4]
  assign RetimeWrapper_31_reset = reset; // @[:@14432.4]
  assign RetimeWrapper_31_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14434.4]
  assign RetimeWrapper_31_io_in = _T_1107 & io_rPort_2_en_0; // @[package.scala 94:16:@14433.4]
  assign RetimeWrapper_32_clock = clock; // @[:@14439.4]
  assign RetimeWrapper_32_reset = reset; // @[:@14440.4]
  assign RetimeWrapper_32_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14442.4]
  assign RetimeWrapper_32_io_in = _T_1199 & io_rPort_2_en_0; // @[package.scala 94:16:@14441.4]
  assign RetimeWrapper_33_clock = clock; // @[:@14447.4]
  assign RetimeWrapper_33_reset = reset; // @[:@14448.4]
  assign RetimeWrapper_33_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14450.4]
  assign RetimeWrapper_33_io_in = _T_1291 & io_rPort_2_en_0; // @[package.scala 94:16:@14449.4]
  assign RetimeWrapper_34_clock = clock; // @[:@14455.4]
  assign RetimeWrapper_34_reset = reset; // @[:@14456.4]
  assign RetimeWrapper_34_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14458.4]
  assign RetimeWrapper_34_io_in = _T_1383 & io_rPort_2_en_0; // @[package.scala 94:16:@14457.4]
  assign RetimeWrapper_35_clock = clock; // @[:@14463.4]
  assign RetimeWrapper_35_reset = reset; // @[:@14464.4]
  assign RetimeWrapper_35_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14466.4]
  assign RetimeWrapper_35_io_in = _T_1475 & io_rPort_2_en_0; // @[package.scala 94:16:@14465.4]
  assign RetimeWrapper_36_clock = clock; // @[:@14519.4]
  assign RetimeWrapper_36_reset = reset; // @[:@14520.4]
  assign RetimeWrapper_36_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14522.4]
  assign RetimeWrapper_36_io_in = _T_469 & io_rPort_3_en_0; // @[package.scala 94:16:@14521.4]
  assign RetimeWrapper_37_clock = clock; // @[:@14527.4]
  assign RetimeWrapper_37_reset = reset; // @[:@14528.4]
  assign RetimeWrapper_37_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14530.4]
  assign RetimeWrapper_37_io_in = _T_561 & io_rPort_3_en_0; // @[package.scala 94:16:@14529.4]
  assign RetimeWrapper_38_clock = clock; // @[:@14535.4]
  assign RetimeWrapper_38_reset = reset; // @[:@14536.4]
  assign RetimeWrapper_38_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14538.4]
  assign RetimeWrapper_38_io_in = _T_653 & io_rPort_3_en_0; // @[package.scala 94:16:@14537.4]
  assign RetimeWrapper_39_clock = clock; // @[:@14543.4]
  assign RetimeWrapper_39_reset = reset; // @[:@14544.4]
  assign RetimeWrapper_39_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14546.4]
  assign RetimeWrapper_39_io_in = _T_745 & io_rPort_3_en_0; // @[package.scala 94:16:@14545.4]
  assign RetimeWrapper_40_clock = clock; // @[:@14551.4]
  assign RetimeWrapper_40_reset = reset; // @[:@14552.4]
  assign RetimeWrapper_40_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14554.4]
  assign RetimeWrapper_40_io_in = _T_837 & io_rPort_3_en_0; // @[package.scala 94:16:@14553.4]
  assign RetimeWrapper_41_clock = clock; // @[:@14559.4]
  assign RetimeWrapper_41_reset = reset; // @[:@14560.4]
  assign RetimeWrapper_41_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14562.4]
  assign RetimeWrapper_41_io_in = _T_929 & io_rPort_3_en_0; // @[package.scala 94:16:@14561.4]
  assign RetimeWrapper_42_clock = clock; // @[:@14567.4]
  assign RetimeWrapper_42_reset = reset; // @[:@14568.4]
  assign RetimeWrapper_42_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14570.4]
  assign RetimeWrapper_42_io_in = _T_1021 & io_rPort_3_en_0; // @[package.scala 94:16:@14569.4]
  assign RetimeWrapper_43_clock = clock; // @[:@14575.4]
  assign RetimeWrapper_43_reset = reset; // @[:@14576.4]
  assign RetimeWrapper_43_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14578.4]
  assign RetimeWrapper_43_io_in = _T_1113 & io_rPort_3_en_0; // @[package.scala 94:16:@14577.4]
  assign RetimeWrapper_44_clock = clock; // @[:@14583.4]
  assign RetimeWrapper_44_reset = reset; // @[:@14584.4]
  assign RetimeWrapper_44_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14586.4]
  assign RetimeWrapper_44_io_in = _T_1205 & io_rPort_3_en_0; // @[package.scala 94:16:@14585.4]
  assign RetimeWrapper_45_clock = clock; // @[:@14591.4]
  assign RetimeWrapper_45_reset = reset; // @[:@14592.4]
  assign RetimeWrapper_45_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14594.4]
  assign RetimeWrapper_45_io_in = _T_1297 & io_rPort_3_en_0; // @[package.scala 94:16:@14593.4]
  assign RetimeWrapper_46_clock = clock; // @[:@14599.4]
  assign RetimeWrapper_46_reset = reset; // @[:@14600.4]
  assign RetimeWrapper_46_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14602.4]
  assign RetimeWrapper_46_io_in = _T_1389 & io_rPort_3_en_0; // @[package.scala 94:16:@14601.4]
  assign RetimeWrapper_47_clock = clock; // @[:@14607.4]
  assign RetimeWrapper_47_reset = reset; // @[:@14608.4]
  assign RetimeWrapper_47_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14610.4]
  assign RetimeWrapper_47_io_in = _T_1481 & io_rPort_3_en_0; // @[package.scala 94:16:@14609.4]
  assign RetimeWrapper_48_clock = clock; // @[:@14663.4]
  assign RetimeWrapper_48_reset = reset; // @[:@14664.4]
  assign RetimeWrapper_48_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14666.4]
  assign RetimeWrapper_48_io_in = _T_475 & io_rPort_4_en_0; // @[package.scala 94:16:@14665.4]
  assign RetimeWrapper_49_clock = clock; // @[:@14671.4]
  assign RetimeWrapper_49_reset = reset; // @[:@14672.4]
  assign RetimeWrapper_49_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14674.4]
  assign RetimeWrapper_49_io_in = _T_567 & io_rPort_4_en_0; // @[package.scala 94:16:@14673.4]
  assign RetimeWrapper_50_clock = clock; // @[:@14679.4]
  assign RetimeWrapper_50_reset = reset; // @[:@14680.4]
  assign RetimeWrapper_50_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14682.4]
  assign RetimeWrapper_50_io_in = _T_659 & io_rPort_4_en_0; // @[package.scala 94:16:@14681.4]
  assign RetimeWrapper_51_clock = clock; // @[:@14687.4]
  assign RetimeWrapper_51_reset = reset; // @[:@14688.4]
  assign RetimeWrapper_51_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14690.4]
  assign RetimeWrapper_51_io_in = _T_751 & io_rPort_4_en_0; // @[package.scala 94:16:@14689.4]
  assign RetimeWrapper_52_clock = clock; // @[:@14695.4]
  assign RetimeWrapper_52_reset = reset; // @[:@14696.4]
  assign RetimeWrapper_52_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14698.4]
  assign RetimeWrapper_52_io_in = _T_843 & io_rPort_4_en_0; // @[package.scala 94:16:@14697.4]
  assign RetimeWrapper_53_clock = clock; // @[:@14703.4]
  assign RetimeWrapper_53_reset = reset; // @[:@14704.4]
  assign RetimeWrapper_53_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14706.4]
  assign RetimeWrapper_53_io_in = _T_935 & io_rPort_4_en_0; // @[package.scala 94:16:@14705.4]
  assign RetimeWrapper_54_clock = clock; // @[:@14711.4]
  assign RetimeWrapper_54_reset = reset; // @[:@14712.4]
  assign RetimeWrapper_54_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14714.4]
  assign RetimeWrapper_54_io_in = _T_1027 & io_rPort_4_en_0; // @[package.scala 94:16:@14713.4]
  assign RetimeWrapper_55_clock = clock; // @[:@14719.4]
  assign RetimeWrapper_55_reset = reset; // @[:@14720.4]
  assign RetimeWrapper_55_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14722.4]
  assign RetimeWrapper_55_io_in = _T_1119 & io_rPort_4_en_0; // @[package.scala 94:16:@14721.4]
  assign RetimeWrapper_56_clock = clock; // @[:@14727.4]
  assign RetimeWrapper_56_reset = reset; // @[:@14728.4]
  assign RetimeWrapper_56_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14730.4]
  assign RetimeWrapper_56_io_in = _T_1211 & io_rPort_4_en_0; // @[package.scala 94:16:@14729.4]
  assign RetimeWrapper_57_clock = clock; // @[:@14735.4]
  assign RetimeWrapper_57_reset = reset; // @[:@14736.4]
  assign RetimeWrapper_57_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14738.4]
  assign RetimeWrapper_57_io_in = _T_1303 & io_rPort_4_en_0; // @[package.scala 94:16:@14737.4]
  assign RetimeWrapper_58_clock = clock; // @[:@14743.4]
  assign RetimeWrapper_58_reset = reset; // @[:@14744.4]
  assign RetimeWrapper_58_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14746.4]
  assign RetimeWrapper_58_io_in = _T_1395 & io_rPort_4_en_0; // @[package.scala 94:16:@14745.4]
  assign RetimeWrapper_59_clock = clock; // @[:@14751.4]
  assign RetimeWrapper_59_reset = reset; // @[:@14752.4]
  assign RetimeWrapper_59_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14754.4]
  assign RetimeWrapper_59_io_in = _T_1487 & io_rPort_4_en_0; // @[package.scala 94:16:@14753.4]
  assign RetimeWrapper_60_clock = clock; // @[:@14807.4]
  assign RetimeWrapper_60_reset = reset; // @[:@14808.4]
  assign RetimeWrapper_60_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14810.4]
  assign RetimeWrapper_60_io_in = _T_481 & io_rPort_5_en_0; // @[package.scala 94:16:@14809.4]
  assign RetimeWrapper_61_clock = clock; // @[:@14815.4]
  assign RetimeWrapper_61_reset = reset; // @[:@14816.4]
  assign RetimeWrapper_61_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14818.4]
  assign RetimeWrapper_61_io_in = _T_573 & io_rPort_5_en_0; // @[package.scala 94:16:@14817.4]
  assign RetimeWrapper_62_clock = clock; // @[:@14823.4]
  assign RetimeWrapper_62_reset = reset; // @[:@14824.4]
  assign RetimeWrapper_62_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14826.4]
  assign RetimeWrapper_62_io_in = _T_665 & io_rPort_5_en_0; // @[package.scala 94:16:@14825.4]
  assign RetimeWrapper_63_clock = clock; // @[:@14831.4]
  assign RetimeWrapper_63_reset = reset; // @[:@14832.4]
  assign RetimeWrapper_63_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14834.4]
  assign RetimeWrapper_63_io_in = _T_757 & io_rPort_5_en_0; // @[package.scala 94:16:@14833.4]
  assign RetimeWrapper_64_clock = clock; // @[:@14839.4]
  assign RetimeWrapper_64_reset = reset; // @[:@14840.4]
  assign RetimeWrapper_64_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14842.4]
  assign RetimeWrapper_64_io_in = _T_849 & io_rPort_5_en_0; // @[package.scala 94:16:@14841.4]
  assign RetimeWrapper_65_clock = clock; // @[:@14847.4]
  assign RetimeWrapper_65_reset = reset; // @[:@14848.4]
  assign RetimeWrapper_65_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14850.4]
  assign RetimeWrapper_65_io_in = _T_941 & io_rPort_5_en_0; // @[package.scala 94:16:@14849.4]
  assign RetimeWrapper_66_clock = clock; // @[:@14855.4]
  assign RetimeWrapper_66_reset = reset; // @[:@14856.4]
  assign RetimeWrapper_66_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14858.4]
  assign RetimeWrapper_66_io_in = _T_1033 & io_rPort_5_en_0; // @[package.scala 94:16:@14857.4]
  assign RetimeWrapper_67_clock = clock; // @[:@14863.4]
  assign RetimeWrapper_67_reset = reset; // @[:@14864.4]
  assign RetimeWrapper_67_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14866.4]
  assign RetimeWrapper_67_io_in = _T_1125 & io_rPort_5_en_0; // @[package.scala 94:16:@14865.4]
  assign RetimeWrapper_68_clock = clock; // @[:@14871.4]
  assign RetimeWrapper_68_reset = reset; // @[:@14872.4]
  assign RetimeWrapper_68_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14874.4]
  assign RetimeWrapper_68_io_in = _T_1217 & io_rPort_5_en_0; // @[package.scala 94:16:@14873.4]
  assign RetimeWrapper_69_clock = clock; // @[:@14879.4]
  assign RetimeWrapper_69_reset = reset; // @[:@14880.4]
  assign RetimeWrapper_69_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14882.4]
  assign RetimeWrapper_69_io_in = _T_1309 & io_rPort_5_en_0; // @[package.scala 94:16:@14881.4]
  assign RetimeWrapper_70_clock = clock; // @[:@14887.4]
  assign RetimeWrapper_70_reset = reset; // @[:@14888.4]
  assign RetimeWrapper_70_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14890.4]
  assign RetimeWrapper_70_io_in = _T_1401 & io_rPort_5_en_0; // @[package.scala 94:16:@14889.4]
  assign RetimeWrapper_71_clock = clock; // @[:@14895.4]
  assign RetimeWrapper_71_reset = reset; // @[:@14896.4]
  assign RetimeWrapper_71_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14898.4]
  assign RetimeWrapper_71_io_in = _T_1493 & io_rPort_5_en_0; // @[package.scala 94:16:@14897.4]
  assign RetimeWrapper_72_clock = clock; // @[:@14951.4]
  assign RetimeWrapper_72_reset = reset; // @[:@14952.4]
  assign RetimeWrapper_72_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14954.4]
  assign RetimeWrapper_72_io_in = _T_487 & io_rPort_6_en_0; // @[package.scala 94:16:@14953.4]
  assign RetimeWrapper_73_clock = clock; // @[:@14959.4]
  assign RetimeWrapper_73_reset = reset; // @[:@14960.4]
  assign RetimeWrapper_73_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14962.4]
  assign RetimeWrapper_73_io_in = _T_579 & io_rPort_6_en_0; // @[package.scala 94:16:@14961.4]
  assign RetimeWrapper_74_clock = clock; // @[:@14967.4]
  assign RetimeWrapper_74_reset = reset; // @[:@14968.4]
  assign RetimeWrapper_74_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14970.4]
  assign RetimeWrapper_74_io_in = _T_671 & io_rPort_6_en_0; // @[package.scala 94:16:@14969.4]
  assign RetimeWrapper_75_clock = clock; // @[:@14975.4]
  assign RetimeWrapper_75_reset = reset; // @[:@14976.4]
  assign RetimeWrapper_75_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14978.4]
  assign RetimeWrapper_75_io_in = _T_763 & io_rPort_6_en_0; // @[package.scala 94:16:@14977.4]
  assign RetimeWrapper_76_clock = clock; // @[:@14983.4]
  assign RetimeWrapper_76_reset = reset; // @[:@14984.4]
  assign RetimeWrapper_76_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14986.4]
  assign RetimeWrapper_76_io_in = _T_855 & io_rPort_6_en_0; // @[package.scala 94:16:@14985.4]
  assign RetimeWrapper_77_clock = clock; // @[:@14991.4]
  assign RetimeWrapper_77_reset = reset; // @[:@14992.4]
  assign RetimeWrapper_77_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14994.4]
  assign RetimeWrapper_77_io_in = _T_947 & io_rPort_6_en_0; // @[package.scala 94:16:@14993.4]
  assign RetimeWrapper_78_clock = clock; // @[:@14999.4]
  assign RetimeWrapper_78_reset = reset; // @[:@15000.4]
  assign RetimeWrapper_78_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15002.4]
  assign RetimeWrapper_78_io_in = _T_1039 & io_rPort_6_en_0; // @[package.scala 94:16:@15001.4]
  assign RetimeWrapper_79_clock = clock; // @[:@15007.4]
  assign RetimeWrapper_79_reset = reset; // @[:@15008.4]
  assign RetimeWrapper_79_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15010.4]
  assign RetimeWrapper_79_io_in = _T_1131 & io_rPort_6_en_0; // @[package.scala 94:16:@15009.4]
  assign RetimeWrapper_80_clock = clock; // @[:@15015.4]
  assign RetimeWrapper_80_reset = reset; // @[:@15016.4]
  assign RetimeWrapper_80_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15018.4]
  assign RetimeWrapper_80_io_in = _T_1223 & io_rPort_6_en_0; // @[package.scala 94:16:@15017.4]
  assign RetimeWrapper_81_clock = clock; // @[:@15023.4]
  assign RetimeWrapper_81_reset = reset; // @[:@15024.4]
  assign RetimeWrapper_81_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15026.4]
  assign RetimeWrapper_81_io_in = _T_1315 & io_rPort_6_en_0; // @[package.scala 94:16:@15025.4]
  assign RetimeWrapper_82_clock = clock; // @[:@15031.4]
  assign RetimeWrapper_82_reset = reset; // @[:@15032.4]
  assign RetimeWrapper_82_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15034.4]
  assign RetimeWrapper_82_io_in = _T_1407 & io_rPort_6_en_0; // @[package.scala 94:16:@15033.4]
  assign RetimeWrapper_83_clock = clock; // @[:@15039.4]
  assign RetimeWrapper_83_reset = reset; // @[:@15040.4]
  assign RetimeWrapper_83_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@15042.4]
  assign RetimeWrapper_83_io_in = _T_1499 & io_rPort_6_en_0; // @[package.scala 94:16:@15041.4]
  assign RetimeWrapper_84_clock = clock; // @[:@15095.4]
  assign RetimeWrapper_84_reset = reset; // @[:@15096.4]
  assign RetimeWrapper_84_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15098.4]
  assign RetimeWrapper_84_io_in = _T_493 & io_rPort_7_en_0; // @[package.scala 94:16:@15097.4]
  assign RetimeWrapper_85_clock = clock; // @[:@15103.4]
  assign RetimeWrapper_85_reset = reset; // @[:@15104.4]
  assign RetimeWrapper_85_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15106.4]
  assign RetimeWrapper_85_io_in = _T_585 & io_rPort_7_en_0; // @[package.scala 94:16:@15105.4]
  assign RetimeWrapper_86_clock = clock; // @[:@15111.4]
  assign RetimeWrapper_86_reset = reset; // @[:@15112.4]
  assign RetimeWrapper_86_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15114.4]
  assign RetimeWrapper_86_io_in = _T_677 & io_rPort_7_en_0; // @[package.scala 94:16:@15113.4]
  assign RetimeWrapper_87_clock = clock; // @[:@15119.4]
  assign RetimeWrapper_87_reset = reset; // @[:@15120.4]
  assign RetimeWrapper_87_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15122.4]
  assign RetimeWrapper_87_io_in = _T_769 & io_rPort_7_en_0; // @[package.scala 94:16:@15121.4]
  assign RetimeWrapper_88_clock = clock; // @[:@15127.4]
  assign RetimeWrapper_88_reset = reset; // @[:@15128.4]
  assign RetimeWrapper_88_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15130.4]
  assign RetimeWrapper_88_io_in = _T_861 & io_rPort_7_en_0; // @[package.scala 94:16:@15129.4]
  assign RetimeWrapper_89_clock = clock; // @[:@15135.4]
  assign RetimeWrapper_89_reset = reset; // @[:@15136.4]
  assign RetimeWrapper_89_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15138.4]
  assign RetimeWrapper_89_io_in = _T_953 & io_rPort_7_en_0; // @[package.scala 94:16:@15137.4]
  assign RetimeWrapper_90_clock = clock; // @[:@15143.4]
  assign RetimeWrapper_90_reset = reset; // @[:@15144.4]
  assign RetimeWrapper_90_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15146.4]
  assign RetimeWrapper_90_io_in = _T_1045 & io_rPort_7_en_0; // @[package.scala 94:16:@15145.4]
  assign RetimeWrapper_91_clock = clock; // @[:@15151.4]
  assign RetimeWrapper_91_reset = reset; // @[:@15152.4]
  assign RetimeWrapper_91_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15154.4]
  assign RetimeWrapper_91_io_in = _T_1137 & io_rPort_7_en_0; // @[package.scala 94:16:@15153.4]
  assign RetimeWrapper_92_clock = clock; // @[:@15159.4]
  assign RetimeWrapper_92_reset = reset; // @[:@15160.4]
  assign RetimeWrapper_92_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15162.4]
  assign RetimeWrapper_92_io_in = _T_1229 & io_rPort_7_en_0; // @[package.scala 94:16:@15161.4]
  assign RetimeWrapper_93_clock = clock; // @[:@15167.4]
  assign RetimeWrapper_93_reset = reset; // @[:@15168.4]
  assign RetimeWrapper_93_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15170.4]
  assign RetimeWrapper_93_io_in = _T_1321 & io_rPort_7_en_0; // @[package.scala 94:16:@15169.4]
  assign RetimeWrapper_94_clock = clock; // @[:@15175.4]
  assign RetimeWrapper_94_reset = reset; // @[:@15176.4]
  assign RetimeWrapper_94_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15178.4]
  assign RetimeWrapper_94_io_in = _T_1413 & io_rPort_7_en_0; // @[package.scala 94:16:@15177.4]
  assign RetimeWrapper_95_clock = clock; // @[:@15183.4]
  assign RetimeWrapper_95_reset = reset; // @[:@15184.4]
  assign RetimeWrapper_95_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@15186.4]
  assign RetimeWrapper_95_io_in = _T_1505 & io_rPort_7_en_0; // @[package.scala 94:16:@15185.4]
  assign RetimeWrapper_96_clock = clock; // @[:@15239.4]
  assign RetimeWrapper_96_reset = reset; // @[:@15240.4]
  assign RetimeWrapper_96_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15242.4]
  assign RetimeWrapper_96_io_in = _T_499 & io_rPort_8_en_0; // @[package.scala 94:16:@15241.4]
  assign RetimeWrapper_97_clock = clock; // @[:@15247.4]
  assign RetimeWrapper_97_reset = reset; // @[:@15248.4]
  assign RetimeWrapper_97_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15250.4]
  assign RetimeWrapper_97_io_in = _T_591 & io_rPort_8_en_0; // @[package.scala 94:16:@15249.4]
  assign RetimeWrapper_98_clock = clock; // @[:@15255.4]
  assign RetimeWrapper_98_reset = reset; // @[:@15256.4]
  assign RetimeWrapper_98_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15258.4]
  assign RetimeWrapper_98_io_in = _T_683 & io_rPort_8_en_0; // @[package.scala 94:16:@15257.4]
  assign RetimeWrapper_99_clock = clock; // @[:@15263.4]
  assign RetimeWrapper_99_reset = reset; // @[:@15264.4]
  assign RetimeWrapper_99_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15266.4]
  assign RetimeWrapper_99_io_in = _T_775 & io_rPort_8_en_0; // @[package.scala 94:16:@15265.4]
  assign RetimeWrapper_100_clock = clock; // @[:@15271.4]
  assign RetimeWrapper_100_reset = reset; // @[:@15272.4]
  assign RetimeWrapper_100_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15274.4]
  assign RetimeWrapper_100_io_in = _T_867 & io_rPort_8_en_0; // @[package.scala 94:16:@15273.4]
  assign RetimeWrapper_101_clock = clock; // @[:@15279.4]
  assign RetimeWrapper_101_reset = reset; // @[:@15280.4]
  assign RetimeWrapper_101_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15282.4]
  assign RetimeWrapper_101_io_in = _T_959 & io_rPort_8_en_0; // @[package.scala 94:16:@15281.4]
  assign RetimeWrapper_102_clock = clock; // @[:@15287.4]
  assign RetimeWrapper_102_reset = reset; // @[:@15288.4]
  assign RetimeWrapper_102_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15290.4]
  assign RetimeWrapper_102_io_in = _T_1051 & io_rPort_8_en_0; // @[package.scala 94:16:@15289.4]
  assign RetimeWrapper_103_clock = clock; // @[:@15295.4]
  assign RetimeWrapper_103_reset = reset; // @[:@15296.4]
  assign RetimeWrapper_103_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15298.4]
  assign RetimeWrapper_103_io_in = _T_1143 & io_rPort_8_en_0; // @[package.scala 94:16:@15297.4]
  assign RetimeWrapper_104_clock = clock; // @[:@15303.4]
  assign RetimeWrapper_104_reset = reset; // @[:@15304.4]
  assign RetimeWrapper_104_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15306.4]
  assign RetimeWrapper_104_io_in = _T_1235 & io_rPort_8_en_0; // @[package.scala 94:16:@15305.4]
  assign RetimeWrapper_105_clock = clock; // @[:@15311.4]
  assign RetimeWrapper_105_reset = reset; // @[:@15312.4]
  assign RetimeWrapper_105_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15314.4]
  assign RetimeWrapper_105_io_in = _T_1327 & io_rPort_8_en_0; // @[package.scala 94:16:@15313.4]
  assign RetimeWrapper_106_clock = clock; // @[:@15319.4]
  assign RetimeWrapper_106_reset = reset; // @[:@15320.4]
  assign RetimeWrapper_106_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15322.4]
  assign RetimeWrapper_106_io_in = _T_1419 & io_rPort_8_en_0; // @[package.scala 94:16:@15321.4]
  assign RetimeWrapper_107_clock = clock; // @[:@15327.4]
  assign RetimeWrapper_107_reset = reset; // @[:@15328.4]
  assign RetimeWrapper_107_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15330.4]
  assign RetimeWrapper_107_io_in = _T_1511 & io_rPort_8_en_0; // @[package.scala 94:16:@15329.4]
endmodule
module RetimeWrapper_171( // @[:@15358.2]
  input         clock, // @[:@15359.4]
  input         reset, // @[:@15360.4]
  input         io_flow, // @[:@15361.4]
  input  [31:0] io_in, // @[:@15361.4]
  output [31:0] io_out // @[:@15361.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15363.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15363.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15363.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15363.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15363.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15363.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@15363.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15376.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15375.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15374.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15373.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15372.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15370.4]
endmodule
module RetimeWrapper_185( // @[:@17063.2]
  input         clock, // @[:@17064.4]
  input         reset, // @[:@17065.4]
  input         io_flow, // @[:@17066.4]
  input  [31:0] io_in, // @[:@17066.4]
  output [31:0] io_out // @[:@17066.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17068.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17068.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17068.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17068.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17068.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17068.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@17068.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17081.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17080.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17079.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17078.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17077.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17075.4]
endmodule
module x323_div( // @[:@17124.2]
  input         clock, // @[:@17125.4]
  input         reset, // @[:@17126.4]
  input  [31:0] io_a, // @[:@17127.4]
  input         io_flow, // @[:@17127.4]
  output [31:0] io_result // @[:@17127.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@17136.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@17136.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@17136.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@17136.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@17136.4]
  wire [31:0] __io_b; // @[Math.scala 709:24:@17149.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@17149.4]
  wire [31:0] _T_15; // @[FixedPoint.scala 24:59:@17133.4]
  wire [32:0] _T_17; // @[BigIPSim.scala 23:39:@17135.4]
  wire [32:0] _T_18; // @[package.scala 94:23:@17139.4]
  wire [31:0] _T_21; // @[package.scala 96:25:@17143.4]
  RetimeWrapper_185 RetimeWrapper ( // @[package.scala 93:22:@17136.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  _ _ ( // @[Math.scala 709:24:@17149.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  assign _T_15 = $signed(io_a); // @[FixedPoint.scala 24:59:@17133.4]
  assign _T_17 = $signed(_T_15) / $signed(32'sh3); // @[BigIPSim.scala 23:39:@17135.4]
  assign _T_18 = $unsigned(_T_17); // @[package.scala 94:23:@17139.4]
  assign _T_21 = $signed(RetimeWrapper_io_out); // @[package.scala 96:25:@17143.4]
  assign io_result = __io_result; // @[Math.scala 290:34:@17157.4]
  assign RetimeWrapper_clock = clock; // @[:@17137.4]
  assign RetimeWrapper_reset = reset; // @[:@17138.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@17141.4]
  assign RetimeWrapper_io_in = _T_18[31:0]; // @[package.scala 94:16:@17140.4]
  assign __io_b = $unsigned(_T_21); // @[Math.scala 710:17:@17152.4]
endmodule
module RetimeWrapper_186( // @[:@17171.2]
  input         clock, // @[:@17172.4]
  input         reset, // @[:@17173.4]
  input         io_flow, // @[:@17174.4]
  input  [31:0] io_in, // @[:@17174.4]
  output [31:0] io_out // @[:@17174.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17176.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17176.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17176.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17176.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17176.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17176.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(17)) sr ( // @[RetimeShiftRegister.scala 15:20:@17176.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17189.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17188.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17187.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17186.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17185.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17183.4]
endmodule
module RetimeWrapper_188( // @[:@17392.2]
  input   clock, // @[:@17393.4]
  input   reset, // @[:@17394.4]
  input   io_flow, // @[:@17395.4]
  input   io_in, // @[:@17395.4]
  output  io_out // @[:@17395.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@17397.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@17397.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@17397.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17397.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17397.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17397.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@17397.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17410.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17409.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@17408.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17407.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17406.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17404.4]
endmodule
module RetimeWrapper_190( // @[:@17456.2]
  input         clock, // @[:@17457.4]
  input         reset, // @[:@17458.4]
  input         io_flow, // @[:@17459.4]
  input  [31:0] io_in, // @[:@17459.4]
  output [31:0] io_out // @[:@17459.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17461.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17461.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17461.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17461.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17461.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17461.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(13)) sr ( // @[RetimeShiftRegister.scala 15:20:@17461.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17474.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17473.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17472.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17471.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17470.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17468.4]
endmodule
module RetimeWrapper_191( // @[:@17488.2]
  input         clock, // @[:@17489.4]
  input         reset, // @[:@17490.4]
  input         io_flow, // @[:@17491.4]
  input  [31:0] io_in, // @[:@17491.4]
  output [31:0] io_out // @[:@17491.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17493.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17493.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17493.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17493.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17493.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17493.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(19)) sr ( // @[RetimeShiftRegister.scala 15:20:@17493.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17506.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17505.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17504.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17503.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17502.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17500.4]
endmodule
module RetimeWrapper_192( // @[:@17520.2]
  input        clock, // @[:@17521.4]
  input        reset, // @[:@17522.4]
  input        io_flow, // @[:@17523.4]
  input  [7:0] io_in, // @[:@17523.4]
  output [7:0] io_out // @[:@17523.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17525.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17525.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17525.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17525.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17525.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17525.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@17525.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17538.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17537.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@17536.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17535.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17534.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17532.4]
endmodule
module RetimeWrapper_194( // @[:@17584.2]
  input         clock, // @[:@17585.4]
  input         reset, // @[:@17586.4]
  input         io_flow, // @[:@17587.4]
  input  [31:0] io_in, // @[:@17587.4]
  output [31:0] io_out // @[:@17587.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17589.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17589.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17589.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17589.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17589.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17589.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(23)) sr ( // @[RetimeShiftRegister.scala 15:20:@17589.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17602.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17601.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17600.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17599.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17598.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17596.4]
endmodule
module RetimeWrapper_200( // @[:@17933.2]
  input         clock, // @[:@17934.4]
  input         reset, // @[:@17935.4]
  input         io_flow, // @[:@17936.4]
  input  [31:0] io_in, // @[:@17936.4]
  output [31:0] io_out // @[:@17936.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@17938.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@17938.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@17938.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@17938.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@17938.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@17938.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(18)) sr ( // @[RetimeShiftRegister.scala 15:20:@17938.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@17951.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@17950.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@17949.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@17948.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@17947.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@17945.4]
endmodule
module RetimeWrapper_203( // @[:@18186.2]
  input   clock, // @[:@18187.4]
  input   reset, // @[:@18188.4]
  input   io_flow, // @[:@18189.4]
  input   io_in, // @[:@18189.4]
  output  io_out // @[:@18189.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@18191.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@18191.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@18191.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18191.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18191.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18191.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(45)) sr ( // @[RetimeShiftRegister.scala 15:20:@18191.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18204.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18203.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@18202.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18201.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18200.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18198.4]
endmodule
module RetimeWrapper_205( // @[:@18250.2]
  input         clock, // @[:@18251.4]
  input         reset, // @[:@18252.4]
  input         io_flow, // @[:@18253.4]
  input  [31:0] io_in, // @[:@18253.4]
  output [31:0] io_out // @[:@18253.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@18255.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@18255.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@18255.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18255.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18255.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18255.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(37)) sr ( // @[RetimeShiftRegister.scala 15:20:@18255.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18268.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18267.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@18266.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18265.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18264.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18262.4]
endmodule
module RetimeWrapper_206( // @[:@18282.2]
  input         clock, // @[:@18283.4]
  input         reset, // @[:@18284.4]
  input         io_flow, // @[:@18285.4]
  input  [31:0] io_in, // @[:@18285.4]
  output [31:0] io_out // @[:@18285.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@18287.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@18287.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@18287.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@18287.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@18287.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@18287.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@18287.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@18300.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@18299.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@18298.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@18297.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@18296.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@18294.4]
endmodule
module RetimeWrapper_230( // @[:@20541.2]
  input         clock, // @[:@20542.4]
  input         reset, // @[:@20543.4]
  input         io_flow, // @[:@20544.4]
  input  [31:0] io_in, // @[:@20544.4]
  output [31:0] io_out // @[:@20544.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@20546.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@20546.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@20546.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@20546.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@20546.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@20546.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(12)) sr ( // @[RetimeShiftRegister.scala 15:20:@20546.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@20559.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@20558.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@20557.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@20556.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@20555.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@20553.4]
endmodule
module RetimeWrapper_231( // @[:@20573.2]
  input   clock, // @[:@20574.4]
  input   reset, // @[:@20575.4]
  input   io_flow, // @[:@20576.4]
  input   io_in, // @[:@20576.4]
  output  io_out // @[:@20576.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@20578.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@20578.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@20578.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@20578.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@20578.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@20578.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@20578.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@20591.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@20590.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@20589.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@20588.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@20587.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@20585.4]
endmodule
module RetimeWrapper_289( // @[:@25492.2]
  input        clock, // @[:@25493.4]
  input        reset, // @[:@25494.4]
  input        io_flow, // @[:@25495.4]
  input  [8:0] io_in, // @[:@25495.4]
  output [8:0] io_out // @[:@25495.4]
);
  wire [8:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@25497.4]
  wire [8:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@25497.4]
  wire [8:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@25497.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@25497.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@25497.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@25497.4]
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@25497.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@25510.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@25509.4]
  assign sr_init = 9'h0; // @[RetimeShiftRegister.scala 19:16:@25508.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@25507.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@25506.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@25504.4]
endmodule
module SimBlackBoxesfix2fixBox_94( // @[:@25672.2]
  input  [7:0] io_a, // @[:@25675.4]
  output [8:0] io_b // @[:@25675.4]
);
  assign io_b = {1'h0,io_a}; // @[SimBlackBoxes.scala 99:40:@25689.4]
endmodule
module __93( // @[:@25691.2]
  input  [7:0] io_b, // @[:@25694.4]
  output [8:0] io_result // @[:@25694.4]
);
  wire [7:0] SimBlackBoxesfix2fixBox_io_a; // @[BigIPSim.scala 239:30:@25699.4]
  wire [8:0] SimBlackBoxesfix2fixBox_io_b; // @[BigIPSim.scala 239:30:@25699.4]
  SimBlackBoxesfix2fixBox_94 SimBlackBoxesfix2fixBox ( // @[BigIPSim.scala 239:30:@25699.4]
    .io_a(SimBlackBoxesfix2fixBox_io_a),
    .io_b(SimBlackBoxesfix2fixBox_io_b)
  );
  assign io_result = SimBlackBoxesfix2fixBox_io_b; // @[Math.scala 706:17:@25712.4]
  assign SimBlackBoxesfix2fixBox_io_a = io_b; // @[BigIPSim.scala 241:23:@25707.4]
endmodule
module fix2fixBox_43( // @[:@25756.2]
  input  [8:0] io_a, // @[:@25759.4]
  output [7:0] io_b // @[:@25759.4]
);
  assign io_b = io_a[7:0]; // @[Converter.scala 95:38:@25772.4]
endmodule
module x403_x15( // @[:@25774.2]
  input  [7:0] io_a, // @[:@25777.4]
  input  [7:0] io_b, // @[:@25777.4]
  output [7:0] io_result // @[:@25777.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@25785.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@25785.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@25792.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@25792.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@25802.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@25802.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@25790.4 Math.scala 713:14:@25791.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@25797.4 Math.scala 713:14:@25798.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@25799.4]
  __93 _ ( // @[Math.scala 709:24:@25785.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __93 __1 ( // @[Math.scala 709:24:@25792.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_43 fix2fixBox ( // @[Math.scala 141:30:@25802.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@25790.4 Math.scala 713:14:@25791.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@25797.4 Math.scala 713:14:@25798.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@25799.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@25810.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@25788.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@25795.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@25805.4]
endmodule
module fix2fixBox_50( // @[:@26864.2]
  input        clock, // @[:@26865.4]
  input        reset, // @[:@26866.4]
  input  [8:0] io_a, // @[:@26867.4]
  input        io_flow, // @[:@26867.4]
  output [7:0] io_b // @[:@26867.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@26880.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@26880.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@26880.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@26880.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@26880.4]
  RetimeWrapper_50 RetimeWrapper ( // @[package.scala 93:22:@26880.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@26887.4]
  assign RetimeWrapper_clock = clock; // @[:@26881.4]
  assign RetimeWrapper_reset = reset; // @[:@26882.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@26884.4]
  assign RetimeWrapper_io_in = io_a[7:0]; // @[package.scala 94:16:@26883.4]
endmodule
module x410_sum( // @[:@26889.2]
  input        clock, // @[:@26890.4]
  input        reset, // @[:@26891.4]
  input  [7:0] io_a, // @[:@26892.4]
  input  [7:0] io_b, // @[:@26892.4]
  input        io_flow, // @[:@26892.4]
  output [7:0] io_result // @[:@26892.4]
);
  wire [7:0] __io_b; // @[Math.scala 709:24:@26900.4]
  wire [8:0] __io_result; // @[Math.scala 709:24:@26900.4]
  wire [7:0] __1_io_b; // @[Math.scala 709:24:@26907.4]
  wire [8:0] __1_io_result; // @[Math.scala 709:24:@26907.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@26917.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@26917.4]
  wire [8:0] fix2fixBox_io_a; // @[Math.scala 141:30:@26917.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@26917.4]
  wire [7:0] fix2fixBox_io_b; // @[Math.scala 141:30:@26917.4]
  wire [8:0] a_upcast_number; // @[Math.scala 712:22:@26905.4 Math.scala 713:14:@26906.4]
  wire [8:0] b_upcast_number; // @[Math.scala 712:22:@26912.4 Math.scala 713:14:@26913.4]
  wire [9:0] _T_21; // @[Math.scala 136:37:@26914.4]
  __93 _ ( // @[Math.scala 709:24:@26900.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __93 __1 ( // @[Math.scala 709:24:@26907.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_50 fix2fixBox ( // @[Math.scala 141:30:@26917.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 712:22:@26905.4 Math.scala 713:14:@26906.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 712:22:@26912.4 Math.scala 713:14:@26913.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@26914.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@26925.4]
  assign __io_b = io_a; // @[Math.scala 710:17:@26903.4]
  assign __1_io_b = io_b; // @[Math.scala 710:17:@26910.4]
  assign fix2fixBox_clock = clock; // @[:@26918.4]
  assign fix2fixBox_reset = reset; // @[:@26919.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@26920.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@26923.4]
endmodule
module RetimeWrapper_299( // @[:@26939.2]
  input        clock, // @[:@26940.4]
  input        reset, // @[:@26941.4]
  input        io_flow, // @[:@26942.4]
  input  [7:0] io_in, // @[:@26942.4]
  output [7:0] io_out // @[:@26942.4]
);
  wire [7:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@26944.4]
  wire [7:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@26944.4]
  wire [7:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@26944.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@26944.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@26944.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@26944.4]
  RetimeShiftRegister #(.WIDTH(8), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@26944.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@26957.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@26956.4]
  assign sr_init = 8'h0; // @[RetimeShiftRegister.scala 19:16:@26955.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@26954.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@26953.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@26951.4]
endmodule
module x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@27055.2]
  input          clock, // @[:@27056.4]
  input          reset, // @[:@27057.4]
  output         io_in_x279_TVALID, // @[:@27058.4]
  input          io_in_x279_TREADY, // @[:@27058.4]
  output [255:0] io_in_x279_TDATA, // @[:@27058.4]
  output         io_in_x278_TREADY, // @[:@27058.4]
  input  [255:0] io_in_x278_TDATA, // @[:@27058.4]
  input  [7:0]   io_in_x278_TID, // @[:@27058.4]
  input  [7:0]   io_in_x278_TDEST, // @[:@27058.4]
  input          io_sigsIn_backpressure, // @[:@27058.4]
  input          io_sigsIn_datapathEn, // @[:@27058.4]
  input          io_sigsIn_break, // @[:@27058.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@27058.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@27058.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@27058.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@27058.4]
  input          io_rr // @[:@27058.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@27072.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@27072.4]
  wire [31:0] __1_io_b; // @[Math.scala 709:24:@27084.4]
  wire [31:0] __1_io_result; // @[Math.scala 709:24:@27084.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@27107.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@27107.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@27107.4]
  wire [7:0] RetimeWrapper_io_in; // @[package.scala 93:22:@27107.4]
  wire [7:0] RetimeWrapper_io_out; // @[package.scala 93:22:@27107.4]
  wire  x311_lb_0_clock; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_reset; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [1:0] x311_lb_0_io_rPort_8_banks_1; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [2:0] x311_lb_0_io_rPort_8_banks_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [9:0] x311_lb_0_io_rPort_8_ofs_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_rPort_8_en_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_rPort_8_backpressure; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [7:0] x311_lb_0_io_rPort_8_output_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [1:0] x311_lb_0_io_rPort_7_banks_1; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [2:0] x311_lb_0_io_rPort_7_banks_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [9:0] x311_lb_0_io_rPort_7_ofs_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_rPort_7_en_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_rPort_7_backpressure; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [7:0] x311_lb_0_io_rPort_7_output_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [1:0] x311_lb_0_io_rPort_6_banks_1; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [2:0] x311_lb_0_io_rPort_6_banks_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [9:0] x311_lb_0_io_rPort_6_ofs_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_rPort_6_en_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_rPort_6_backpressure; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [7:0] x311_lb_0_io_rPort_6_output_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [1:0] x311_lb_0_io_rPort_5_banks_1; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [2:0] x311_lb_0_io_rPort_5_banks_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [9:0] x311_lb_0_io_rPort_5_ofs_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_rPort_5_en_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_rPort_5_backpressure; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [7:0] x311_lb_0_io_rPort_5_output_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [1:0] x311_lb_0_io_rPort_4_banks_1; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [2:0] x311_lb_0_io_rPort_4_banks_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [9:0] x311_lb_0_io_rPort_4_ofs_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_rPort_4_en_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_rPort_4_backpressure; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [7:0] x311_lb_0_io_rPort_4_output_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [1:0] x311_lb_0_io_rPort_3_banks_1; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [2:0] x311_lb_0_io_rPort_3_banks_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [9:0] x311_lb_0_io_rPort_3_ofs_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_rPort_3_en_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_rPort_3_backpressure; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [7:0] x311_lb_0_io_rPort_3_output_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [1:0] x311_lb_0_io_rPort_2_banks_1; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [2:0] x311_lb_0_io_rPort_2_banks_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [9:0] x311_lb_0_io_rPort_2_ofs_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_rPort_2_en_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_rPort_2_backpressure; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [7:0] x311_lb_0_io_rPort_2_output_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [1:0] x311_lb_0_io_rPort_1_banks_1; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [2:0] x311_lb_0_io_rPort_1_banks_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [9:0] x311_lb_0_io_rPort_1_ofs_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_rPort_1_en_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_rPort_1_backpressure; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [7:0] x311_lb_0_io_rPort_1_output_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [1:0] x311_lb_0_io_rPort_0_banks_1; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [2:0] x311_lb_0_io_rPort_0_banks_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [9:0] x311_lb_0_io_rPort_0_ofs_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_rPort_0_en_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_rPort_0_backpressure; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [7:0] x311_lb_0_io_rPort_0_output_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [1:0] x311_lb_0_io_wPort_0_banks_1; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [2:0] x311_lb_0_io_wPort_0_banks_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [9:0] x311_lb_0_io_wPort_0_ofs_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire [7:0] x311_lb_0_io_wPort_0_data_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  x311_lb_0_io_wPort_0_en_0; // @[m_x311_lb_0.scala 35:17:@27117.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@27239.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@27239.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@27239.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@27239.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@27239.4]
  wire  x474_sum_1_clock; // @[Math.scala 150:24:@27279.4]
  wire  x474_sum_1_reset; // @[Math.scala 150:24:@27279.4]
  wire [31:0] x474_sum_1_io_a; // @[Math.scala 150:24:@27279.4]
  wire [31:0] x474_sum_1_io_b; // @[Math.scala 150:24:@27279.4]
  wire  x474_sum_1_io_flow; // @[Math.scala 150:24:@27279.4]
  wire [31:0] x474_sum_1_io_result; // @[Math.scala 150:24:@27279.4]
  wire  x477_sum_1_clock; // @[Math.scala 150:24:@27309.4]
  wire  x477_sum_1_reset; // @[Math.scala 150:24:@27309.4]
  wire [31:0] x477_sum_1_io_a; // @[Math.scala 150:24:@27309.4]
  wire [31:0] x477_sum_1_io_b; // @[Math.scala 150:24:@27309.4]
  wire  x477_sum_1_io_flow; // @[Math.scala 150:24:@27309.4]
  wire [31:0] x477_sum_1_io_result; // @[Math.scala 150:24:@27309.4]
  wire  x480_sum_1_clock; // @[Math.scala 150:24:@27339.4]
  wire  x480_sum_1_reset; // @[Math.scala 150:24:@27339.4]
  wire [31:0] x480_sum_1_io_a; // @[Math.scala 150:24:@27339.4]
  wire [31:0] x480_sum_1_io_b; // @[Math.scala 150:24:@27339.4]
  wire  x480_sum_1_io_flow; // @[Math.scala 150:24:@27339.4]
  wire [31:0] x480_sum_1_io_result; // @[Math.scala 150:24:@27339.4]
  wire  x483_sum_1_clock; // @[Math.scala 150:24:@27369.4]
  wire  x483_sum_1_reset; // @[Math.scala 150:24:@27369.4]
  wire [31:0] x483_sum_1_io_a; // @[Math.scala 150:24:@27369.4]
  wire [31:0] x483_sum_1_io_b; // @[Math.scala 150:24:@27369.4]
  wire  x483_sum_1_io_flow; // @[Math.scala 150:24:@27369.4]
  wire [31:0] x483_sum_1_io_result; // @[Math.scala 150:24:@27369.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@27385.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@27385.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@27385.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@27385.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@27385.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@27402.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@27402.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@27402.4]
  wire [31:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@27402.4]
  wire [31:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@27402.4]
  wire  x486_sum_1_clock; // @[Math.scala 150:24:@27415.4]
  wire  x486_sum_1_reset; // @[Math.scala 150:24:@27415.4]
  wire [31:0] x486_sum_1_io_a; // @[Math.scala 150:24:@27415.4]
  wire [31:0] x486_sum_1_io_b; // @[Math.scala 150:24:@27415.4]
  wire  x486_sum_1_io_flow; // @[Math.scala 150:24:@27415.4]
  wire [31:0] x486_sum_1_io_result; // @[Math.scala 150:24:@27415.4]
  wire  x489_sum_1_clock; // @[Math.scala 150:24:@27445.4]
  wire  x489_sum_1_reset; // @[Math.scala 150:24:@27445.4]
  wire [31:0] x489_sum_1_io_a; // @[Math.scala 150:24:@27445.4]
  wire [31:0] x489_sum_1_io_b; // @[Math.scala 150:24:@27445.4]
  wire  x489_sum_1_io_flow; // @[Math.scala 150:24:@27445.4]
  wire [31:0] x489_sum_1_io_result; // @[Math.scala 150:24:@27445.4]
  wire  x492_sub_1_clock; // @[Math.scala 191:24:@27471.4]
  wire  x492_sub_1_reset; // @[Math.scala 191:24:@27471.4]
  wire [31:0] x492_sub_1_io_a; // @[Math.scala 191:24:@27471.4]
  wire [31:0] x492_sub_1_io_b; // @[Math.scala 191:24:@27471.4]
  wire  x492_sub_1_io_flow; // @[Math.scala 191:24:@27471.4]
  wire [31:0] x492_sub_1_io_result; // @[Math.scala 191:24:@27471.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@27481.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@27481.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@27481.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@27481.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@27481.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@27490.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@27490.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@27490.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@27490.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@27490.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@27499.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@27499.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@27499.4]
  wire [31:0] RetimeWrapper_6_io_in; // @[package.scala 93:22:@27499.4]
  wire [31:0] RetimeWrapper_6_io_out; // @[package.scala 93:22:@27499.4]
  wire  x496_sum_1_clock; // @[Math.scala 150:24:@27530.4]
  wire  x496_sum_1_reset; // @[Math.scala 150:24:@27530.4]
  wire [31:0] x496_sum_1_io_a; // @[Math.scala 150:24:@27530.4]
  wire [31:0] x496_sum_1_io_b; // @[Math.scala 150:24:@27530.4]
  wire  x496_sum_1_io_flow; // @[Math.scala 150:24:@27530.4]
  wire [31:0] x496_sum_1_io_result; // @[Math.scala 150:24:@27530.4]
  wire  x323_div_1_clock; // @[Math.scala 327:24:@27542.4]
  wire  x323_div_1_reset; // @[Math.scala 327:24:@27542.4]
  wire [31:0] x323_div_1_io_a; // @[Math.scala 327:24:@27542.4]
  wire  x323_div_1_io_flow; // @[Math.scala 327:24:@27542.4]
  wire [31:0] x323_div_1_io_result; // @[Math.scala 327:24:@27542.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@27552.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@27552.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@27552.4]
  wire [31:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@27552.4]
  wire [31:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@27552.4]
  wire  x324_sum_1_clock; // @[Math.scala 150:24:@27561.4]
  wire  x324_sum_1_reset; // @[Math.scala 150:24:@27561.4]
  wire [31:0] x324_sum_1_io_a; // @[Math.scala 150:24:@27561.4]
  wire [31:0] x324_sum_1_io_b; // @[Math.scala 150:24:@27561.4]
  wire  x324_sum_1_io_flow; // @[Math.scala 150:24:@27561.4]
  wire [31:0] x324_sum_1_io_result; // @[Math.scala 150:24:@27561.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@27571.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@27571.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@27571.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@27571.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@27571.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@27580.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@27580.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@27580.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@27580.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@27580.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@27589.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@27589.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@27589.4]
  wire [31:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@27589.4]
  wire [31:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@27589.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@27598.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@27598.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@27598.4]
  wire [31:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@27598.4]
  wire [31:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@27598.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@27607.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@27607.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@27607.4]
  wire [7:0] RetimeWrapper_12_io_in; // @[package.scala 93:22:@27607.4]
  wire [7:0] RetimeWrapper_12_io_out; // @[package.scala 93:22:@27607.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@27618.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@27618.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@27618.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@27618.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@27618.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@27639.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@27639.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@27639.4]
  wire [31:0] RetimeWrapper_14_io_in; // @[package.scala 93:22:@27639.4]
  wire [31:0] RetimeWrapper_14_io_out; // @[package.scala 93:22:@27639.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@27657.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@27657.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@27657.4]
  wire [31:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@27657.4]
  wire [31:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@27657.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@27675.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@27675.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@27675.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@27675.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@27675.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@27684.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@27684.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@27684.4]
  wire [31:0] RetimeWrapper_17_io_in; // @[package.scala 93:22:@27684.4]
  wire [31:0] RetimeWrapper_17_io_out; // @[package.scala 93:22:@27684.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@27698.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@27698.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@27698.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@27698.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@27698.4]
  wire  x501_sum_1_clock; // @[Math.scala 150:24:@27743.4]
  wire  x501_sum_1_reset; // @[Math.scala 150:24:@27743.4]
  wire [31:0] x501_sum_1_io_a; // @[Math.scala 150:24:@27743.4]
  wire [31:0] x501_sum_1_io_b; // @[Math.scala 150:24:@27743.4]
  wire  x501_sum_1_io_flow; // @[Math.scala 150:24:@27743.4]
  wire [31:0] x501_sum_1_io_result; // @[Math.scala 150:24:@27743.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@27753.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@27753.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@27753.4]
  wire [31:0] RetimeWrapper_19_io_in; // @[package.scala 93:22:@27753.4]
  wire [31:0] RetimeWrapper_19_io_out; // @[package.scala 93:22:@27753.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@27762.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@27762.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@27762.4]
  wire [31:0] RetimeWrapper_20_io_in; // @[package.scala 93:22:@27762.4]
  wire [31:0] RetimeWrapper_20_io_out; // @[package.scala 93:22:@27762.4]
  wire  x335_sum_1_clock; // @[Math.scala 150:24:@27771.4]
  wire  x335_sum_1_reset; // @[Math.scala 150:24:@27771.4]
  wire [31:0] x335_sum_1_io_a; // @[Math.scala 150:24:@27771.4]
  wire [31:0] x335_sum_1_io_b; // @[Math.scala 150:24:@27771.4]
  wire  x335_sum_1_io_flow; // @[Math.scala 150:24:@27771.4]
  wire [31:0] x335_sum_1_io_result; // @[Math.scala 150:24:@27771.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@27781.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@27781.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@27781.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@27781.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@27781.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@27790.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@27790.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@27790.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@27790.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@27790.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@27799.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@27799.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@27799.4]
  wire [31:0] RetimeWrapper_23_io_in; // @[package.scala 93:22:@27799.4]
  wire [31:0] RetimeWrapper_23_io_out; // @[package.scala 93:22:@27799.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@27808.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@27808.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@27808.4]
  wire [31:0] RetimeWrapper_24_io_in; // @[package.scala 93:22:@27808.4]
  wire [31:0] RetimeWrapper_24_io_out; // @[package.scala 93:22:@27808.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@27817.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@27817.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@27817.4]
  wire [31:0] RetimeWrapper_25_io_in; // @[package.scala 93:22:@27817.4]
  wire [31:0] RetimeWrapper_25_io_out; // @[package.scala 93:22:@27817.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@27826.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@27826.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@27826.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@27826.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@27826.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@27838.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@27838.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@27838.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@27838.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@27838.4]
  wire  x338_rdcol_1_clock; // @[Math.scala 191:24:@27861.4]
  wire  x338_rdcol_1_reset; // @[Math.scala 191:24:@27861.4]
  wire [31:0] x338_rdcol_1_io_a; // @[Math.scala 191:24:@27861.4]
  wire [31:0] x338_rdcol_1_io_b; // @[Math.scala 191:24:@27861.4]
  wire  x338_rdcol_1_io_flow; // @[Math.scala 191:24:@27861.4]
  wire [31:0] x338_rdcol_1_io_result; // @[Math.scala 191:24:@27861.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@27876.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@27876.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@27876.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@27876.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@27876.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@27885.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@27885.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@27885.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@27885.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@27885.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@27906.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@27906.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@27906.4]
  wire [31:0] RetimeWrapper_30_io_in; // @[package.scala 93:22:@27906.4]
  wire [31:0] RetimeWrapper_30_io_out; // @[package.scala 93:22:@27906.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@27923.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@27923.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@27923.4]
  wire [31:0] RetimeWrapper_31_io_in; // @[package.scala 93:22:@27923.4]
  wire [31:0] RetimeWrapper_31_io_out; // @[package.scala 93:22:@27923.4]
  wire  x504_sum_1_clock; // @[Math.scala 150:24:@27936.4]
  wire  x504_sum_1_reset; // @[Math.scala 150:24:@27936.4]
  wire [31:0] x504_sum_1_io_a; // @[Math.scala 150:24:@27936.4]
  wire [31:0] x504_sum_1_io_b; // @[Math.scala 150:24:@27936.4]
  wire  x504_sum_1_io_flow; // @[Math.scala 150:24:@27936.4]
  wire [31:0] x504_sum_1_io_result; // @[Math.scala 150:24:@27936.4]
  wire  x507_sum_1_clock; // @[Math.scala 150:24:@27966.4]
  wire  x507_sum_1_reset; // @[Math.scala 150:24:@27966.4]
  wire [31:0] x507_sum_1_io_a; // @[Math.scala 150:24:@27966.4]
  wire [31:0] x507_sum_1_io_b; // @[Math.scala 150:24:@27966.4]
  wire  x507_sum_1_io_flow; // @[Math.scala 150:24:@27966.4]
  wire [31:0] x507_sum_1_io_result; // @[Math.scala 150:24:@27966.4]
  wire  x510_sum_1_clock; // @[Math.scala 150:24:@27996.4]
  wire  x510_sum_1_reset; // @[Math.scala 150:24:@27996.4]
  wire [31:0] x510_sum_1_io_a; // @[Math.scala 150:24:@27996.4]
  wire [31:0] x510_sum_1_io_b; // @[Math.scala 150:24:@27996.4]
  wire  x510_sum_1_io_flow; // @[Math.scala 150:24:@27996.4]
  wire [31:0] x510_sum_1_io_result; // @[Math.scala 150:24:@27996.4]
  wire  x513_sum_1_clock; // @[Math.scala 150:24:@28026.4]
  wire  x513_sum_1_reset; // @[Math.scala 150:24:@28026.4]
  wire [31:0] x513_sum_1_io_a; // @[Math.scala 150:24:@28026.4]
  wire [31:0] x513_sum_1_io_b; // @[Math.scala 150:24:@28026.4]
  wire  x513_sum_1_io_flow; // @[Math.scala 150:24:@28026.4]
  wire [31:0] x513_sum_1_io_result; // @[Math.scala 150:24:@28026.4]
  wire  x516_sum_1_clock; // @[Math.scala 150:24:@28056.4]
  wire  x516_sum_1_reset; // @[Math.scala 150:24:@28056.4]
  wire [31:0] x516_sum_1_io_a; // @[Math.scala 150:24:@28056.4]
  wire [31:0] x516_sum_1_io_b; // @[Math.scala 150:24:@28056.4]
  wire  x516_sum_1_io_flow; // @[Math.scala 150:24:@28056.4]
  wire [31:0] x516_sum_1_io_result; // @[Math.scala 150:24:@28056.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@28072.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@28072.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@28072.4]
  wire [31:0] RetimeWrapper_32_io_in; // @[package.scala 93:22:@28072.4]
  wire [31:0] RetimeWrapper_32_io_out; // @[package.scala 93:22:@28072.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@28089.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@28089.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@28089.4]
  wire [31:0] RetimeWrapper_33_io_in; // @[package.scala 93:22:@28089.4]
  wire [31:0] RetimeWrapper_33_io_out; // @[package.scala 93:22:@28089.4]
  wire  x519_sum_1_clock; // @[Math.scala 150:24:@28102.4]
  wire  x519_sum_1_reset; // @[Math.scala 150:24:@28102.4]
  wire [31:0] x519_sum_1_io_a; // @[Math.scala 150:24:@28102.4]
  wire [31:0] x519_sum_1_io_b; // @[Math.scala 150:24:@28102.4]
  wire  x519_sum_1_io_flow; // @[Math.scala 150:24:@28102.4]
  wire [31:0] x519_sum_1_io_result; // @[Math.scala 150:24:@28102.4]
  wire  x522_sub_1_clock; // @[Math.scala 191:24:@28130.4]
  wire  x522_sub_1_reset; // @[Math.scala 191:24:@28130.4]
  wire [31:0] x522_sub_1_io_a; // @[Math.scala 191:24:@28130.4]
  wire [31:0] x522_sub_1_io_b; // @[Math.scala 191:24:@28130.4]
  wire  x522_sub_1_io_flow; // @[Math.scala 191:24:@28130.4]
  wire [31:0] x522_sub_1_io_result; // @[Math.scala 191:24:@28130.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@28140.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@28140.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@28140.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@28140.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@28140.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@28149.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@28149.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@28149.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@28149.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@28149.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@28158.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@28158.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@28158.4]
  wire [31:0] RetimeWrapper_36_io_in; // @[package.scala 93:22:@28158.4]
  wire [31:0] RetimeWrapper_36_io_out; // @[package.scala 93:22:@28158.4]
  wire  x343_div_1_clock; // @[Math.scala 327:24:@28172.4]
  wire  x343_div_1_reset; // @[Math.scala 327:24:@28172.4]
  wire [31:0] x343_div_1_io_a; // @[Math.scala 327:24:@28172.4]
  wire  x343_div_1_io_flow; // @[Math.scala 327:24:@28172.4]
  wire [31:0] x343_div_1_io_result; // @[Math.scala 327:24:@28172.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@28182.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@28182.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@28182.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@28182.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@28182.4]
  wire  x344_sum_1_clock; // @[Math.scala 150:24:@28191.4]
  wire  x344_sum_1_reset; // @[Math.scala 150:24:@28191.4]
  wire [31:0] x344_sum_1_io_a; // @[Math.scala 150:24:@28191.4]
  wire [31:0] x344_sum_1_io_b; // @[Math.scala 150:24:@28191.4]
  wire  x344_sum_1_io_flow; // @[Math.scala 150:24:@28191.4]
  wire [31:0] x344_sum_1_io_result; // @[Math.scala 150:24:@28191.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@28201.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@28201.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@28201.4]
  wire [31:0] RetimeWrapper_38_io_in; // @[package.scala 93:22:@28201.4]
  wire [31:0] RetimeWrapper_38_io_out; // @[package.scala 93:22:@28201.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@28210.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@28210.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@28210.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@28210.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@28210.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@28222.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@28222.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@28222.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@28222.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@28222.4]
  wire  x347_rdcol_1_clock; // @[Math.scala 191:24:@28245.4]
  wire  x347_rdcol_1_reset; // @[Math.scala 191:24:@28245.4]
  wire [31:0] x347_rdcol_1_io_a; // @[Math.scala 191:24:@28245.4]
  wire [31:0] x347_rdcol_1_io_b; // @[Math.scala 191:24:@28245.4]
  wire  x347_rdcol_1_io_flow; // @[Math.scala 191:24:@28245.4]
  wire [31:0] x347_rdcol_1_io_result; // @[Math.scala 191:24:@28245.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@28260.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@28260.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@28260.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@28260.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@28260.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@28281.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@28281.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@28281.4]
  wire [31:0] RetimeWrapper_42_io_in; // @[package.scala 93:22:@28281.4]
  wire [31:0] RetimeWrapper_42_io_out; // @[package.scala 93:22:@28281.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@28298.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@28298.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@28298.4]
  wire [31:0] RetimeWrapper_43_io_in; // @[package.scala 93:22:@28298.4]
  wire [31:0] RetimeWrapper_43_io_out; // @[package.scala 93:22:@28298.4]
  wire  x526_sum_1_clock; // @[Math.scala 150:24:@28311.4]
  wire  x526_sum_1_reset; // @[Math.scala 150:24:@28311.4]
  wire [31:0] x526_sum_1_io_a; // @[Math.scala 150:24:@28311.4]
  wire [31:0] x526_sum_1_io_b; // @[Math.scala 150:24:@28311.4]
  wire  x526_sum_1_io_flow; // @[Math.scala 150:24:@28311.4]
  wire [31:0] x526_sum_1_io_result; // @[Math.scala 150:24:@28311.4]
  wire  x529_sum_1_clock; // @[Math.scala 150:24:@28341.4]
  wire  x529_sum_1_reset; // @[Math.scala 150:24:@28341.4]
  wire [31:0] x529_sum_1_io_a; // @[Math.scala 150:24:@28341.4]
  wire [31:0] x529_sum_1_io_b; // @[Math.scala 150:24:@28341.4]
  wire  x529_sum_1_io_flow; // @[Math.scala 150:24:@28341.4]
  wire [31:0] x529_sum_1_io_result; // @[Math.scala 150:24:@28341.4]
  wire  x532_sum_1_clock; // @[Math.scala 150:24:@28371.4]
  wire  x532_sum_1_reset; // @[Math.scala 150:24:@28371.4]
  wire [31:0] x532_sum_1_io_a; // @[Math.scala 150:24:@28371.4]
  wire [31:0] x532_sum_1_io_b; // @[Math.scala 150:24:@28371.4]
  wire  x532_sum_1_io_flow; // @[Math.scala 150:24:@28371.4]
  wire [31:0] x532_sum_1_io_result; // @[Math.scala 150:24:@28371.4]
  wire  x535_sum_1_clock; // @[Math.scala 150:24:@28401.4]
  wire  x535_sum_1_reset; // @[Math.scala 150:24:@28401.4]
  wire [31:0] x535_sum_1_io_a; // @[Math.scala 150:24:@28401.4]
  wire [31:0] x535_sum_1_io_b; // @[Math.scala 150:24:@28401.4]
  wire  x535_sum_1_io_flow; // @[Math.scala 150:24:@28401.4]
  wire [31:0] x535_sum_1_io_result; // @[Math.scala 150:24:@28401.4]
  wire  x538_sum_1_clock; // @[Math.scala 150:24:@28431.4]
  wire  x538_sum_1_reset; // @[Math.scala 150:24:@28431.4]
  wire [31:0] x538_sum_1_io_a; // @[Math.scala 150:24:@28431.4]
  wire [31:0] x538_sum_1_io_b; // @[Math.scala 150:24:@28431.4]
  wire  x538_sum_1_io_flow; // @[Math.scala 150:24:@28431.4]
  wire [31:0] x538_sum_1_io_result; // @[Math.scala 150:24:@28431.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@28447.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@28447.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@28447.4]
  wire [31:0] RetimeWrapper_44_io_in; // @[package.scala 93:22:@28447.4]
  wire [31:0] RetimeWrapper_44_io_out; // @[package.scala 93:22:@28447.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@28464.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@28464.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@28464.4]
  wire [31:0] RetimeWrapper_45_io_in; // @[package.scala 93:22:@28464.4]
  wire [31:0] RetimeWrapper_45_io_out; // @[package.scala 93:22:@28464.4]
  wire  x541_sum_1_clock; // @[Math.scala 150:24:@28477.4]
  wire  x541_sum_1_reset; // @[Math.scala 150:24:@28477.4]
  wire [31:0] x541_sum_1_io_a; // @[Math.scala 150:24:@28477.4]
  wire [31:0] x541_sum_1_io_b; // @[Math.scala 150:24:@28477.4]
  wire  x541_sum_1_io_flow; // @[Math.scala 150:24:@28477.4]
  wire [31:0] x541_sum_1_io_result; // @[Math.scala 150:24:@28477.4]
  wire  x544_sub_1_clock; // @[Math.scala 191:24:@28503.4]
  wire  x544_sub_1_reset; // @[Math.scala 191:24:@28503.4]
  wire [31:0] x544_sub_1_io_a; // @[Math.scala 191:24:@28503.4]
  wire [31:0] x544_sub_1_io_b; // @[Math.scala 191:24:@28503.4]
  wire  x544_sub_1_io_flow; // @[Math.scala 191:24:@28503.4]
  wire [31:0] x544_sub_1_io_result; // @[Math.scala 191:24:@28503.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@28513.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@28513.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@28513.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@28513.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@28513.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@28522.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@28522.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@28522.4]
  wire [31:0] RetimeWrapper_47_io_in; // @[package.scala 93:22:@28522.4]
  wire [31:0] RetimeWrapper_47_io_out; // @[package.scala 93:22:@28522.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@28531.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@28531.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@28531.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@28531.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@28531.4]
  wire  x352_div_1_clock; // @[Math.scala 327:24:@28545.4]
  wire  x352_div_1_reset; // @[Math.scala 327:24:@28545.4]
  wire [31:0] x352_div_1_io_a; // @[Math.scala 327:24:@28545.4]
  wire  x352_div_1_io_flow; // @[Math.scala 327:24:@28545.4]
  wire [31:0] x352_div_1_io_result; // @[Math.scala 327:24:@28545.4]
  wire  x353_sum_1_clock; // @[Math.scala 150:24:@28555.4]
  wire  x353_sum_1_reset; // @[Math.scala 150:24:@28555.4]
  wire [31:0] x353_sum_1_io_a; // @[Math.scala 150:24:@28555.4]
  wire [31:0] x353_sum_1_io_b; // @[Math.scala 150:24:@28555.4]
  wire  x353_sum_1_io_flow; // @[Math.scala 150:24:@28555.4]
  wire [31:0] x353_sum_1_io_result; // @[Math.scala 150:24:@28555.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@28565.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@28565.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@28565.4]
  wire [31:0] RetimeWrapper_49_io_in; // @[package.scala 93:22:@28565.4]
  wire [31:0] RetimeWrapper_49_io_out; // @[package.scala 93:22:@28565.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@28574.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@28574.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@28574.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@28574.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@28574.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@28586.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@28586.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@28586.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@28586.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@28586.4]
  wire  x356_rdrow_1_clock; // @[Math.scala 191:24:@28611.4]
  wire  x356_rdrow_1_reset; // @[Math.scala 191:24:@28611.4]
  wire [31:0] x356_rdrow_1_io_a; // @[Math.scala 191:24:@28611.4]
  wire [31:0] x356_rdrow_1_io_b; // @[Math.scala 191:24:@28611.4]
  wire  x356_rdrow_1_io_flow; // @[Math.scala 191:24:@28611.4]
  wire [31:0] x356_rdrow_1_io_result; // @[Math.scala 191:24:@28611.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@28628.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@28628.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@28628.4]
  wire [31:0] RetimeWrapper_52_io_in; // @[package.scala 93:22:@28628.4]
  wire [31:0] RetimeWrapper_52_io_out; // @[package.scala 93:22:@28628.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@28646.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@28646.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@28646.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@28646.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@28646.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@28655.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@28655.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@28655.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@28655.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@28655.4]
  wire  x550_sum_1_clock; // @[Math.scala 150:24:@28700.4]
  wire  x550_sum_1_reset; // @[Math.scala 150:24:@28700.4]
  wire [31:0] x550_sum_1_io_a; // @[Math.scala 150:24:@28700.4]
  wire [31:0] x550_sum_1_io_b; // @[Math.scala 150:24:@28700.4]
  wire  x550_sum_1_io_flow; // @[Math.scala 150:24:@28700.4]
  wire [31:0] x550_sum_1_io_result; // @[Math.scala 150:24:@28700.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@28710.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@28710.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@28710.4]
  wire [31:0] RetimeWrapper_55_io_in; // @[package.scala 93:22:@28710.4]
  wire [31:0] RetimeWrapper_55_io_out; // @[package.scala 93:22:@28710.4]
  wire  x364_sum_1_clock; // @[Math.scala 150:24:@28719.4]
  wire  x364_sum_1_reset; // @[Math.scala 150:24:@28719.4]
  wire [31:0] x364_sum_1_io_a; // @[Math.scala 150:24:@28719.4]
  wire [31:0] x364_sum_1_io_b; // @[Math.scala 150:24:@28719.4]
  wire  x364_sum_1_io_flow; // @[Math.scala 150:24:@28719.4]
  wire [31:0] x364_sum_1_io_result; // @[Math.scala 150:24:@28719.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@28729.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@28729.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@28729.4]
  wire [31:0] RetimeWrapper_56_io_in; // @[package.scala 93:22:@28729.4]
  wire [31:0] RetimeWrapper_56_io_out; // @[package.scala 93:22:@28729.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@28738.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@28738.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@28738.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@28738.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@28738.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@28747.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@28747.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@28747.4]
  wire [31:0] RetimeWrapper_58_io_in; // @[package.scala 93:22:@28747.4]
  wire [31:0] RetimeWrapper_58_io_out; // @[package.scala 93:22:@28747.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@28759.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@28759.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@28759.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@28759.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@28759.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@28786.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@28786.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@28786.4]
  wire [31:0] RetimeWrapper_60_io_in; // @[package.scala 93:22:@28786.4]
  wire [31:0] RetimeWrapper_60_io_out; // @[package.scala 93:22:@28786.4]
  wire  x369_sum_1_clock; // @[Math.scala 150:24:@28795.4]
  wire  x369_sum_1_reset; // @[Math.scala 150:24:@28795.4]
  wire [31:0] x369_sum_1_io_a; // @[Math.scala 150:24:@28795.4]
  wire [31:0] x369_sum_1_io_b; // @[Math.scala 150:24:@28795.4]
  wire  x369_sum_1_io_flow; // @[Math.scala 150:24:@28795.4]
  wire [31:0] x369_sum_1_io_result; // @[Math.scala 150:24:@28795.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@28805.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@28805.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@28805.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@28805.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@28805.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@28817.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@28817.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@28817.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@28817.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@28817.4]
  wire  x374_sum_1_clock; // @[Math.scala 150:24:@28844.4]
  wire  x374_sum_1_reset; // @[Math.scala 150:24:@28844.4]
  wire [31:0] x374_sum_1_io_a; // @[Math.scala 150:24:@28844.4]
  wire [31:0] x374_sum_1_io_b; // @[Math.scala 150:24:@28844.4]
  wire  x374_sum_1_io_flow; // @[Math.scala 150:24:@28844.4]
  wire [31:0] x374_sum_1_io_result; // @[Math.scala 150:24:@28844.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@28854.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@28854.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@28854.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@28854.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@28854.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@28866.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@28866.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@28866.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@28866.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@28866.4]
  wire  x377_rdrow_1_clock; // @[Math.scala 191:24:@28889.4]
  wire  x377_rdrow_1_reset; // @[Math.scala 191:24:@28889.4]
  wire [31:0] x377_rdrow_1_io_a; // @[Math.scala 191:24:@28889.4]
  wire [31:0] x377_rdrow_1_io_b; // @[Math.scala 191:24:@28889.4]
  wire  x377_rdrow_1_io_flow; // @[Math.scala 191:24:@28889.4]
  wire [31:0] x377_rdrow_1_io_result; // @[Math.scala 191:24:@28889.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@28906.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@28906.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@28906.4]
  wire [31:0] RetimeWrapper_65_io_in; // @[package.scala 93:22:@28906.4]
  wire [31:0] RetimeWrapper_65_io_out; // @[package.scala 93:22:@28906.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@28924.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@28924.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@28924.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@28924.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@28924.4]
  wire  x555_sum_1_clock; // @[Math.scala 150:24:@28969.4]
  wire  x555_sum_1_reset; // @[Math.scala 150:24:@28969.4]
  wire [31:0] x555_sum_1_io_a; // @[Math.scala 150:24:@28969.4]
  wire [31:0] x555_sum_1_io_b; // @[Math.scala 150:24:@28969.4]
  wire  x555_sum_1_io_flow; // @[Math.scala 150:24:@28969.4]
  wire [31:0] x555_sum_1_io_result; // @[Math.scala 150:24:@28969.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@28979.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@28979.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@28979.4]
  wire [31:0] RetimeWrapper_67_io_in; // @[package.scala 93:22:@28979.4]
  wire [31:0] RetimeWrapper_67_io_out; // @[package.scala 93:22:@28979.4]
  wire  x385_sum_1_clock; // @[Math.scala 150:24:@28988.4]
  wire  x385_sum_1_reset; // @[Math.scala 150:24:@28988.4]
  wire [31:0] x385_sum_1_io_a; // @[Math.scala 150:24:@28988.4]
  wire [31:0] x385_sum_1_io_b; // @[Math.scala 150:24:@28988.4]
  wire  x385_sum_1_io_flow; // @[Math.scala 150:24:@28988.4]
  wire [31:0] x385_sum_1_io_result; // @[Math.scala 150:24:@28988.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@28998.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@28998.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@28998.4]
  wire [31:0] RetimeWrapper_68_io_in; // @[package.scala 93:22:@28998.4]
  wire [31:0] RetimeWrapper_68_io_out; // @[package.scala 93:22:@28998.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@29007.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@29007.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@29007.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@29007.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@29007.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@29016.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@29016.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@29016.4]
  wire [31:0] RetimeWrapper_70_io_in; // @[package.scala 93:22:@29016.4]
  wire [31:0] RetimeWrapper_70_io_out; // @[package.scala 93:22:@29016.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@29028.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@29028.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@29028.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@29028.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@29028.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@29055.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@29055.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@29055.4]
  wire [31:0] RetimeWrapper_72_io_in; // @[package.scala 93:22:@29055.4]
  wire [31:0] RetimeWrapper_72_io_out; // @[package.scala 93:22:@29055.4]
  wire  x390_sum_1_clock; // @[Math.scala 150:24:@29066.4]
  wire  x390_sum_1_reset; // @[Math.scala 150:24:@29066.4]
  wire [31:0] x390_sum_1_io_a; // @[Math.scala 150:24:@29066.4]
  wire [31:0] x390_sum_1_io_b; // @[Math.scala 150:24:@29066.4]
  wire  x390_sum_1_io_flow; // @[Math.scala 150:24:@29066.4]
  wire [31:0] x390_sum_1_io_result; // @[Math.scala 150:24:@29066.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@29076.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@29076.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@29076.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@29076.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@29076.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@29088.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@29088.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@29088.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@29088.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@29088.4]
  wire  x395_sum_1_clock; // @[Math.scala 150:24:@29115.4]
  wire  x395_sum_1_reset; // @[Math.scala 150:24:@29115.4]
  wire [31:0] x395_sum_1_io_a; // @[Math.scala 150:24:@29115.4]
  wire [31:0] x395_sum_1_io_b; // @[Math.scala 150:24:@29115.4]
  wire  x395_sum_1_io_flow; // @[Math.scala 150:24:@29115.4]
  wire [31:0] x395_sum_1_io_result; // @[Math.scala 150:24:@29115.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@29125.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@29125.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@29125.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@29125.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@29125.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@29137.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@29137.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@29137.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@29137.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@29137.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@29160.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@29160.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@29160.4]
  wire [8:0] RetimeWrapper_77_io_in; // @[package.scala 93:22:@29160.4]
  wire [8:0] RetimeWrapper_77_io_out; // @[package.scala 93:22:@29160.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@29172.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@29172.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@29172.4]
  wire [8:0] RetimeWrapper_78_io_in; // @[package.scala 93:22:@29172.4]
  wire [8:0] RetimeWrapper_78_io_out; // @[package.scala 93:22:@29172.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@29184.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@29184.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@29184.4]
  wire [9:0] RetimeWrapper_79_io_in; // @[package.scala 93:22:@29184.4]
  wire [9:0] RetimeWrapper_79_io_out; // @[package.scala 93:22:@29184.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@29196.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@29196.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@29196.4]
  wire [8:0] RetimeWrapper_80_io_in; // @[package.scala 93:22:@29196.4]
  wire [8:0] RetimeWrapper_80_io_out; // @[package.scala 93:22:@29196.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@29208.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@29208.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@29208.4]
  wire [8:0] RetimeWrapper_81_io_in; // @[package.scala 93:22:@29208.4]
  wire [8:0] RetimeWrapper_81_io_out; // @[package.scala 93:22:@29208.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@29218.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@29218.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@29218.4]
  wire [7:0] RetimeWrapper_82_io_in; // @[package.scala 93:22:@29218.4]
  wire [7:0] RetimeWrapper_82_io_out; // @[package.scala 93:22:@29218.4]
  wire [7:0] x403_x15_1_io_a; // @[Math.scala 150:24:@29227.4]
  wire [7:0] x403_x15_1_io_b; // @[Math.scala 150:24:@29227.4]
  wire [7:0] x403_x15_1_io_result; // @[Math.scala 150:24:@29227.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@29237.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@29237.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@29237.4]
  wire [7:0] RetimeWrapper_83_io_in; // @[package.scala 93:22:@29237.4]
  wire [7:0] RetimeWrapper_83_io_out; // @[package.scala 93:22:@29237.4]
  wire [7:0] x404_x16_1_io_a; // @[Math.scala 150:24:@29246.4]
  wire [7:0] x404_x16_1_io_b; // @[Math.scala 150:24:@29246.4]
  wire [7:0] x404_x16_1_io_result; // @[Math.scala 150:24:@29246.4]
  wire [7:0] x405_x15_1_io_a; // @[Math.scala 150:24:@29256.4]
  wire [7:0] x405_x15_1_io_b; // @[Math.scala 150:24:@29256.4]
  wire [7:0] x405_x15_1_io_result; // @[Math.scala 150:24:@29256.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@29266.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@29266.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@29266.4]
  wire [7:0] RetimeWrapper_84_io_in; // @[package.scala 93:22:@29266.4]
  wire [7:0] RetimeWrapper_84_io_out; // @[package.scala 93:22:@29266.4]
  wire [7:0] x406_x16_1_io_a; // @[Math.scala 150:24:@29275.4]
  wire [7:0] x406_x16_1_io_b; // @[Math.scala 150:24:@29275.4]
  wire [7:0] x406_x16_1_io_result; // @[Math.scala 150:24:@29275.4]
  wire [7:0] x407_x15_1_io_a; // @[Math.scala 150:24:@29285.4]
  wire [7:0] x407_x15_1_io_b; // @[Math.scala 150:24:@29285.4]
  wire [7:0] x407_x15_1_io_result; // @[Math.scala 150:24:@29285.4]
  wire [7:0] x408_x16_1_io_a; // @[Math.scala 150:24:@29295.4]
  wire [7:0] x408_x16_1_io_b; // @[Math.scala 150:24:@29295.4]
  wire [7:0] x408_x16_1_io_result; // @[Math.scala 150:24:@29295.4]
  wire [7:0] x409_x15_1_io_a; // @[Math.scala 150:24:@29305.4]
  wire [7:0] x409_x15_1_io_b; // @[Math.scala 150:24:@29305.4]
  wire [7:0] x409_x15_1_io_result; // @[Math.scala 150:24:@29305.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@29315.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@29315.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@29315.4]
  wire [7:0] RetimeWrapper_85_io_in; // @[package.scala 93:22:@29315.4]
  wire [7:0] RetimeWrapper_85_io_out; // @[package.scala 93:22:@29315.4]
  wire  x410_sum_1_clock; // @[Math.scala 150:24:@29324.4]
  wire  x410_sum_1_reset; // @[Math.scala 150:24:@29324.4]
  wire [7:0] x410_sum_1_io_a; // @[Math.scala 150:24:@29324.4]
  wire [7:0] x410_sum_1_io_b; // @[Math.scala 150:24:@29324.4]
  wire  x410_sum_1_io_flow; // @[Math.scala 150:24:@29324.4]
  wire [7:0] x410_sum_1_io_result; // @[Math.scala 150:24:@29324.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@29345.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@29345.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@29345.4]
  wire [7:0] RetimeWrapper_86_io_in; // @[package.scala 93:22:@29345.4]
  wire [7:0] RetimeWrapper_86_io_out; // @[package.scala 93:22:@29345.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@29354.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@29354.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@29354.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@29354.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@29354.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@29363.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@29363.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@29363.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@29363.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@29363.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@29372.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@29372.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@29372.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@29372.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@29372.4]
  wire  b307; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 62:18:@27092.4]
  wire  b308; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 63:18:@27093.4]
  wire  _T_205; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 67:30:@27095.4]
  wire  _T_206; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 67:37:@27096.4]
  wire  _T_210; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 69:76:@27101.4]
  wire  _T_211; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 69:62:@27102.4]
  wire  _T_213; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 69:101:@27103.4]
  wire [31:0] b305_number; // @[Math.scala 712:22:@27077.4 Math.scala 713:14:@27078.4]
  wire [31:0] _T_240; // @[Math.scala 499:52:@27193.4]
  wire  x314; // @[Math.scala 499:44:@27201.4]
  wire  x315; // @[Math.scala 499:44:@27208.4]
  wire  x316; // @[Math.scala 499:44:@27215.4]
  wire [31:0] _T_287; // @[Mux.scala 19:72:@27227.4]
  wire [31:0] _T_289; // @[Mux.scala 19:72:@27228.4]
  wire [31:0] _T_291; // @[Mux.scala 19:72:@27229.4]
  wire [31:0] _T_293; // @[Mux.scala 19:72:@27231.4]
  wire [31:0] x562_x317_D2_number; // @[package.scala 96:25:@27244.4 package.scala 96:25:@27245.4]
  wire [31:0] _T_308; // @[Math.scala 406:49:@27251.4]
  wire [31:0] _T_310; // @[Math.scala 406:56:@27253.4]
  wire [31:0] _T_311; // @[Math.scala 406:56:@27254.4]
  wire [31:0] b306_number; // @[Math.scala 712:22:@27089.4 Math.scala 713:14:@27090.4]
  wire  _T_316; // @[FixedPoint.scala 50:25:@27260.4]
  wire [15:0] _T_320; // @[Bitwise.scala 72:12:@27262.4]
  wire [15:0] _T_321; // @[FixedPoint.scala 18:52:@27263.4]
  wire [31:0] _T_330; // @[Math.scala 406:49:@27271.4]
  wire [31:0] _T_332; // @[Math.scala 406:56:@27273.4]
  wire [31:0] _T_333; // @[Math.scala 406:56:@27274.4]
  wire [31:0] x474_sum_number; // @[Math.scala 154:22:@27285.4 Math.scala 155:14:@27286.4]
  wire  _T_341; // @[FixedPoint.scala 50:25:@27290.4]
  wire [7:0] _T_345; // @[Bitwise.scala 72:12:@27292.4]
  wire [23:0] _T_346; // @[FixedPoint.scala 18:52:@27293.4]
  wire [31:0] _T_355; // @[Math.scala 406:49:@27301.4]
  wire [31:0] _T_357; // @[Math.scala 406:56:@27303.4]
  wire [31:0] _T_358; // @[Math.scala 406:56:@27304.4]
  wire [31:0] x477_sum_number; // @[Math.scala 154:22:@27315.4 Math.scala 155:14:@27316.4]
  wire  _T_366; // @[FixedPoint.scala 50:25:@27320.4]
  wire [3:0] _T_370; // @[Bitwise.scala 72:12:@27322.4]
  wire [27:0] _T_371; // @[FixedPoint.scala 18:52:@27323.4]
  wire [31:0] _T_380; // @[Math.scala 406:49:@27331.4]
  wire [31:0] _T_382; // @[Math.scala 406:56:@27333.4]
  wire [31:0] _T_383; // @[Math.scala 406:56:@27334.4]
  wire [31:0] x480_sum_number; // @[Math.scala 154:22:@27345.4 Math.scala 155:14:@27346.4]
  wire  _T_391; // @[FixedPoint.scala 50:25:@27350.4]
  wire [1:0] _T_395; // @[Bitwise.scala 72:12:@27352.4]
  wire [29:0] _T_396; // @[FixedPoint.scala 18:52:@27353.4]
  wire [31:0] _T_405; // @[Math.scala 406:49:@27361.4]
  wire [31:0] _T_407; // @[Math.scala 406:56:@27363.4]
  wire [31:0] _T_408; // @[Math.scala 406:56:@27364.4]
  wire [31:0] x483_sum_number; // @[Math.scala 154:22:@27375.4 Math.scala 155:14:@27376.4]
  wire  _T_416; // @[FixedPoint.scala 50:25:@27380.4]
  wire [1:0] _T_420; // @[Bitwise.scala 72:12:@27382.4]
  wire [29:0] _T_421; // @[FixedPoint.scala 18:52:@27383.4]
  wire [31:0] _T_432; // @[Math.scala 406:49:@27398.4]
  wire [31:0] _T_434; // @[Math.scala 406:56:@27400.4]
  wire [31:0] _T_435; // @[Math.scala 406:56:@27401.4]
  wire [31:0] _T_439; // @[package.scala 96:25:@27409.4]
  wire [31:0] x486_sum_number; // @[Math.scala 154:22:@27421.4 Math.scala 155:14:@27422.4]
  wire  _T_447; // @[FixedPoint.scala 50:25:@27426.4]
  wire [1:0] _T_451; // @[Bitwise.scala 72:12:@27428.4]
  wire [29:0] _T_452; // @[FixedPoint.scala 18:52:@27429.4]
  wire [31:0] _T_461; // @[Math.scala 406:49:@27437.4]
  wire [31:0] _T_463; // @[Math.scala 406:56:@27439.4]
  wire [31:0] _T_464; // @[Math.scala 406:56:@27440.4]
  wire [31:0] x489_sum_number; // @[Math.scala 154:22:@27451.4 Math.scala 155:14:@27452.4]
  wire [31:0] _T_474; // @[Math.scala 465:37:@27457.4]
  wire  x564_x490_D1; // @[package.scala 96:25:@27495.4 package.scala 96:25:@27496.4]
  wire [31:0] x565_x489_sum_D1_number; // @[package.scala 96:25:@27504.4 package.scala 96:25:@27505.4]
  wire [31:0] x492_sub_number; // @[Math.scala 195:22:@27477.4 Math.scala 196:14:@27478.4]
  wire  _T_506; // @[FixedPoint.scala 50:25:@27512.4]
  wire [1:0] _T_510; // @[Bitwise.scala 72:12:@27514.4]
  wire [29:0] _T_511; // @[FixedPoint.scala 18:52:@27515.4]
  wire [31:0] x321_number; // @[Cat.scala 30:58:@27516.4]
  wire [40:0] _GEN_0; // @[Math.scala 450:32:@27521.4]
  wire [40:0] _T_516; // @[Math.scala 450:32:@27521.4]
  wire [38:0] _GEN_1; // @[Math.scala 450:32:@27526.4]
  wire [38:0] _T_520; // @[Math.scala 450:32:@27526.4]
  wire  _T_553; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 179:149:@27615.4]
  wire  _T_557; // @[package.scala 96:25:@27623.4 package.scala 96:25:@27624.4]
  wire  _T_559; // @[implicits.scala 55:10:@27625.4]
  wire  _T_560; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 179:166:@27626.4]
  wire  _T_562; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 179:255:@27628.4]
  wire  _T_563; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 179:274:@27629.4]
  wire  x568_b307_D21; // @[package.scala 96:25:@27585.4 package.scala 96:25:@27586.4]
  wire  _T_564; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 179:300:@27630.4]
  wire  x567_b308_D21; // @[package.scala 96:25:@27576.4 package.scala 96:25:@27577.4]
  wire [31:0] x572_b305_D23_number; // @[package.scala 96:25:@27644.4 package.scala 96:25:@27645.4]
  wire [31:0] _T_578; // @[Math.scala 406:49:@27653.4]
  wire [31:0] _T_580; // @[Math.scala 406:56:@27655.4]
  wire [31:0] _T_581; // @[Math.scala 406:56:@27656.4]
  wire [31:0] _T_585; // @[package.scala 96:25:@27664.4]
  wire [31:0] x497_number; // @[implicits.scala 133:21:@27666.4]
  wire [31:0] x573_b306_D23_number; // @[package.scala 96:25:@27689.4 package.scala 96:25:@27690.4]
  wire [31:0] _T_605; // @[Math.scala 465:37:@27695.4]
  wire  x328; // @[package.scala 96:25:@27680.4 package.scala 96:25:@27681.4]
  wire  x329; // @[package.scala 96:25:@27703.4 package.scala 96:25:@27704.4]
  wire  x330; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 194:24:@27707.4]
  wire [31:0] _T_621; // @[Math.scala 406:49:@27716.4]
  wire [31:0] _T_623; // @[Math.scala 406:56:@27718.4]
  wire [31:0] _T_624; // @[Math.scala 406:56:@27719.4]
  wire  _T_629; // @[FixedPoint.scala 50:25:@27725.4]
  wire [1:0] _T_633; // @[Bitwise.scala 72:12:@27727.4]
  wire [29:0] _T_634; // @[FixedPoint.scala 18:52:@27728.4]
  wire [31:0] x333_number; // @[Cat.scala 30:58:@27729.4]
  wire [40:0] _GEN_2; // @[Math.scala 450:32:@27734.4]
  wire [40:0] _T_639; // @[Math.scala 450:32:@27734.4]
  wire [38:0] _GEN_3; // @[Math.scala 450:32:@27739.4]
  wire [38:0] _T_643; // @[Math.scala 450:32:@27739.4]
  wire  _T_685; // @[package.scala 96:25:@27843.4 package.scala 96:25:@27844.4]
  wire  _T_687; // @[implicits.scala 55:10:@27845.4]
  wire  _T_688; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 229:194:@27846.4]
  wire  x581_x331_D21; // @[package.scala 96:25:@27831.4 package.scala 96:25:@27832.4]
  wire  _T_689; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 229:283:@27847.4]
  wire  x577_b307_D45; // @[package.scala 96:25:@27795.4 package.scala 96:25:@27796.4]
  wire  _T_690; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 229:291:@27848.4]
  wire  x576_b308_D45; // @[package.scala 96:25:@27786.4 package.scala 96:25:@27787.4]
  wire [31:0] x338_rdcol_number; // @[Math.scala 195:22:@27867.4 Math.scala 196:14:@27868.4]
  wire [31:0] _T_705; // @[Math.scala 465:37:@27873.4]
  wire  x582_x328_D1; // @[package.scala 96:25:@27890.4 package.scala 96:25:@27891.4]
  wire  x339; // @[package.scala 96:25:@27881.4 package.scala 96:25:@27882.4]
  wire  x340; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 239:24:@27894.4]
  wire  _T_720; // @[FixedPoint.scala 50:25:@27901.4]
  wire [15:0] _T_724; // @[Bitwise.scala 72:12:@27903.4]
  wire [15:0] _T_725; // @[FixedPoint.scala 18:52:@27904.4]
  wire [31:0] _T_738; // @[Math.scala 406:56:@27921.4]
  wire [31:0] _T_739; // @[Math.scala 406:56:@27922.4]
  wire [31:0] _T_743; // @[package.scala 96:25:@27930.4]
  wire [31:0] x504_sum_number; // @[Math.scala 154:22:@27942.4 Math.scala 155:14:@27943.4]
  wire  _T_751; // @[FixedPoint.scala 50:25:@27947.4]
  wire [7:0] _T_755; // @[Bitwise.scala 72:12:@27949.4]
  wire [23:0] _T_756; // @[FixedPoint.scala 18:52:@27950.4]
  wire [31:0] _T_765; // @[Math.scala 406:49:@27958.4]
  wire [31:0] _T_767; // @[Math.scala 406:56:@27960.4]
  wire [31:0] _T_768; // @[Math.scala 406:56:@27961.4]
  wire [31:0] x507_sum_number; // @[Math.scala 154:22:@27972.4 Math.scala 155:14:@27973.4]
  wire  _T_776; // @[FixedPoint.scala 50:25:@27977.4]
  wire [3:0] _T_780; // @[Bitwise.scala 72:12:@27979.4]
  wire [27:0] _T_781; // @[FixedPoint.scala 18:52:@27980.4]
  wire [31:0] _T_790; // @[Math.scala 406:49:@27988.4]
  wire [31:0] _T_792; // @[Math.scala 406:56:@27990.4]
  wire [31:0] _T_793; // @[Math.scala 406:56:@27991.4]
  wire [31:0] x510_sum_number; // @[Math.scala 154:22:@28002.4 Math.scala 155:14:@28003.4]
  wire  _T_801; // @[FixedPoint.scala 50:25:@28007.4]
  wire [1:0] _T_805; // @[Bitwise.scala 72:12:@28009.4]
  wire [29:0] _T_806; // @[FixedPoint.scala 18:52:@28010.4]
  wire [31:0] _T_815; // @[Math.scala 406:49:@28018.4]
  wire [31:0] _T_817; // @[Math.scala 406:56:@28020.4]
  wire [31:0] _T_818; // @[Math.scala 406:56:@28021.4]
  wire [31:0] x513_sum_number; // @[Math.scala 154:22:@28032.4 Math.scala 155:14:@28033.4]
  wire  _T_826; // @[FixedPoint.scala 50:25:@28037.4]
  wire [1:0] _T_830; // @[Bitwise.scala 72:12:@28039.4]
  wire [29:0] _T_831; // @[FixedPoint.scala 18:52:@28040.4]
  wire [31:0] _T_840; // @[Math.scala 406:49:@28048.4]
  wire [31:0] _T_842; // @[Math.scala 406:56:@28050.4]
  wire [31:0] _T_843; // @[Math.scala 406:56:@28051.4]
  wire [31:0] x516_sum_number; // @[Math.scala 154:22:@28062.4 Math.scala 155:14:@28063.4]
  wire  _T_851; // @[FixedPoint.scala 50:25:@28067.4]
  wire [1:0] _T_855; // @[Bitwise.scala 72:12:@28069.4]
  wire [29:0] _T_856; // @[FixedPoint.scala 18:52:@28070.4]
  wire [31:0] _T_867; // @[Math.scala 406:49:@28085.4]
  wire [31:0] _T_869; // @[Math.scala 406:56:@28087.4]
  wire [31:0] _T_870; // @[Math.scala 406:56:@28088.4]
  wire [31:0] _T_874; // @[package.scala 96:25:@28096.4]
  wire [31:0] x519_sum_number; // @[Math.scala 154:22:@28108.4 Math.scala 155:14:@28109.4]
  wire [31:0] _T_886; // @[Math.scala 465:37:@28116.4]
  wire  x584_x520_D1; // @[package.scala 96:25:@28154.4 package.scala 96:25:@28155.4]
  wire [31:0] x585_x519_sum_D1_number; // @[package.scala 96:25:@28163.4 package.scala 96:25:@28164.4]
  wire [31:0] x522_sub_number; // @[Math.scala 195:22:@28136.4 Math.scala 196:14:@28137.4]
  wire  _T_945; // @[package.scala 96:25:@28227.4 package.scala 96:25:@28228.4]
  wire  _T_947; // @[implicits.scala 55:10:@28229.4]
  wire  _T_948; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 314:194:@28230.4]
  wire  x588_x341_D20; // @[package.scala 96:25:@28215.4 package.scala 96:25:@28216.4]
  wire  _T_949; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 314:283:@28231.4]
  wire  _T_950; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 314:291:@28232.4]
  wire [31:0] x347_rdcol_number; // @[Math.scala 195:22:@28251.4 Math.scala 196:14:@28252.4]
  wire [31:0] _T_965; // @[Math.scala 465:37:@28257.4]
  wire  x348; // @[package.scala 96:25:@28265.4 package.scala 96:25:@28266.4]
  wire  x349; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 322:59:@28269.4]
  wire  _T_977; // @[FixedPoint.scala 50:25:@28276.4]
  wire [15:0] _T_981; // @[Bitwise.scala 72:12:@28278.4]
  wire [15:0] _T_982; // @[FixedPoint.scala 18:52:@28279.4]
  wire [31:0] _T_995; // @[Math.scala 406:56:@28296.4]
  wire [31:0] _T_996; // @[Math.scala 406:56:@28297.4]
  wire [31:0] _T_1000; // @[package.scala 96:25:@28305.4]
  wire [31:0] x526_sum_number; // @[Math.scala 154:22:@28317.4 Math.scala 155:14:@28318.4]
  wire  _T_1008; // @[FixedPoint.scala 50:25:@28322.4]
  wire [7:0] _T_1012; // @[Bitwise.scala 72:12:@28324.4]
  wire [23:0] _T_1013; // @[FixedPoint.scala 18:52:@28325.4]
  wire [31:0] _T_1022; // @[Math.scala 406:49:@28333.4]
  wire [31:0] _T_1024; // @[Math.scala 406:56:@28335.4]
  wire [31:0] _T_1025; // @[Math.scala 406:56:@28336.4]
  wire [31:0] x529_sum_number; // @[Math.scala 154:22:@28347.4 Math.scala 155:14:@28348.4]
  wire  _T_1033; // @[FixedPoint.scala 50:25:@28352.4]
  wire [3:0] _T_1037; // @[Bitwise.scala 72:12:@28354.4]
  wire [27:0] _T_1038; // @[FixedPoint.scala 18:52:@28355.4]
  wire [31:0] _T_1047; // @[Math.scala 406:49:@28363.4]
  wire [31:0] _T_1049; // @[Math.scala 406:56:@28365.4]
  wire [31:0] _T_1050; // @[Math.scala 406:56:@28366.4]
  wire [31:0] x532_sum_number; // @[Math.scala 154:22:@28377.4 Math.scala 155:14:@28378.4]
  wire  _T_1058; // @[FixedPoint.scala 50:25:@28382.4]
  wire [1:0] _T_1062; // @[Bitwise.scala 72:12:@28384.4]
  wire [29:0] _T_1063; // @[FixedPoint.scala 18:52:@28385.4]
  wire [31:0] _T_1072; // @[Math.scala 406:49:@28393.4]
  wire [31:0] _T_1074; // @[Math.scala 406:56:@28395.4]
  wire [31:0] _T_1075; // @[Math.scala 406:56:@28396.4]
  wire [31:0] x535_sum_number; // @[Math.scala 154:22:@28407.4 Math.scala 155:14:@28408.4]
  wire  _T_1083; // @[FixedPoint.scala 50:25:@28412.4]
  wire [1:0] _T_1087; // @[Bitwise.scala 72:12:@28414.4]
  wire [29:0] _T_1088; // @[FixedPoint.scala 18:52:@28415.4]
  wire [31:0] _T_1097; // @[Math.scala 406:49:@28423.4]
  wire [31:0] _T_1099; // @[Math.scala 406:56:@28425.4]
  wire [31:0] _T_1100; // @[Math.scala 406:56:@28426.4]
  wire [31:0] x538_sum_number; // @[Math.scala 154:22:@28437.4 Math.scala 155:14:@28438.4]
  wire  _T_1108; // @[FixedPoint.scala 50:25:@28442.4]
  wire [1:0] _T_1112; // @[Bitwise.scala 72:12:@28444.4]
  wire [29:0] _T_1113; // @[FixedPoint.scala 18:52:@28445.4]
  wire [31:0] _T_1124; // @[Math.scala 406:49:@28460.4]
  wire [31:0] _T_1126; // @[Math.scala 406:56:@28462.4]
  wire [31:0] _T_1127; // @[Math.scala 406:56:@28463.4]
  wire [31:0] _T_1131; // @[package.scala 96:25:@28471.4]
  wire [31:0] x541_sum_number; // @[Math.scala 154:22:@28483.4 Math.scala 155:14:@28484.4]
  wire [31:0] _T_1141; // @[Math.scala 465:37:@28489.4]
  wire  x591_x542_D1; // @[package.scala 96:25:@28536.4 package.scala 96:25:@28537.4]
  wire [31:0] x590_x541_sum_D1_number; // @[package.scala 96:25:@28527.4 package.scala 96:25:@28528.4]
  wire [31:0] x544_sub_number; // @[Math.scala 195:22:@28509.4 Math.scala 196:14:@28510.4]
  wire  _T_1197; // @[package.scala 96:25:@28591.4 package.scala 96:25:@28592.4]
  wire  _T_1199; // @[implicits.scala 55:10:@28593.4]
  wire  _T_1200; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 387:194:@28594.4]
  wire  x593_x350_D20; // @[package.scala 96:25:@28579.4 package.scala 96:25:@28580.4]
  wire  _T_1201; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 387:283:@28595.4]
  wire  _T_1202; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 387:291:@28596.4]
  wire [31:0] x356_rdrow_number; // @[Math.scala 195:22:@28617.4 Math.scala 196:14:@28618.4]
  wire [31:0] _T_1221; // @[Math.scala 406:49:@28624.4]
  wire [31:0] _T_1223; // @[Math.scala 406:56:@28626.4]
  wire [31:0] _T_1224; // @[Math.scala 406:56:@28627.4]
  wire [31:0] _T_1228; // @[package.scala 96:25:@28635.4]
  wire [31:0] x546_number; // @[implicits.scala 133:21:@28637.4]
  wire  x358; // @[package.scala 96:25:@28651.4 package.scala 96:25:@28652.4]
  wire  x594_x329_D1; // @[package.scala 96:25:@28660.4 package.scala 96:25:@28661.4]
  wire  x359; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 407:24:@28664.4]
  wire [31:0] _T_1254; // @[Math.scala 406:49:@28673.4]
  wire [31:0] _T_1256; // @[Math.scala 406:56:@28675.4]
  wire [31:0] _T_1257; // @[Math.scala 406:56:@28676.4]
  wire  _T_1262; // @[FixedPoint.scala 50:25:@28682.4]
  wire [1:0] _T_1266; // @[Bitwise.scala 72:12:@28684.4]
  wire [29:0] _T_1267; // @[FixedPoint.scala 18:52:@28685.4]
  wire [31:0] x362_number; // @[Cat.scala 30:58:@28686.4]
  wire [40:0] _GEN_4; // @[Math.scala 450:32:@28691.4]
  wire [40:0] _T_1272; // @[Math.scala 450:32:@28691.4]
  wire [38:0] _GEN_5; // @[Math.scala 450:32:@28696.4]
  wire [38:0] _T_1276; // @[Math.scala 450:32:@28696.4]
  wire  _T_1306; // @[package.scala 96:25:@28764.4 package.scala 96:25:@28765.4]
  wire  _T_1308; // @[implicits.scala 55:10:@28766.4]
  wire  _T_1309; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 434:194:@28767.4]
  wire  x597_x360_D20; // @[package.scala 96:25:@28743.4 package.scala 96:25:@28744.4]
  wire  _T_1310; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 434:283:@28768.4]
  wire  _T_1311; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 434:291:@28769.4]
  wire  x367; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 438:24:@28780.4]
  wire  _T_1338; // @[package.scala 96:25:@28822.4 package.scala 96:25:@28823.4]
  wire  _T_1340; // @[implicits.scala 55:10:@28824.4]
  wire  _T_1341; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 451:194:@28825.4]
  wire  x600_x368_D20; // @[package.scala 96:25:@28810.4 package.scala 96:25:@28811.4]
  wire  _T_1342; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 451:283:@28826.4]
  wire  _T_1343; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 451:291:@28827.4]
  wire  x372; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 455:24:@28838.4]
  wire  _T_1367; // @[package.scala 96:25:@28871.4 package.scala 96:25:@28872.4]
  wire  _T_1369; // @[implicits.scala 55:10:@28873.4]
  wire  _T_1370; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 466:194:@28874.4]
  wire  x601_x373_D20; // @[package.scala 96:25:@28859.4 package.scala 96:25:@28860.4]
  wire  _T_1371; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 466:283:@28875.4]
  wire  _T_1372; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 466:291:@28876.4]
  wire [31:0] x377_rdrow_number; // @[Math.scala 195:22:@28895.4 Math.scala 196:14:@28896.4]
  wire [31:0] _T_1389; // @[Math.scala 406:49:@28902.4]
  wire [31:0] _T_1391; // @[Math.scala 406:56:@28904.4]
  wire [31:0] _T_1392; // @[Math.scala 406:56:@28905.4]
  wire [31:0] _T_1396; // @[package.scala 96:25:@28913.4]
  wire [31:0] x551_number; // @[implicits.scala 133:21:@28915.4]
  wire  x379; // @[package.scala 96:25:@28929.4 package.scala 96:25:@28930.4]
  wire  x380; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 476:24:@28933.4]
  wire [31:0] _T_1419; // @[Math.scala 406:49:@28942.4]
  wire [31:0] _T_1421; // @[Math.scala 406:56:@28944.4]
  wire [31:0] _T_1422; // @[Math.scala 406:56:@28945.4]
  wire  _T_1427; // @[FixedPoint.scala 50:25:@28951.4]
  wire [1:0] _T_1431; // @[Bitwise.scala 72:12:@28953.4]
  wire [29:0] _T_1432; // @[FixedPoint.scala 18:52:@28954.4]
  wire [31:0] x383_number; // @[Cat.scala 30:58:@28955.4]
  wire [40:0] _GEN_6; // @[Math.scala 450:32:@28960.4]
  wire [40:0] _T_1437; // @[Math.scala 450:32:@28960.4]
  wire [38:0] _GEN_7; // @[Math.scala 450:32:@28965.4]
  wire [38:0] _T_1441; // @[Math.scala 450:32:@28965.4]
  wire  _T_1471; // @[package.scala 96:25:@29033.4 package.scala 96:25:@29034.4]
  wire  _T_1473; // @[implicits.scala 55:10:@29035.4]
  wire  _T_1474; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 503:194:@29036.4]
  wire  x604_x381_D20; // @[package.scala 96:25:@29012.4 package.scala 96:25:@29013.4]
  wire  _T_1475; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 503:283:@29037.4]
  wire  _T_1476; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 503:291:@29038.4]
  wire  x388; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 507:24:@29049.4]
  wire  _T_1505; // @[package.scala 96:25:@29093.4 package.scala 96:25:@29094.4]
  wire  _T_1507; // @[implicits.scala 55:10:@29095.4]
  wire  _T_1508; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 528:194:@29096.4]
  wire  x607_x389_D20; // @[package.scala 96:25:@29081.4 package.scala 96:25:@29082.4]
  wire  _T_1509; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 528:283:@29097.4]
  wire  _T_1510; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 528:291:@29098.4]
  wire  x393; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 532:59:@29109.4]
  wire  _T_1534; // @[package.scala 96:25:@29142.4 package.scala 96:25:@29143.4]
  wire  _T_1536; // @[implicits.scala 55:10:@29144.4]
  wire  _T_1537; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 543:194:@29145.4]
  wire  x608_x394_D20; // @[package.scala 96:25:@29130.4 package.scala 96:25:@29131.4]
  wire  _T_1538; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 543:283:@29146.4]
  wire  _T_1539; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 543:291:@29147.4]
  wire [7:0] x345_rd_0_number; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 310:29:@28218.4 sm_x416_inr_Foreach_SAMPLER_BOX.scala 314:408:@28239.4]
  wire [8:0] _GEN_8; // @[Math.scala 450:32:@29159.4]
  wire [7:0] x365_rd_0_number; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 430:29:@28755.4 sm_x416_inr_Foreach_SAMPLER_BOX.scala 434:408:@28776.4]
  wire [8:0] _GEN_9; // @[Math.scala 450:32:@29171.4]
  wire [7:0] x370_rd_0_number; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 447:29:@28813.4 sm_x416_inr_Foreach_SAMPLER_BOX.scala 451:408:@28834.4]
  wire [9:0] _GEN_10; // @[Math.scala 450:32:@29183.4]
  wire [7:0] x375_rd_0_number; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 462:29:@28862.4 sm_x416_inr_Foreach_SAMPLER_BOX.scala 466:408:@28883.4]
  wire [8:0] _GEN_11; // @[Math.scala 450:32:@29195.4]
  wire [7:0] x391_rd_0_number; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 524:29:@29084.4 sm_x416_inr_Foreach_SAMPLER_BOX.scala 528:408:@29105.4]
  wire [8:0] _GEN_12; // @[Math.scala 450:32:@29207.4]
  wire [7:0] x410_sum_number; // @[Math.scala 154:22:@29330.4 Math.scala 155:14:@29331.4]
  wire [3:0] _T_1616; // @[FixedPoint.scala 18:52:@29336.4]
  wire  _T_1637; // @[package.scala 96:25:@29377.4 package.scala 96:25:@29378.4]
  wire  _T_1639; // @[implicits.scala 55:10:@29379.4]
  wire  x613_b307_D52; // @[package.scala 96:25:@29359.4 package.scala 96:25:@29360.4]
  wire  _T_1640; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 591:117:@29380.4]
  wire  x614_b308_D52; // @[package.scala 96:25:@29368.4 package.scala 96:25:@29369.4]
  wire  _T_1641; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 591:123:@29381.4]
  wire [31:0] x324_sum_number; // @[Math.scala 154:22:@27567.4 Math.scala 155:14:@27568.4]
  wire [31:0] x569_x493_D13_number; // @[package.scala 96:25:@27594.4 package.scala 96:25:@27595.4]
  wire [31:0] x570_x471_D19_number; // @[package.scala 96:25:@27603.4 package.scala 96:25:@27604.4]
  wire [31:0] x578_x493_D37_number; // @[package.scala 96:25:@27804.4 package.scala 96:25:@27805.4]
  wire [31:0] x579_x498_D21_number; // @[package.scala 96:25:@27813.4 package.scala 96:25:@27814.4]
  wire [31:0] x580_x335_sum_D1_number; // @[package.scala 96:25:@27822.4 package.scala 96:25:@27823.4]
  wire [31:0] x344_sum_number; // @[Math.scala 154:22:@28197.4 Math.scala 155:14:@28198.4]
  wire [31:0] x587_x523_D12_number; // @[package.scala 96:25:@28206.4 package.scala 96:25:@28207.4]
  wire [31:0] x353_sum_number; // @[Math.scala 154:22:@28561.4 Math.scala 155:14:@28562.4]
  wire [31:0] x592_x545_D12_number; // @[package.scala 96:25:@28570.4 package.scala 96:25:@28571.4]
  wire [31:0] x596_x547_D20_number; // @[package.scala 96:25:@28734.4 package.scala 96:25:@28735.4]
  wire [31:0] x598_x364_sum_D1_number; // @[package.scala 96:25:@28752.4 package.scala 96:25:@28753.4]
  wire [31:0] x369_sum_number; // @[Math.scala 154:22:@28801.4 Math.scala 155:14:@28802.4]
  wire [31:0] x374_sum_number; // @[Math.scala 154:22:@28850.4 Math.scala 155:14:@28851.4]
  wire [31:0] x603_x385_sum_D1_number; // @[package.scala 96:25:@29003.4 package.scala 96:25:@29004.4]
  wire [31:0] x605_x552_D20_number; // @[package.scala 96:25:@29021.4 package.scala 96:25:@29022.4]
  wire [31:0] x390_sum_number; // @[Math.scala 154:22:@29072.4 Math.scala 155:14:@29073.4]
  wire [31:0] x395_sum_number; // @[Math.scala 154:22:@29121.4 Math.scala 155:14:@29122.4]
  wire [8:0] _T_1547; // @[package.scala 96:25:@29165.4 package.scala 96:25:@29166.4]
  wire [8:0] _T_1553; // @[package.scala 96:25:@29177.4 package.scala 96:25:@29178.4]
  wire [9:0] _T_1559; // @[package.scala 96:25:@29189.4 package.scala 96:25:@29190.4]
  wire [8:0] _T_1565; // @[package.scala 96:25:@29201.4 package.scala 96:25:@29202.4]
  wire [8:0] _T_1571; // @[package.scala 96:25:@29213.4 package.scala 96:25:@29214.4]
  _ _ ( // @[Math.scala 709:24:@27072.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 709:24:@27084.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  RetimeWrapper_50 RetimeWrapper ( // @[package.scala 93:22:@27107.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x311_lb_0 x311_lb_0 ( // @[m_x311_lb_0.scala 35:17:@27117.4]
    .clock(x311_lb_0_clock),
    .reset(x311_lb_0_reset),
    .io_rPort_8_banks_1(x311_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x311_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x311_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x311_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x311_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x311_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x311_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x311_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x311_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x311_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x311_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x311_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x311_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x311_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x311_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x311_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x311_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x311_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x311_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x311_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x311_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x311_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x311_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x311_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x311_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x311_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x311_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x311_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x311_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x311_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x311_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x311_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x311_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x311_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x311_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x311_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x311_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x311_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x311_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x311_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x311_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x311_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x311_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x311_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x311_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x311_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x311_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x311_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x311_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x311_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x311_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x311_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x311_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x311_lb_0_io_rPort_0_output_0),
    .io_wPort_0_banks_1(x311_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x311_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x311_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x311_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x311_lb_0_io_wPort_0_en_0)
  );
  RetimeWrapper_171 RetimeWrapper_1 ( // @[package.scala 93:22:@27239.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x292_sum x474_sum_1 ( // @[Math.scala 150:24:@27279.4]
    .clock(x474_sum_1_clock),
    .reset(x474_sum_1_reset),
    .io_a(x474_sum_1_io_a),
    .io_b(x474_sum_1_io_b),
    .io_flow(x474_sum_1_io_flow),
    .io_result(x474_sum_1_io_result)
  );
  x292_sum x477_sum_1 ( // @[Math.scala 150:24:@27309.4]
    .clock(x477_sum_1_clock),
    .reset(x477_sum_1_reset),
    .io_a(x477_sum_1_io_a),
    .io_b(x477_sum_1_io_b),
    .io_flow(x477_sum_1_io_flow),
    .io_result(x477_sum_1_io_result)
  );
  x292_sum x480_sum_1 ( // @[Math.scala 150:24:@27339.4]
    .clock(x480_sum_1_clock),
    .reset(x480_sum_1_reset),
    .io_a(x480_sum_1_io_a),
    .io_b(x480_sum_1_io_b),
    .io_flow(x480_sum_1_io_flow),
    .io_result(x480_sum_1_io_result)
  );
  x292_sum x483_sum_1 ( // @[Math.scala 150:24:@27369.4]
    .clock(x483_sum_1_clock),
    .reset(x483_sum_1_reset),
    .io_a(x483_sum_1_io_a),
    .io_b(x483_sum_1_io_b),
    .io_flow(x483_sum_1_io_flow),
    .io_result(x483_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_2 ( // @[package.scala 93:22:@27385.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_3 ( // @[package.scala 93:22:@27402.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x292_sum x486_sum_1 ( // @[Math.scala 150:24:@27415.4]
    .clock(x486_sum_1_clock),
    .reset(x486_sum_1_reset),
    .io_a(x486_sum_1_io_a),
    .io_b(x486_sum_1_io_b),
    .io_flow(x486_sum_1_io_flow),
    .io_result(x486_sum_1_io_result)
  );
  x292_sum x489_sum_1 ( // @[Math.scala 150:24:@27445.4]
    .clock(x489_sum_1_clock),
    .reset(x489_sum_1_reset),
    .io_a(x489_sum_1_io_a),
    .io_b(x489_sum_1_io_b),
    .io_flow(x489_sum_1_io_flow),
    .io_result(x489_sum_1_io_result)
  );
  x467_sub x492_sub_1 ( // @[Math.scala 191:24:@27471.4]
    .clock(x492_sub_1_clock),
    .reset(x492_sub_1_reset),
    .io_a(x492_sub_1_io_a),
    .io_b(x492_sub_1_io_b),
    .io_flow(x492_sub_1_io_flow),
    .io_result(x492_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@27481.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@27490.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_6 ( // @[package.scala 93:22:@27499.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x292_sum x496_sum_1 ( // @[Math.scala 150:24:@27530.4]
    .clock(x496_sum_1_clock),
    .reset(x496_sum_1_reset),
    .io_a(x496_sum_1_io_a),
    .io_b(x496_sum_1_io_b),
    .io_flow(x496_sum_1_io_flow),
    .io_result(x496_sum_1_io_result)
  );
  x323_div x323_div_1 ( // @[Math.scala 327:24:@27542.4]
    .clock(x323_div_1_clock),
    .reset(x323_div_1_reset),
    .io_a(x323_div_1_io_a),
    .io_flow(x323_div_1_io_flow),
    .io_result(x323_div_1_io_result)
  );
  RetimeWrapper_186 RetimeWrapper_7 ( // @[package.scala 93:22:@27552.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  x292_sum x324_sum_1 ( // @[Math.scala 150:24:@27561.4]
    .clock(x324_sum_1_clock),
    .reset(x324_sum_1_reset),
    .io_a(x324_sum_1_io_a),
    .io_b(x324_sum_1_io_b),
    .io_flow(x324_sum_1_io_flow),
    .io_result(x324_sum_1_io_result)
  );
  RetimeWrapper_188 RetimeWrapper_8 ( // @[package.scala 93:22:@27571.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_188 RetimeWrapper_9 ( // @[package.scala 93:22:@27580.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_190 RetimeWrapper_10 ( // @[package.scala 93:22:@27589.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_191 RetimeWrapper_11 ( // @[package.scala 93:22:@27598.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_192 RetimeWrapper_12 ( // @[package.scala 93:22:@27607.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_188 RetimeWrapper_13 ( // @[package.scala 93:22:@27618.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_194 RetimeWrapper_14 ( // @[package.scala 93:22:@27639.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_15 ( // @[package.scala 93:22:@27657.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper RetimeWrapper_16 ( // @[package.scala 93:22:@27675.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_194 RetimeWrapper_17 ( // @[package.scala 93:22:@27684.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper RetimeWrapper_18 ( // @[package.scala 93:22:@27698.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  x292_sum x501_sum_1 ( // @[Math.scala 150:24:@27743.4]
    .clock(x501_sum_1_clock),
    .reset(x501_sum_1_reset),
    .io_a(x501_sum_1_io_a),
    .io_b(x501_sum_1_io_b),
    .io_flow(x501_sum_1_io_flow),
    .io_result(x501_sum_1_io_result)
  );
  RetimeWrapper_200 RetimeWrapper_19 ( // @[package.scala 93:22:@27753.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_194 RetimeWrapper_20 ( // @[package.scala 93:22:@27762.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  x292_sum x335_sum_1 ( // @[Math.scala 150:24:@27771.4]
    .clock(x335_sum_1_clock),
    .reset(x335_sum_1_reset),
    .io_a(x335_sum_1_io_a),
    .io_b(x335_sum_1_io_b),
    .io_flow(x335_sum_1_io_flow),
    .io_result(x335_sum_1_io_result)
  );
  RetimeWrapper_203 RetimeWrapper_21 ( // @[package.scala 93:22:@27781.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_203 RetimeWrapper_22 ( // @[package.scala 93:22:@27790.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_205 RetimeWrapper_23 ( // @[package.scala 93:22:@27799.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_206 RetimeWrapper_24 ( // @[package.scala 93:22:@27808.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_25 ( // @[package.scala 93:22:@27817.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_188 RetimeWrapper_26 ( // @[package.scala 93:22:@27826.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_203 RetimeWrapper_27 ( // @[package.scala 93:22:@27838.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  x467_sub x338_rdcol_1 ( // @[Math.scala 191:24:@27861.4]
    .clock(x338_rdcol_1_clock),
    .reset(x338_rdcol_1_reset),
    .io_a(x338_rdcol_1_io_a),
    .io_b(x338_rdcol_1_io_b),
    .io_flow(x338_rdcol_1_io_flow),
    .io_result(x338_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_28 ( // @[package.scala 93:22:@27876.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper RetimeWrapper_29 ( // @[package.scala 93:22:@27885.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_30 ( // @[package.scala 93:22:@27906.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_31 ( // @[package.scala 93:22:@27923.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  x292_sum x504_sum_1 ( // @[Math.scala 150:24:@27936.4]
    .clock(x504_sum_1_clock),
    .reset(x504_sum_1_reset),
    .io_a(x504_sum_1_io_a),
    .io_b(x504_sum_1_io_b),
    .io_flow(x504_sum_1_io_flow),
    .io_result(x504_sum_1_io_result)
  );
  x292_sum x507_sum_1 ( // @[Math.scala 150:24:@27966.4]
    .clock(x507_sum_1_clock),
    .reset(x507_sum_1_reset),
    .io_a(x507_sum_1_io_a),
    .io_b(x507_sum_1_io_b),
    .io_flow(x507_sum_1_io_flow),
    .io_result(x507_sum_1_io_result)
  );
  x292_sum x510_sum_1 ( // @[Math.scala 150:24:@27996.4]
    .clock(x510_sum_1_clock),
    .reset(x510_sum_1_reset),
    .io_a(x510_sum_1_io_a),
    .io_b(x510_sum_1_io_b),
    .io_flow(x510_sum_1_io_flow),
    .io_result(x510_sum_1_io_result)
  );
  x292_sum x513_sum_1 ( // @[Math.scala 150:24:@28026.4]
    .clock(x513_sum_1_clock),
    .reset(x513_sum_1_reset),
    .io_a(x513_sum_1_io_a),
    .io_b(x513_sum_1_io_b),
    .io_flow(x513_sum_1_io_flow),
    .io_result(x513_sum_1_io_result)
  );
  x292_sum x516_sum_1 ( // @[Math.scala 150:24:@28056.4]
    .clock(x516_sum_1_clock),
    .reset(x516_sum_1_reset),
    .io_a(x516_sum_1_io_a),
    .io_b(x516_sum_1_io_b),
    .io_flow(x516_sum_1_io_flow),
    .io_result(x516_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_32 ( // @[package.scala 93:22:@28072.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_33 ( // @[package.scala 93:22:@28089.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  x292_sum x519_sum_1 ( // @[Math.scala 150:24:@28102.4]
    .clock(x519_sum_1_clock),
    .reset(x519_sum_1_reset),
    .io_a(x519_sum_1_io_a),
    .io_b(x519_sum_1_io_b),
    .io_flow(x519_sum_1_io_flow),
    .io_result(x519_sum_1_io_result)
  );
  x467_sub x522_sub_1 ( // @[Math.scala 191:24:@28130.4]
    .clock(x522_sub_1_clock),
    .reset(x522_sub_1_reset),
    .io_a(x522_sub_1_io_a),
    .io_b(x522_sub_1_io_b),
    .io_flow(x522_sub_1_io_flow),
    .io_result(x522_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_34 ( // @[package.scala 93:22:@28140.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper RetimeWrapper_35 ( // @[package.scala 93:22:@28149.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_36 ( // @[package.scala 93:22:@28158.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  x323_div x343_div_1 ( // @[Math.scala 327:24:@28172.4]
    .clock(x343_div_1_clock),
    .reset(x343_div_1_reset),
    .io_a(x343_div_1_io_a),
    .io_flow(x343_div_1_io_flow),
    .io_result(x343_div_1_io_result)
  );
  RetimeWrapper_191 RetimeWrapper_37 ( // @[package.scala 93:22:@28182.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  x292_sum x344_sum_1 ( // @[Math.scala 150:24:@28191.4]
    .clock(x344_sum_1_clock),
    .reset(x344_sum_1_reset),
    .io_a(x344_sum_1_io_a),
    .io_b(x344_sum_1_io_b),
    .io_flow(x344_sum_1_io_flow),
    .io_result(x344_sum_1_io_result)
  );
  RetimeWrapper_230 RetimeWrapper_38 ( // @[package.scala 93:22:@28201.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_231 RetimeWrapper_39 ( // @[package.scala 93:22:@28210.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_203 RetimeWrapper_40 ( // @[package.scala 93:22:@28222.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  x467_sub x347_rdcol_1 ( // @[Math.scala 191:24:@28245.4]
    .clock(x347_rdcol_1_clock),
    .reset(x347_rdcol_1_reset),
    .io_a(x347_rdcol_1_io_a),
    .io_b(x347_rdcol_1_io_b),
    .io_flow(x347_rdcol_1_io_flow),
    .io_result(x347_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_41 ( // @[package.scala 93:22:@28260.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_42 ( // @[package.scala 93:22:@28281.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_43 ( // @[package.scala 93:22:@28298.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  x292_sum x526_sum_1 ( // @[Math.scala 150:24:@28311.4]
    .clock(x526_sum_1_clock),
    .reset(x526_sum_1_reset),
    .io_a(x526_sum_1_io_a),
    .io_b(x526_sum_1_io_b),
    .io_flow(x526_sum_1_io_flow),
    .io_result(x526_sum_1_io_result)
  );
  x292_sum x529_sum_1 ( // @[Math.scala 150:24:@28341.4]
    .clock(x529_sum_1_clock),
    .reset(x529_sum_1_reset),
    .io_a(x529_sum_1_io_a),
    .io_b(x529_sum_1_io_b),
    .io_flow(x529_sum_1_io_flow),
    .io_result(x529_sum_1_io_result)
  );
  x292_sum x532_sum_1 ( // @[Math.scala 150:24:@28371.4]
    .clock(x532_sum_1_clock),
    .reset(x532_sum_1_reset),
    .io_a(x532_sum_1_io_a),
    .io_b(x532_sum_1_io_b),
    .io_flow(x532_sum_1_io_flow),
    .io_result(x532_sum_1_io_result)
  );
  x292_sum x535_sum_1 ( // @[Math.scala 150:24:@28401.4]
    .clock(x535_sum_1_clock),
    .reset(x535_sum_1_reset),
    .io_a(x535_sum_1_io_a),
    .io_b(x535_sum_1_io_b),
    .io_flow(x535_sum_1_io_flow),
    .io_result(x535_sum_1_io_result)
  );
  x292_sum x538_sum_1 ( // @[Math.scala 150:24:@28431.4]
    .clock(x538_sum_1_clock),
    .reset(x538_sum_1_reset),
    .io_a(x538_sum_1_io_a),
    .io_b(x538_sum_1_io_b),
    .io_flow(x538_sum_1_io_flow),
    .io_result(x538_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_44 ( // @[package.scala 93:22:@28447.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_45 ( // @[package.scala 93:22:@28464.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  x292_sum x541_sum_1 ( // @[Math.scala 150:24:@28477.4]
    .clock(x541_sum_1_clock),
    .reset(x541_sum_1_reset),
    .io_a(x541_sum_1_io_a),
    .io_b(x541_sum_1_io_b),
    .io_flow(x541_sum_1_io_flow),
    .io_result(x541_sum_1_io_result)
  );
  x467_sub x544_sub_1 ( // @[Math.scala 191:24:@28503.4]
    .clock(x544_sub_1_clock),
    .reset(x544_sub_1_reset),
    .io_a(x544_sub_1_io_a),
    .io_b(x544_sub_1_io_b),
    .io_flow(x544_sub_1_io_flow),
    .io_result(x544_sub_1_io_result)
  );
  RetimeWrapper RetimeWrapper_46 ( // @[package.scala 93:22:@28513.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_47 ( // @[package.scala 93:22:@28522.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper RetimeWrapper_48 ( // @[package.scala 93:22:@28531.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  x323_div x352_div_1 ( // @[Math.scala 327:24:@28545.4]
    .clock(x352_div_1_clock),
    .reset(x352_div_1_reset),
    .io_a(x352_div_1_io_a),
    .io_flow(x352_div_1_io_flow),
    .io_result(x352_div_1_io_result)
  );
  x292_sum x353_sum_1 ( // @[Math.scala 150:24:@28555.4]
    .clock(x353_sum_1_clock),
    .reset(x353_sum_1_reset),
    .io_a(x353_sum_1_io_a),
    .io_b(x353_sum_1_io_b),
    .io_flow(x353_sum_1_io_flow),
    .io_result(x353_sum_1_io_result)
  );
  RetimeWrapper_230 RetimeWrapper_49 ( // @[package.scala 93:22:@28565.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_231 RetimeWrapper_50 ( // @[package.scala 93:22:@28574.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_203 RetimeWrapper_51 ( // @[package.scala 93:22:@28586.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  x467_sub x356_rdrow_1 ( // @[Math.scala 191:24:@28611.4]
    .clock(x356_rdrow_1_clock),
    .reset(x356_rdrow_1_reset),
    .io_a(x356_rdrow_1_io_a),
    .io_b(x356_rdrow_1_io_b),
    .io_flow(x356_rdrow_1_io_flow),
    .io_result(x356_rdrow_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_52 ( // @[package.scala 93:22:@28628.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper RetimeWrapper_53 ( // @[package.scala 93:22:@28646.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper RetimeWrapper_54 ( // @[package.scala 93:22:@28655.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  x292_sum x550_sum_1 ( // @[Math.scala 150:24:@28700.4]
    .clock(x550_sum_1_clock),
    .reset(x550_sum_1_reset),
    .io_a(x550_sum_1_io_a),
    .io_b(x550_sum_1_io_b),
    .io_flow(x550_sum_1_io_flow),
    .io_result(x550_sum_1_io_result)
  );
  RetimeWrapper_186 RetimeWrapper_55 ( // @[package.scala 93:22:@28710.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  x292_sum x364_sum_1 ( // @[Math.scala 150:24:@28719.4]
    .clock(x364_sum_1_clock),
    .reset(x364_sum_1_reset),
    .io_a(x364_sum_1_io_a),
    .io_b(x364_sum_1_io_b),
    .io_flow(x364_sum_1_io_flow),
    .io_result(x364_sum_1_io_result)
  );
  RetimeWrapper_185 RetimeWrapper_56 ( // @[package.scala 93:22:@28729.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_231 RetimeWrapper_57 ( // @[package.scala 93:22:@28738.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_58 ( // @[package.scala 93:22:@28747.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_203 RetimeWrapper_59 ( // @[package.scala 93:22:@28759.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_200 RetimeWrapper_60 ( // @[package.scala 93:22:@28786.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  x292_sum x369_sum_1 ( // @[Math.scala 150:24:@28795.4]
    .clock(x369_sum_1_clock),
    .reset(x369_sum_1_reset),
    .io_a(x369_sum_1_io_a),
    .io_b(x369_sum_1_io_b),
    .io_flow(x369_sum_1_io_flow),
    .io_result(x369_sum_1_io_result)
  );
  RetimeWrapper_231 RetimeWrapper_61 ( // @[package.scala 93:22:@28805.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_203 RetimeWrapper_62 ( // @[package.scala 93:22:@28817.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  x292_sum x374_sum_1 ( // @[Math.scala 150:24:@28844.4]
    .clock(x374_sum_1_clock),
    .reset(x374_sum_1_reset),
    .io_a(x374_sum_1_io_a),
    .io_b(x374_sum_1_io_b),
    .io_flow(x374_sum_1_io_flow),
    .io_result(x374_sum_1_io_result)
  );
  RetimeWrapper_231 RetimeWrapper_63 ( // @[package.scala 93:22:@28854.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_203 RetimeWrapper_64 ( // @[package.scala 93:22:@28866.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  x467_sub x377_rdrow_1 ( // @[Math.scala 191:24:@28889.4]
    .clock(x377_rdrow_1_clock),
    .reset(x377_rdrow_1_reset),
    .io_a(x377_rdrow_1_io_a),
    .io_b(x377_rdrow_1_io_b),
    .io_flow(x377_rdrow_1_io_flow),
    .io_result(x377_rdrow_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_65 ( // @[package.scala 93:22:@28906.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper RetimeWrapper_66 ( // @[package.scala 93:22:@28924.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  x292_sum x555_sum_1 ( // @[Math.scala 150:24:@28969.4]
    .clock(x555_sum_1_clock),
    .reset(x555_sum_1_reset),
    .io_a(x555_sum_1_io_a),
    .io_b(x555_sum_1_io_b),
    .io_flow(x555_sum_1_io_flow),
    .io_result(x555_sum_1_io_result)
  );
  RetimeWrapper_186 RetimeWrapper_67 ( // @[package.scala 93:22:@28979.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  x292_sum x385_sum_1 ( // @[Math.scala 150:24:@28988.4]
    .clock(x385_sum_1_clock),
    .reset(x385_sum_1_reset),
    .io_a(x385_sum_1_io_a),
    .io_b(x385_sum_1_io_b),
    .io_flow(x385_sum_1_io_flow),
    .io_result(x385_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_68 ( // @[package.scala 93:22:@28998.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_231 RetimeWrapper_69 ( // @[package.scala 93:22:@29007.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_185 RetimeWrapper_70 ( // @[package.scala 93:22:@29016.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_203 RetimeWrapper_71 ( // @[package.scala 93:22:@29028.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_200 RetimeWrapper_72 ( // @[package.scala 93:22:@29055.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  x292_sum x390_sum_1 ( // @[Math.scala 150:24:@29066.4]
    .clock(x390_sum_1_clock),
    .reset(x390_sum_1_reset),
    .io_a(x390_sum_1_io_a),
    .io_b(x390_sum_1_io_b),
    .io_flow(x390_sum_1_io_flow),
    .io_result(x390_sum_1_io_result)
  );
  RetimeWrapper_231 RetimeWrapper_73 ( // @[package.scala 93:22:@29076.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_203 RetimeWrapper_74 ( // @[package.scala 93:22:@29088.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  x292_sum x395_sum_1 ( // @[Math.scala 150:24:@29115.4]
    .clock(x395_sum_1_clock),
    .reset(x395_sum_1_reset),
    .io_a(x395_sum_1_io_a),
    .io_b(x395_sum_1_io_b),
    .io_flow(x395_sum_1_io_flow),
    .io_result(x395_sum_1_io_result)
  );
  RetimeWrapper_231 RetimeWrapper_75 ( // @[package.scala 93:22:@29125.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_203 RetimeWrapper_76 ( // @[package.scala 93:22:@29137.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_289 RetimeWrapper_77 ( // @[package.scala 93:22:@29160.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_289 RetimeWrapper_78 ( // @[package.scala 93:22:@29172.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_51 RetimeWrapper_79 ( // @[package.scala 93:22:@29184.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_289 RetimeWrapper_80 ( // @[package.scala 93:22:@29196.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_289 RetimeWrapper_81 ( // @[package.scala 93:22:@29208.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_50 RetimeWrapper_82 ( // @[package.scala 93:22:@29218.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  x403_x15 x403_x15_1 ( // @[Math.scala 150:24:@29227.4]
    .io_a(x403_x15_1_io_a),
    .io_b(x403_x15_1_io_b),
    .io_result(x403_x15_1_io_result)
  );
  RetimeWrapper_50 RetimeWrapper_83 ( // @[package.scala 93:22:@29237.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  x403_x15 x404_x16_1 ( // @[Math.scala 150:24:@29246.4]
    .io_a(x404_x16_1_io_a),
    .io_b(x404_x16_1_io_b),
    .io_result(x404_x16_1_io_result)
  );
  x403_x15 x405_x15_1 ( // @[Math.scala 150:24:@29256.4]
    .io_a(x405_x15_1_io_a),
    .io_b(x405_x15_1_io_b),
    .io_result(x405_x15_1_io_result)
  );
  RetimeWrapper_50 RetimeWrapper_84 ( // @[package.scala 93:22:@29266.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  x403_x15 x406_x16_1 ( // @[Math.scala 150:24:@29275.4]
    .io_a(x406_x16_1_io_a),
    .io_b(x406_x16_1_io_b),
    .io_result(x406_x16_1_io_result)
  );
  x403_x15 x407_x15_1 ( // @[Math.scala 150:24:@29285.4]
    .io_a(x407_x15_1_io_a),
    .io_b(x407_x15_1_io_b),
    .io_result(x407_x15_1_io_result)
  );
  x403_x15 x408_x16_1 ( // @[Math.scala 150:24:@29295.4]
    .io_a(x408_x16_1_io_a),
    .io_b(x408_x16_1_io_b),
    .io_result(x408_x16_1_io_result)
  );
  x403_x15 x409_x15_1 ( // @[Math.scala 150:24:@29305.4]
    .io_a(x409_x15_1_io_a),
    .io_b(x409_x15_1_io_b),
    .io_result(x409_x15_1_io_result)
  );
  RetimeWrapper_50 RetimeWrapper_85 ( // @[package.scala 93:22:@29315.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  x410_sum x410_sum_1 ( // @[Math.scala 150:24:@29324.4]
    .clock(x410_sum_1_clock),
    .reset(x410_sum_1_reset),
    .io_a(x410_sum_1_io_a),
    .io_b(x410_sum_1_io_b),
    .io_flow(x410_sum_1_io_flow),
    .io_result(x410_sum_1_io_result)
  );
  RetimeWrapper_299 RetimeWrapper_86 ( // @[package.scala 93:22:@29345.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_42 RetimeWrapper_87 ( // @[package.scala 93:22:@29354.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_42 RetimeWrapper_88 ( // @[package.scala 93:22:@29363.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_42 RetimeWrapper_89 ( // @[package.scala 93:22:@29372.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  assign b307 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 62:18:@27092.4]
  assign b308 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 63:18:@27093.4]
  assign _T_205 = b307 & b308; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 67:30:@27095.4]
  assign _T_206 = _T_205 & io_sigsIn_datapathEn; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 67:37:@27096.4]
  assign _T_210 = io_in_x278_TID == 8'h0; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 69:76:@27101.4]
  assign _T_211 = _T_206 & _T_210; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 69:62:@27102.4]
  assign _T_213 = io_in_x278_TDEST == 8'h0; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 69:101:@27103.4]
  assign b305_number = __io_result; // @[Math.scala 712:22:@27077.4 Math.scala 713:14:@27078.4]
  assign _T_240 = $signed(b305_number); // @[Math.scala 499:52:@27193.4]
  assign x314 = $signed(32'sh1) == $signed(_T_240); // @[Math.scala 499:44:@27201.4]
  assign x315 = $signed(32'sh2) == $signed(_T_240); // @[Math.scala 499:44:@27208.4]
  assign x316 = $signed(32'sh3) == $signed(_T_240); // @[Math.scala 499:44:@27215.4]
  assign _T_287 = x314 ? 32'h1 : 32'h0; // @[Mux.scala 19:72:@27227.4]
  assign _T_289 = x315 ? 32'h2 : 32'h0; // @[Mux.scala 19:72:@27228.4]
  assign _T_291 = x316 ? 32'h3 : 32'h0; // @[Mux.scala 19:72:@27229.4]
  assign _T_293 = _T_287 | _T_289; // @[Mux.scala 19:72:@27231.4]
  assign x562_x317_D2_number = RetimeWrapper_1_io_out; // @[package.scala 96:25:@27244.4 package.scala 96:25:@27245.4]
  assign _T_308 = $signed(x562_x317_D2_number); // @[Math.scala 406:49:@27251.4]
  assign _T_310 = $signed(_T_308) & $signed(32'sh3); // @[Math.scala 406:56:@27253.4]
  assign _T_311 = $signed(_T_310); // @[Math.scala 406:56:@27254.4]
  assign b306_number = __1_io_result; // @[Math.scala 712:22:@27089.4 Math.scala 713:14:@27090.4]
  assign _T_316 = b306_number[31]; // @[FixedPoint.scala 50:25:@27260.4]
  assign _T_320 = _T_316 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@27262.4]
  assign _T_321 = b306_number[31:16]; // @[FixedPoint.scala 18:52:@27263.4]
  assign _T_330 = $signed(b306_number); // @[Math.scala 406:49:@27271.4]
  assign _T_332 = $signed(_T_330) & $signed(32'shffff); // @[Math.scala 406:56:@27273.4]
  assign _T_333 = $signed(_T_332); // @[Math.scala 406:56:@27274.4]
  assign x474_sum_number = x474_sum_1_io_result; // @[Math.scala 154:22:@27285.4 Math.scala 155:14:@27286.4]
  assign _T_341 = x474_sum_number[31]; // @[FixedPoint.scala 50:25:@27290.4]
  assign _T_345 = _T_341 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@27292.4]
  assign _T_346 = x474_sum_number[31:8]; // @[FixedPoint.scala 18:52:@27293.4]
  assign _T_355 = $signed(x474_sum_number); // @[Math.scala 406:49:@27301.4]
  assign _T_357 = $signed(_T_355) & $signed(32'shff); // @[Math.scala 406:56:@27303.4]
  assign _T_358 = $signed(_T_357); // @[Math.scala 406:56:@27304.4]
  assign x477_sum_number = x477_sum_1_io_result; // @[Math.scala 154:22:@27315.4 Math.scala 155:14:@27316.4]
  assign _T_366 = x477_sum_number[31]; // @[FixedPoint.scala 50:25:@27320.4]
  assign _T_370 = _T_366 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@27322.4]
  assign _T_371 = x477_sum_number[31:4]; // @[FixedPoint.scala 18:52:@27323.4]
  assign _T_380 = $signed(x477_sum_number); // @[Math.scala 406:49:@27331.4]
  assign _T_382 = $signed(_T_380) & $signed(32'shf); // @[Math.scala 406:56:@27333.4]
  assign _T_383 = $signed(_T_382); // @[Math.scala 406:56:@27334.4]
  assign x480_sum_number = x480_sum_1_io_result; // @[Math.scala 154:22:@27345.4 Math.scala 155:14:@27346.4]
  assign _T_391 = x480_sum_number[31]; // @[FixedPoint.scala 50:25:@27350.4]
  assign _T_395 = _T_391 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27352.4]
  assign _T_396 = x480_sum_number[31:2]; // @[FixedPoint.scala 18:52:@27353.4]
  assign _T_405 = $signed(x480_sum_number); // @[Math.scala 406:49:@27361.4]
  assign _T_407 = $signed(_T_405) & $signed(32'sh3); // @[Math.scala 406:56:@27363.4]
  assign _T_408 = $signed(_T_407); // @[Math.scala 406:56:@27364.4]
  assign x483_sum_number = x483_sum_1_io_result; // @[Math.scala 154:22:@27375.4 Math.scala 155:14:@27376.4]
  assign _T_416 = x483_sum_number[31]; // @[FixedPoint.scala 50:25:@27380.4]
  assign _T_420 = _T_416 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27382.4]
  assign _T_421 = x483_sum_number[31:2]; // @[FixedPoint.scala 18:52:@27383.4]
  assign _T_432 = $signed(x483_sum_number); // @[Math.scala 406:49:@27398.4]
  assign _T_434 = $signed(_T_432) & $signed(32'sh3); // @[Math.scala 406:56:@27400.4]
  assign _T_435 = $signed(_T_434); // @[Math.scala 406:56:@27401.4]
  assign _T_439 = $signed(RetimeWrapper_3_io_out); // @[package.scala 96:25:@27409.4]
  assign x486_sum_number = x486_sum_1_io_result; // @[Math.scala 154:22:@27421.4 Math.scala 155:14:@27422.4]
  assign _T_447 = x486_sum_number[31]; // @[FixedPoint.scala 50:25:@27426.4]
  assign _T_451 = _T_447 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27428.4]
  assign _T_452 = x486_sum_number[31:2]; // @[FixedPoint.scala 18:52:@27429.4]
  assign _T_461 = $signed(x486_sum_number); // @[Math.scala 406:49:@27437.4]
  assign _T_463 = $signed(_T_461) & $signed(32'sh3); // @[Math.scala 406:56:@27439.4]
  assign _T_464 = $signed(_T_463); // @[Math.scala 406:56:@27440.4]
  assign x489_sum_number = x489_sum_1_io_result; // @[Math.scala 154:22:@27451.4 Math.scala 155:14:@27452.4]
  assign _T_474 = $signed(x489_sum_number); // @[Math.scala 465:37:@27457.4]
  assign x564_x490_D1 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@27495.4 package.scala 96:25:@27496.4]
  assign x565_x489_sum_D1_number = RetimeWrapper_6_io_out; // @[package.scala 96:25:@27504.4 package.scala 96:25:@27505.4]
  assign x492_sub_number = x492_sub_1_io_result; // @[Math.scala 195:22:@27477.4 Math.scala 196:14:@27478.4]
  assign _T_506 = x562_x317_D2_number[31]; // @[FixedPoint.scala 50:25:@27512.4]
  assign _T_510 = _T_506 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27514.4]
  assign _T_511 = x562_x317_D2_number[31:2]; // @[FixedPoint.scala 18:52:@27515.4]
  assign x321_number = {_T_510,_T_511}; // @[Cat.scala 30:58:@27516.4]
  assign _GEN_0 = {{9'd0}, x321_number}; // @[Math.scala 450:32:@27521.4]
  assign _T_516 = _GEN_0 << 9; // @[Math.scala 450:32:@27521.4]
  assign _GEN_1 = {{7'd0}, x321_number}; // @[Math.scala 450:32:@27526.4]
  assign _T_520 = _GEN_1 << 7; // @[Math.scala 450:32:@27526.4]
  assign _T_553 = ~ io_sigsIn_break; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 179:149:@27615.4]
  assign _T_557 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@27623.4 package.scala 96:25:@27624.4]
  assign _T_559 = io_rr ? _T_557 : 1'h0; // @[implicits.scala 55:10:@27625.4]
  assign _T_560 = _T_553 & _T_559; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 179:166:@27626.4]
  assign _T_562 = _T_560 & _T_553; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 179:255:@27628.4]
  assign _T_563 = _T_562 & io_sigsIn_backpressure; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 179:274:@27629.4]
  assign x568_b307_D21 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@27585.4 package.scala 96:25:@27586.4]
  assign _T_564 = _T_563 & x568_b307_D21; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 179:300:@27630.4]
  assign x567_b308_D21 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@27576.4 package.scala 96:25:@27577.4]
  assign x572_b305_D23_number = RetimeWrapper_14_io_out; // @[package.scala 96:25:@27644.4 package.scala 96:25:@27645.4]
  assign _T_578 = $signed(x572_b305_D23_number); // @[Math.scala 406:49:@27653.4]
  assign _T_580 = $signed(_T_578) & $signed(32'sh3); // @[Math.scala 406:56:@27655.4]
  assign _T_581 = $signed(_T_580); // @[Math.scala 406:56:@27656.4]
  assign _T_585 = $signed(RetimeWrapper_15_io_out); // @[package.scala 96:25:@27664.4]
  assign x497_number = $unsigned(_T_585); // @[implicits.scala 133:21:@27666.4]
  assign x573_b306_D23_number = RetimeWrapper_17_io_out; // @[package.scala 96:25:@27689.4 package.scala 96:25:@27690.4]
  assign _T_605 = $signed(x573_b306_D23_number); // @[Math.scala 465:37:@27695.4]
  assign x328 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@27680.4 package.scala 96:25:@27681.4]
  assign x329 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@27703.4 package.scala 96:25:@27704.4]
  assign x330 = x328 | x329; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 194:24:@27707.4]
  assign _T_621 = $signed(x497_number); // @[Math.scala 406:49:@27716.4]
  assign _T_623 = $signed(_T_621) & $signed(32'sh3); // @[Math.scala 406:56:@27718.4]
  assign _T_624 = $signed(_T_623); // @[Math.scala 406:56:@27719.4]
  assign _T_629 = x497_number[31]; // @[FixedPoint.scala 50:25:@27725.4]
  assign _T_633 = _T_629 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@27727.4]
  assign _T_634 = x497_number[31:2]; // @[FixedPoint.scala 18:52:@27728.4]
  assign x333_number = {_T_633,_T_634}; // @[Cat.scala 30:58:@27729.4]
  assign _GEN_2 = {{9'd0}, x333_number}; // @[Math.scala 450:32:@27734.4]
  assign _T_639 = _GEN_2 << 9; // @[Math.scala 450:32:@27734.4]
  assign _GEN_3 = {{7'd0}, x333_number}; // @[Math.scala 450:32:@27739.4]
  assign _T_643 = _GEN_3 << 7; // @[Math.scala 450:32:@27739.4]
  assign _T_685 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@27843.4 package.scala 96:25:@27844.4]
  assign _T_687 = io_rr ? _T_685 : 1'h0; // @[implicits.scala 55:10:@27845.4]
  assign _T_688 = _T_553 & _T_687; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 229:194:@27846.4]
  assign x581_x331_D21 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@27831.4 package.scala 96:25:@27832.4]
  assign _T_689 = _T_688 & x581_x331_D21; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 229:283:@27847.4]
  assign x577_b307_D45 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@27795.4 package.scala 96:25:@27796.4]
  assign _T_690 = _T_689 & x577_b307_D45; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 229:291:@27848.4]
  assign x576_b308_D45 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@27786.4 package.scala 96:25:@27787.4]
  assign x338_rdcol_number = x338_rdcol_1_io_result; // @[Math.scala 195:22:@27867.4 Math.scala 196:14:@27868.4]
  assign _T_705 = $signed(x338_rdcol_number); // @[Math.scala 465:37:@27873.4]
  assign x582_x328_D1 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@27890.4 package.scala 96:25:@27891.4]
  assign x339 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@27881.4 package.scala 96:25:@27882.4]
  assign x340 = x582_x328_D1 | x339; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 239:24:@27894.4]
  assign _T_720 = x338_rdcol_number[31]; // @[FixedPoint.scala 50:25:@27901.4]
  assign _T_724 = _T_720 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@27903.4]
  assign _T_725 = x338_rdcol_number[31:16]; // @[FixedPoint.scala 18:52:@27904.4]
  assign _T_738 = $signed(_T_705) & $signed(32'shffff); // @[Math.scala 406:56:@27921.4]
  assign _T_739 = $signed(_T_738); // @[Math.scala 406:56:@27922.4]
  assign _T_743 = $signed(RetimeWrapper_31_io_out); // @[package.scala 96:25:@27930.4]
  assign x504_sum_number = x504_sum_1_io_result; // @[Math.scala 154:22:@27942.4 Math.scala 155:14:@27943.4]
  assign _T_751 = x504_sum_number[31]; // @[FixedPoint.scala 50:25:@27947.4]
  assign _T_755 = _T_751 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@27949.4]
  assign _T_756 = x504_sum_number[31:8]; // @[FixedPoint.scala 18:52:@27950.4]
  assign _T_765 = $signed(x504_sum_number); // @[Math.scala 406:49:@27958.4]
  assign _T_767 = $signed(_T_765) & $signed(32'shff); // @[Math.scala 406:56:@27960.4]
  assign _T_768 = $signed(_T_767); // @[Math.scala 406:56:@27961.4]
  assign x507_sum_number = x507_sum_1_io_result; // @[Math.scala 154:22:@27972.4 Math.scala 155:14:@27973.4]
  assign _T_776 = x507_sum_number[31]; // @[FixedPoint.scala 50:25:@27977.4]
  assign _T_780 = _T_776 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@27979.4]
  assign _T_781 = x507_sum_number[31:4]; // @[FixedPoint.scala 18:52:@27980.4]
  assign _T_790 = $signed(x507_sum_number); // @[Math.scala 406:49:@27988.4]
  assign _T_792 = $signed(_T_790) & $signed(32'shf); // @[Math.scala 406:56:@27990.4]
  assign _T_793 = $signed(_T_792); // @[Math.scala 406:56:@27991.4]
  assign x510_sum_number = x510_sum_1_io_result; // @[Math.scala 154:22:@28002.4 Math.scala 155:14:@28003.4]
  assign _T_801 = x510_sum_number[31]; // @[FixedPoint.scala 50:25:@28007.4]
  assign _T_805 = _T_801 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28009.4]
  assign _T_806 = x510_sum_number[31:2]; // @[FixedPoint.scala 18:52:@28010.4]
  assign _T_815 = $signed(x510_sum_number); // @[Math.scala 406:49:@28018.4]
  assign _T_817 = $signed(_T_815) & $signed(32'sh3); // @[Math.scala 406:56:@28020.4]
  assign _T_818 = $signed(_T_817); // @[Math.scala 406:56:@28021.4]
  assign x513_sum_number = x513_sum_1_io_result; // @[Math.scala 154:22:@28032.4 Math.scala 155:14:@28033.4]
  assign _T_826 = x513_sum_number[31]; // @[FixedPoint.scala 50:25:@28037.4]
  assign _T_830 = _T_826 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28039.4]
  assign _T_831 = x513_sum_number[31:2]; // @[FixedPoint.scala 18:52:@28040.4]
  assign _T_840 = $signed(x513_sum_number); // @[Math.scala 406:49:@28048.4]
  assign _T_842 = $signed(_T_840) & $signed(32'sh3); // @[Math.scala 406:56:@28050.4]
  assign _T_843 = $signed(_T_842); // @[Math.scala 406:56:@28051.4]
  assign x516_sum_number = x516_sum_1_io_result; // @[Math.scala 154:22:@28062.4 Math.scala 155:14:@28063.4]
  assign _T_851 = x516_sum_number[31]; // @[FixedPoint.scala 50:25:@28067.4]
  assign _T_855 = _T_851 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28069.4]
  assign _T_856 = x516_sum_number[31:2]; // @[FixedPoint.scala 18:52:@28070.4]
  assign _T_867 = $signed(x516_sum_number); // @[Math.scala 406:49:@28085.4]
  assign _T_869 = $signed(_T_867) & $signed(32'sh3); // @[Math.scala 406:56:@28087.4]
  assign _T_870 = $signed(_T_869); // @[Math.scala 406:56:@28088.4]
  assign _T_874 = $signed(RetimeWrapper_33_io_out); // @[package.scala 96:25:@28096.4]
  assign x519_sum_number = x519_sum_1_io_result; // @[Math.scala 154:22:@28108.4 Math.scala 155:14:@28109.4]
  assign _T_886 = $signed(x519_sum_number); // @[Math.scala 465:37:@28116.4]
  assign x584_x520_D1 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@28154.4 package.scala 96:25:@28155.4]
  assign x585_x519_sum_D1_number = RetimeWrapper_36_io_out; // @[package.scala 96:25:@28163.4 package.scala 96:25:@28164.4]
  assign x522_sub_number = x522_sub_1_io_result; // @[Math.scala 195:22:@28136.4 Math.scala 196:14:@28137.4]
  assign _T_945 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@28227.4 package.scala 96:25:@28228.4]
  assign _T_947 = io_rr ? _T_945 : 1'h0; // @[implicits.scala 55:10:@28229.4]
  assign _T_948 = _T_553 & _T_947; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 314:194:@28230.4]
  assign x588_x341_D20 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@28215.4 package.scala 96:25:@28216.4]
  assign _T_949 = _T_948 & x588_x341_D20; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 314:283:@28231.4]
  assign _T_950 = _T_949 & x577_b307_D45; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 314:291:@28232.4]
  assign x347_rdcol_number = x347_rdcol_1_io_result; // @[Math.scala 195:22:@28251.4 Math.scala 196:14:@28252.4]
  assign _T_965 = $signed(x347_rdcol_number); // @[Math.scala 465:37:@28257.4]
  assign x348 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@28265.4 package.scala 96:25:@28266.4]
  assign x349 = x582_x328_D1 | x348; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 322:59:@28269.4]
  assign _T_977 = x347_rdcol_number[31]; // @[FixedPoint.scala 50:25:@28276.4]
  assign _T_981 = _T_977 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12:@28278.4]
  assign _T_982 = x347_rdcol_number[31:16]; // @[FixedPoint.scala 18:52:@28279.4]
  assign _T_995 = $signed(_T_965) & $signed(32'shffff); // @[Math.scala 406:56:@28296.4]
  assign _T_996 = $signed(_T_995); // @[Math.scala 406:56:@28297.4]
  assign _T_1000 = $signed(RetimeWrapper_43_io_out); // @[package.scala 96:25:@28305.4]
  assign x526_sum_number = x526_sum_1_io_result; // @[Math.scala 154:22:@28317.4 Math.scala 155:14:@28318.4]
  assign _T_1008 = x526_sum_number[31]; // @[FixedPoint.scala 50:25:@28322.4]
  assign _T_1012 = _T_1008 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:@28324.4]
  assign _T_1013 = x526_sum_number[31:8]; // @[FixedPoint.scala 18:52:@28325.4]
  assign _T_1022 = $signed(x526_sum_number); // @[Math.scala 406:49:@28333.4]
  assign _T_1024 = $signed(_T_1022) & $signed(32'shff); // @[Math.scala 406:56:@28335.4]
  assign _T_1025 = $signed(_T_1024); // @[Math.scala 406:56:@28336.4]
  assign x529_sum_number = x529_sum_1_io_result; // @[Math.scala 154:22:@28347.4 Math.scala 155:14:@28348.4]
  assign _T_1033 = x529_sum_number[31]; // @[FixedPoint.scala 50:25:@28352.4]
  assign _T_1037 = _T_1033 ? 4'hf : 4'h0; // @[Bitwise.scala 72:12:@28354.4]
  assign _T_1038 = x529_sum_number[31:4]; // @[FixedPoint.scala 18:52:@28355.4]
  assign _T_1047 = $signed(x529_sum_number); // @[Math.scala 406:49:@28363.4]
  assign _T_1049 = $signed(_T_1047) & $signed(32'shf); // @[Math.scala 406:56:@28365.4]
  assign _T_1050 = $signed(_T_1049); // @[Math.scala 406:56:@28366.4]
  assign x532_sum_number = x532_sum_1_io_result; // @[Math.scala 154:22:@28377.4 Math.scala 155:14:@28378.4]
  assign _T_1058 = x532_sum_number[31]; // @[FixedPoint.scala 50:25:@28382.4]
  assign _T_1062 = _T_1058 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28384.4]
  assign _T_1063 = x532_sum_number[31:2]; // @[FixedPoint.scala 18:52:@28385.4]
  assign _T_1072 = $signed(x532_sum_number); // @[Math.scala 406:49:@28393.4]
  assign _T_1074 = $signed(_T_1072) & $signed(32'sh3); // @[Math.scala 406:56:@28395.4]
  assign _T_1075 = $signed(_T_1074); // @[Math.scala 406:56:@28396.4]
  assign x535_sum_number = x535_sum_1_io_result; // @[Math.scala 154:22:@28407.4 Math.scala 155:14:@28408.4]
  assign _T_1083 = x535_sum_number[31]; // @[FixedPoint.scala 50:25:@28412.4]
  assign _T_1087 = _T_1083 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28414.4]
  assign _T_1088 = x535_sum_number[31:2]; // @[FixedPoint.scala 18:52:@28415.4]
  assign _T_1097 = $signed(x535_sum_number); // @[Math.scala 406:49:@28423.4]
  assign _T_1099 = $signed(_T_1097) & $signed(32'sh3); // @[Math.scala 406:56:@28425.4]
  assign _T_1100 = $signed(_T_1099); // @[Math.scala 406:56:@28426.4]
  assign x538_sum_number = x538_sum_1_io_result; // @[Math.scala 154:22:@28437.4 Math.scala 155:14:@28438.4]
  assign _T_1108 = x538_sum_number[31]; // @[FixedPoint.scala 50:25:@28442.4]
  assign _T_1112 = _T_1108 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28444.4]
  assign _T_1113 = x538_sum_number[31:2]; // @[FixedPoint.scala 18:52:@28445.4]
  assign _T_1124 = $signed(x538_sum_number); // @[Math.scala 406:49:@28460.4]
  assign _T_1126 = $signed(_T_1124) & $signed(32'sh3); // @[Math.scala 406:56:@28462.4]
  assign _T_1127 = $signed(_T_1126); // @[Math.scala 406:56:@28463.4]
  assign _T_1131 = $signed(RetimeWrapper_45_io_out); // @[package.scala 96:25:@28471.4]
  assign x541_sum_number = x541_sum_1_io_result; // @[Math.scala 154:22:@28483.4 Math.scala 155:14:@28484.4]
  assign _T_1141 = $signed(x541_sum_number); // @[Math.scala 465:37:@28489.4]
  assign x591_x542_D1 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@28536.4 package.scala 96:25:@28537.4]
  assign x590_x541_sum_D1_number = RetimeWrapper_47_io_out; // @[package.scala 96:25:@28527.4 package.scala 96:25:@28528.4]
  assign x544_sub_number = x544_sub_1_io_result; // @[Math.scala 195:22:@28509.4 Math.scala 196:14:@28510.4]
  assign _T_1197 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@28591.4 package.scala 96:25:@28592.4]
  assign _T_1199 = io_rr ? _T_1197 : 1'h0; // @[implicits.scala 55:10:@28593.4]
  assign _T_1200 = _T_553 & _T_1199; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 387:194:@28594.4]
  assign x593_x350_D20 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@28579.4 package.scala 96:25:@28580.4]
  assign _T_1201 = _T_1200 & x593_x350_D20; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 387:283:@28595.4]
  assign _T_1202 = _T_1201 & x577_b307_D45; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 387:291:@28596.4]
  assign x356_rdrow_number = x356_rdrow_1_io_result; // @[Math.scala 195:22:@28617.4 Math.scala 196:14:@28618.4]
  assign _T_1221 = $signed(x356_rdrow_number); // @[Math.scala 406:49:@28624.4]
  assign _T_1223 = $signed(_T_1221) & $signed(32'sh3); // @[Math.scala 406:56:@28626.4]
  assign _T_1224 = $signed(_T_1223); // @[Math.scala 406:56:@28627.4]
  assign _T_1228 = $signed(RetimeWrapper_52_io_out); // @[package.scala 96:25:@28635.4]
  assign x546_number = $unsigned(_T_1228); // @[implicits.scala 133:21:@28637.4]
  assign x358 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@28651.4 package.scala 96:25:@28652.4]
  assign x594_x329_D1 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@28660.4 package.scala 96:25:@28661.4]
  assign x359 = x358 | x594_x329_D1; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 407:24:@28664.4]
  assign _T_1254 = $signed(x546_number); // @[Math.scala 406:49:@28673.4]
  assign _T_1256 = $signed(_T_1254) & $signed(32'sh3); // @[Math.scala 406:56:@28675.4]
  assign _T_1257 = $signed(_T_1256); // @[Math.scala 406:56:@28676.4]
  assign _T_1262 = x546_number[31]; // @[FixedPoint.scala 50:25:@28682.4]
  assign _T_1266 = _T_1262 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28684.4]
  assign _T_1267 = x546_number[31:2]; // @[FixedPoint.scala 18:52:@28685.4]
  assign x362_number = {_T_1266,_T_1267}; // @[Cat.scala 30:58:@28686.4]
  assign _GEN_4 = {{9'd0}, x362_number}; // @[Math.scala 450:32:@28691.4]
  assign _T_1272 = _GEN_4 << 9; // @[Math.scala 450:32:@28691.4]
  assign _GEN_5 = {{7'd0}, x362_number}; // @[Math.scala 450:32:@28696.4]
  assign _T_1276 = _GEN_5 << 7; // @[Math.scala 450:32:@28696.4]
  assign _T_1306 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@28764.4 package.scala 96:25:@28765.4]
  assign _T_1308 = io_rr ? _T_1306 : 1'h0; // @[implicits.scala 55:10:@28766.4]
  assign _T_1309 = _T_553 & _T_1308; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 434:194:@28767.4]
  assign x597_x360_D20 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@28743.4 package.scala 96:25:@28744.4]
  assign _T_1310 = _T_1309 & x597_x360_D20; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 434:283:@28768.4]
  assign _T_1311 = _T_1310 & x577_b307_D45; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 434:291:@28769.4]
  assign x367 = x358 | x339; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 438:24:@28780.4]
  assign _T_1338 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@28822.4 package.scala 96:25:@28823.4]
  assign _T_1340 = io_rr ? _T_1338 : 1'h0; // @[implicits.scala 55:10:@28824.4]
  assign _T_1341 = _T_553 & _T_1340; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 451:194:@28825.4]
  assign x600_x368_D20 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@28810.4 package.scala 96:25:@28811.4]
  assign _T_1342 = _T_1341 & x600_x368_D20; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 451:283:@28826.4]
  assign _T_1343 = _T_1342 & x577_b307_D45; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 451:291:@28827.4]
  assign x372 = x358 | x348; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 455:24:@28838.4]
  assign _T_1367 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@28871.4 package.scala 96:25:@28872.4]
  assign _T_1369 = io_rr ? _T_1367 : 1'h0; // @[implicits.scala 55:10:@28873.4]
  assign _T_1370 = _T_553 & _T_1369; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 466:194:@28874.4]
  assign x601_x373_D20 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@28859.4 package.scala 96:25:@28860.4]
  assign _T_1371 = _T_1370 & x601_x373_D20; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 466:283:@28875.4]
  assign _T_1372 = _T_1371 & x577_b307_D45; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 466:291:@28876.4]
  assign x377_rdrow_number = x377_rdrow_1_io_result; // @[Math.scala 195:22:@28895.4 Math.scala 196:14:@28896.4]
  assign _T_1389 = $signed(x377_rdrow_number); // @[Math.scala 406:49:@28902.4]
  assign _T_1391 = $signed(_T_1389) & $signed(32'sh3); // @[Math.scala 406:56:@28904.4]
  assign _T_1392 = $signed(_T_1391); // @[Math.scala 406:56:@28905.4]
  assign _T_1396 = $signed(RetimeWrapper_65_io_out); // @[package.scala 96:25:@28913.4]
  assign x551_number = $unsigned(_T_1396); // @[implicits.scala 133:21:@28915.4]
  assign x379 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@28929.4 package.scala 96:25:@28930.4]
  assign x380 = x379 | x594_x329_D1; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 476:24:@28933.4]
  assign _T_1419 = $signed(x551_number); // @[Math.scala 406:49:@28942.4]
  assign _T_1421 = $signed(_T_1419) & $signed(32'sh3); // @[Math.scala 406:56:@28944.4]
  assign _T_1422 = $signed(_T_1421); // @[Math.scala 406:56:@28945.4]
  assign _T_1427 = x551_number[31]; // @[FixedPoint.scala 50:25:@28951.4]
  assign _T_1431 = _T_1427 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@28953.4]
  assign _T_1432 = x551_number[31:2]; // @[FixedPoint.scala 18:52:@28954.4]
  assign x383_number = {_T_1431,_T_1432}; // @[Cat.scala 30:58:@28955.4]
  assign _GEN_6 = {{9'd0}, x383_number}; // @[Math.scala 450:32:@28960.4]
  assign _T_1437 = _GEN_6 << 9; // @[Math.scala 450:32:@28960.4]
  assign _GEN_7 = {{7'd0}, x383_number}; // @[Math.scala 450:32:@28965.4]
  assign _T_1441 = _GEN_7 << 7; // @[Math.scala 450:32:@28965.4]
  assign _T_1471 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@29033.4 package.scala 96:25:@29034.4]
  assign _T_1473 = io_rr ? _T_1471 : 1'h0; // @[implicits.scala 55:10:@29035.4]
  assign _T_1474 = _T_553 & _T_1473; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 503:194:@29036.4]
  assign x604_x381_D20 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@29012.4 package.scala 96:25:@29013.4]
  assign _T_1475 = _T_1474 & x604_x381_D20; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 503:283:@29037.4]
  assign _T_1476 = _T_1475 & x577_b307_D45; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 503:291:@29038.4]
  assign x388 = x379 | x339; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 507:24:@29049.4]
  assign _T_1505 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@29093.4 package.scala 96:25:@29094.4]
  assign _T_1507 = io_rr ? _T_1505 : 1'h0; // @[implicits.scala 55:10:@29095.4]
  assign _T_1508 = _T_553 & _T_1507; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 528:194:@29096.4]
  assign x607_x389_D20 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@29081.4 package.scala 96:25:@29082.4]
  assign _T_1509 = _T_1508 & x607_x389_D20; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 528:283:@29097.4]
  assign _T_1510 = _T_1509 & x577_b307_D45; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 528:291:@29098.4]
  assign x393 = x379 | x348; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 532:59:@29109.4]
  assign _T_1534 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@29142.4 package.scala 96:25:@29143.4]
  assign _T_1536 = io_rr ? _T_1534 : 1'h0; // @[implicits.scala 55:10:@29144.4]
  assign _T_1537 = _T_553 & _T_1536; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 543:194:@29145.4]
  assign x608_x394_D20 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@29130.4 package.scala 96:25:@29131.4]
  assign _T_1538 = _T_1537 & x608_x394_D20; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 543:283:@29146.4]
  assign _T_1539 = _T_1538 & x577_b307_D45; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 543:291:@29147.4]
  assign x345_rd_0_number = x311_lb_0_io_rPort_4_output_0; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 310:29:@28218.4 sm_x416_inr_Foreach_SAMPLER_BOX.scala 314:408:@28239.4]
  assign _GEN_8 = {{1'd0}, x345_rd_0_number}; // @[Math.scala 450:32:@29159.4]
  assign x365_rd_0_number = x311_lb_0_io_rPort_0_output_0; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 430:29:@28755.4 sm_x416_inr_Foreach_SAMPLER_BOX.scala 434:408:@28776.4]
  assign _GEN_9 = {{1'd0}, x365_rd_0_number}; // @[Math.scala 450:32:@29171.4]
  assign x370_rd_0_number = x311_lb_0_io_rPort_5_output_0; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 447:29:@28813.4 sm_x416_inr_Foreach_SAMPLER_BOX.scala 451:408:@28834.4]
  assign _GEN_10 = {{2'd0}, x370_rd_0_number}; // @[Math.scala 450:32:@29183.4]
  assign x375_rd_0_number = x311_lb_0_io_rPort_2_output_0; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 462:29:@28862.4 sm_x416_inr_Foreach_SAMPLER_BOX.scala 466:408:@28883.4]
  assign _GEN_11 = {{1'd0}, x375_rd_0_number}; // @[Math.scala 450:32:@29195.4]
  assign x391_rd_0_number = x311_lb_0_io_rPort_3_output_0; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 524:29:@29084.4 sm_x416_inr_Foreach_SAMPLER_BOX.scala 528:408:@29105.4]
  assign _GEN_12 = {{1'd0}, x391_rd_0_number}; // @[Math.scala 450:32:@29207.4]
  assign x410_sum_number = x410_sum_1_io_result; // @[Math.scala 154:22:@29330.4 Math.scala 155:14:@29331.4]
  assign _T_1616 = x410_sum_number[7:4]; // @[FixedPoint.scala 18:52:@29336.4]
  assign _T_1637 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@29377.4 package.scala 96:25:@29378.4]
  assign _T_1639 = io_rr ? _T_1637 : 1'h0; // @[implicits.scala 55:10:@29379.4]
  assign x613_b307_D52 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@29359.4 package.scala 96:25:@29360.4]
  assign _T_1640 = _T_1639 & x613_b307_D52; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 591:117:@29380.4]
  assign x614_b308_D52 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@29368.4 package.scala 96:25:@29369.4]
  assign _T_1641 = _T_1640 & x614_b308_D52; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 591:123:@29381.4]
  assign x324_sum_number = x324_sum_1_io_result; // @[Math.scala 154:22:@27567.4 Math.scala 155:14:@27568.4]
  assign x569_x493_D13_number = RetimeWrapper_10_io_out; // @[package.scala 96:25:@27594.4 package.scala 96:25:@27595.4]
  assign x570_x471_D19_number = RetimeWrapper_11_io_out; // @[package.scala 96:25:@27603.4 package.scala 96:25:@27604.4]
  assign x578_x493_D37_number = RetimeWrapper_23_io_out; // @[package.scala 96:25:@27804.4 package.scala 96:25:@27805.4]
  assign x579_x498_D21_number = RetimeWrapper_24_io_out; // @[package.scala 96:25:@27813.4 package.scala 96:25:@27814.4]
  assign x580_x335_sum_D1_number = RetimeWrapper_25_io_out; // @[package.scala 96:25:@27822.4 package.scala 96:25:@27823.4]
  assign x344_sum_number = x344_sum_1_io_result; // @[Math.scala 154:22:@28197.4 Math.scala 155:14:@28198.4]
  assign x587_x523_D12_number = RetimeWrapper_38_io_out; // @[package.scala 96:25:@28206.4 package.scala 96:25:@28207.4]
  assign x353_sum_number = x353_sum_1_io_result; // @[Math.scala 154:22:@28561.4 Math.scala 155:14:@28562.4]
  assign x592_x545_D12_number = RetimeWrapper_49_io_out; // @[package.scala 96:25:@28570.4 package.scala 96:25:@28571.4]
  assign x596_x547_D20_number = RetimeWrapper_56_io_out; // @[package.scala 96:25:@28734.4 package.scala 96:25:@28735.4]
  assign x598_x364_sum_D1_number = RetimeWrapper_58_io_out; // @[package.scala 96:25:@28752.4 package.scala 96:25:@28753.4]
  assign x369_sum_number = x369_sum_1_io_result; // @[Math.scala 154:22:@28801.4 Math.scala 155:14:@28802.4]
  assign x374_sum_number = x374_sum_1_io_result; // @[Math.scala 154:22:@28850.4 Math.scala 155:14:@28851.4]
  assign x603_x385_sum_D1_number = RetimeWrapper_68_io_out; // @[package.scala 96:25:@29003.4 package.scala 96:25:@29004.4]
  assign x605_x552_D20_number = RetimeWrapper_70_io_out; // @[package.scala 96:25:@29021.4 package.scala 96:25:@29022.4]
  assign x390_sum_number = x390_sum_1_io_result; // @[Math.scala 154:22:@29072.4 Math.scala 155:14:@29073.4]
  assign x395_sum_number = x395_sum_1_io_result; // @[Math.scala 154:22:@29121.4 Math.scala 155:14:@29122.4]
  assign _T_1547 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@29165.4 package.scala 96:25:@29166.4]
  assign _T_1553 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@29177.4 package.scala 96:25:@29178.4]
  assign _T_1559 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@29189.4 package.scala 96:25:@29190.4]
  assign _T_1565 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@29201.4 package.scala 96:25:@29202.4]
  assign _T_1571 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@29213.4 package.scala 96:25:@29214.4]
  assign io_in_x279_TVALID = _T_1641 & io_sigsIn_backpressure; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 591:22:@29383.4]
  assign io_in_x279_TDATA = {{248'd0}, RetimeWrapper_86_io_out}; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 592:24:@29384.4]
  assign io_in_x278_TREADY = _T_211 & _T_213; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 67:22:@27097.4 sm_x416_inr_Foreach_SAMPLER_BOX.scala 69:22:@27105.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@27075.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 710:17:@27087.4]
  assign RetimeWrapper_clock = clock; // @[:@27108.4]
  assign RetimeWrapper_reset = reset; // @[:@27109.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27111.4]
  assign RetimeWrapper_io_in = io_in_x278_TDATA[7:0]; // @[package.scala 94:16:@27110.4]
  assign x311_lb_0_clock = clock; // @[:@27118.4]
  assign x311_lb_0_reset = reset; // @[:@27119.4]
  assign x311_lb_0_io_rPort_8_banks_1 = x592_x545_D12_number[1:0]; // @[MemInterfaceType.scala 106:58:@28599.4]
  assign x311_lb_0_io_rPort_8_banks_0 = x579_x498_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@28598.4]
  assign x311_lb_0_io_rPort_8_ofs_0 = x353_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@28600.4]
  assign x311_lb_0_io_rPort_8_en_0 = _T_1202 & x576_b308_D45; // @[MemInterfaceType.scala 110:79:@28602.4]
  assign x311_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28601.4]
  assign x311_lb_0_io_rPort_7_banks_1 = x578_x493_D37_number[1:0]; // @[MemInterfaceType.scala 106:58:@29041.4]
  assign x311_lb_0_io_rPort_7_banks_0 = x605_x552_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@29040.4]
  assign x311_lb_0_io_rPort_7_ofs_0 = x603_x385_sum_D1_number[9:0]; // @[MemInterfaceType.scala 107:54:@29042.4]
  assign x311_lb_0_io_rPort_7_en_0 = _T_1476 & x576_b308_D45; // @[MemInterfaceType.scala 110:79:@29044.4]
  assign x311_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@29043.4]
  assign x311_lb_0_io_rPort_6_banks_1 = x578_x493_D37_number[1:0]; // @[MemInterfaceType.scala 106:58:@27851.4]
  assign x311_lb_0_io_rPort_6_banks_0 = x579_x498_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@27850.4]
  assign x311_lb_0_io_rPort_6_ofs_0 = x580_x335_sum_D1_number[9:0]; // @[MemInterfaceType.scala 107:54:@27852.4]
  assign x311_lb_0_io_rPort_6_en_0 = _T_690 & x576_b308_D45; // @[MemInterfaceType.scala 110:79:@27854.4]
  assign x311_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@27853.4]
  assign x311_lb_0_io_rPort_5_banks_1 = x587_x523_D12_number[1:0]; // @[MemInterfaceType.scala 106:58:@28830.4]
  assign x311_lb_0_io_rPort_5_banks_0 = x596_x547_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@28829.4]
  assign x311_lb_0_io_rPort_5_ofs_0 = x369_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@28831.4]
  assign x311_lb_0_io_rPort_5_en_0 = _T_1343 & x576_b308_D45; // @[MemInterfaceType.scala 110:79:@28833.4]
  assign x311_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28832.4]
  assign x311_lb_0_io_rPort_4_banks_1 = x587_x523_D12_number[1:0]; // @[MemInterfaceType.scala 106:58:@28235.4]
  assign x311_lb_0_io_rPort_4_banks_0 = x579_x498_D21_number[2:0]; // @[MemInterfaceType.scala 106:58:@28234.4]
  assign x311_lb_0_io_rPort_4_ofs_0 = x344_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@28236.4]
  assign x311_lb_0_io_rPort_4_en_0 = _T_950 & x576_b308_D45; // @[MemInterfaceType.scala 110:79:@28238.4]
  assign x311_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28237.4]
  assign x311_lb_0_io_rPort_3_banks_1 = x587_x523_D12_number[1:0]; // @[MemInterfaceType.scala 106:58:@29101.4]
  assign x311_lb_0_io_rPort_3_banks_0 = x605_x552_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@29100.4]
  assign x311_lb_0_io_rPort_3_ofs_0 = x390_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@29102.4]
  assign x311_lb_0_io_rPort_3_en_0 = _T_1510 & x576_b308_D45; // @[MemInterfaceType.scala 110:79:@29104.4]
  assign x311_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@29103.4]
  assign x311_lb_0_io_rPort_2_banks_1 = x592_x545_D12_number[1:0]; // @[MemInterfaceType.scala 106:58:@28879.4]
  assign x311_lb_0_io_rPort_2_banks_0 = x596_x547_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@28878.4]
  assign x311_lb_0_io_rPort_2_ofs_0 = x374_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@28880.4]
  assign x311_lb_0_io_rPort_2_en_0 = _T_1372 & x576_b308_D45; // @[MemInterfaceType.scala 110:79:@28882.4]
  assign x311_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28881.4]
  assign x311_lb_0_io_rPort_1_banks_1 = x592_x545_D12_number[1:0]; // @[MemInterfaceType.scala 106:58:@29150.4]
  assign x311_lb_0_io_rPort_1_banks_0 = x605_x552_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@29149.4]
  assign x311_lb_0_io_rPort_1_ofs_0 = x395_sum_number[9:0]; // @[MemInterfaceType.scala 107:54:@29151.4]
  assign x311_lb_0_io_rPort_1_en_0 = _T_1539 & x576_b308_D45; // @[MemInterfaceType.scala 110:79:@29153.4]
  assign x311_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@29152.4]
  assign x311_lb_0_io_rPort_0_banks_1 = x578_x493_D37_number[1:0]; // @[MemInterfaceType.scala 106:58:@28772.4]
  assign x311_lb_0_io_rPort_0_banks_0 = x596_x547_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@28771.4]
  assign x311_lb_0_io_rPort_0_ofs_0 = x598_x364_sum_D1_number[9:0]; // @[MemInterfaceType.scala 107:54:@28773.4]
  assign x311_lb_0_io_rPort_0_en_0 = _T_1311 & x576_b308_D45; // @[MemInterfaceType.scala 110:79:@28775.4]
  assign x311_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@28774.4]
  assign x311_lb_0_io_wPort_0_banks_1 = x569_x493_D13_number[1:0]; // @[MemInterfaceType.scala 88:58:@27633.4]
  assign x311_lb_0_io_wPort_0_banks_0 = x570_x471_D19_number[2:0]; // @[MemInterfaceType.scala 88:58:@27632.4]
  assign x311_lb_0_io_wPort_0_ofs_0 = x324_sum_number[9:0]; // @[MemInterfaceType.scala 89:54:@27634.4]
  assign x311_lb_0_io_wPort_0_data_0 = RetimeWrapper_12_io_out; // @[MemInterfaceType.scala 90:56:@27635.4]
  assign x311_lb_0_io_wPort_0_en_0 = _T_564 & x567_b308_D21; // @[MemInterfaceType.scala 93:57:@27637.4]
  assign RetimeWrapper_1_clock = clock; // @[:@27240.4]
  assign RetimeWrapper_1_reset = reset; // @[:@27241.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27243.4]
  assign RetimeWrapper_1_io_in = _T_293 | _T_291; // @[package.scala 94:16:@27242.4]
  assign x474_sum_1_clock = clock; // @[:@27280.4]
  assign x474_sum_1_reset = reset; // @[:@27281.4]
  assign x474_sum_1_io_a = {_T_320,_T_321}; // @[Math.scala 151:17:@27282.4]
  assign x474_sum_1_io_b = $unsigned(_T_333); // @[Math.scala 152:17:@27283.4]
  assign x474_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@27284.4]
  assign x477_sum_1_clock = clock; // @[:@27310.4]
  assign x477_sum_1_reset = reset; // @[:@27311.4]
  assign x477_sum_1_io_a = {_T_345,_T_346}; // @[Math.scala 151:17:@27312.4]
  assign x477_sum_1_io_b = $unsigned(_T_358); // @[Math.scala 152:17:@27313.4]
  assign x477_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@27314.4]
  assign x480_sum_1_clock = clock; // @[:@27340.4]
  assign x480_sum_1_reset = reset; // @[:@27341.4]
  assign x480_sum_1_io_a = {_T_370,_T_371}; // @[Math.scala 151:17:@27342.4]
  assign x480_sum_1_io_b = $unsigned(_T_383); // @[Math.scala 152:17:@27343.4]
  assign x480_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@27344.4]
  assign x483_sum_1_clock = clock; // @[:@27370.4]
  assign x483_sum_1_reset = reset; // @[:@27371.4]
  assign x483_sum_1_io_a = {_T_395,_T_396}; // @[Math.scala 151:17:@27372.4]
  assign x483_sum_1_io_b = $unsigned(_T_408); // @[Math.scala 152:17:@27373.4]
  assign x483_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@27374.4]
  assign RetimeWrapper_2_clock = clock; // @[:@27386.4]
  assign RetimeWrapper_2_reset = reset; // @[:@27387.4]
  assign RetimeWrapper_2_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@27389.4]
  assign RetimeWrapper_2_io_in = {_T_420,_T_421}; // @[package.scala 94:16:@27388.4]
  assign RetimeWrapper_3_clock = clock; // @[:@27403.4]
  assign RetimeWrapper_3_reset = reset; // @[:@27404.4]
  assign RetimeWrapper_3_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@27407.4]
  assign RetimeWrapper_3_io_in = $unsigned(_T_435); // @[package.scala 94:16:@27406.4]
  assign x486_sum_1_clock = clock; // @[:@27416.4]
  assign x486_sum_1_reset = reset; // @[:@27417.4]
  assign x486_sum_1_io_a = RetimeWrapper_2_io_out; // @[Math.scala 151:17:@27418.4]
  assign x486_sum_1_io_b = $unsigned(_T_439); // @[Math.scala 152:17:@27419.4]
  assign x486_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@27420.4]
  assign x489_sum_1_clock = clock; // @[:@27446.4]
  assign x489_sum_1_reset = reset; // @[:@27447.4]
  assign x489_sum_1_io_a = {_T_451,_T_452}; // @[Math.scala 151:17:@27448.4]
  assign x489_sum_1_io_b = $unsigned(_T_464); // @[Math.scala 152:17:@27449.4]
  assign x489_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@27450.4]
  assign x492_sub_1_clock = clock; // @[:@27472.4]
  assign x492_sub_1_reset = reset; // @[:@27473.4]
  assign x492_sub_1_io_a = x489_sum_1_io_result; // @[Math.scala 192:17:@27474.4]
  assign x492_sub_1_io_b = 32'h3; // @[Math.scala 193:17:@27475.4]
  assign x492_sub_1_io_flow = io_in_x279_TREADY; // @[Math.scala 194:20:@27476.4]
  assign RetimeWrapper_4_clock = clock; // @[:@27482.4]
  assign RetimeWrapper_4_reset = reset; // @[:@27483.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27485.4]
  assign RetimeWrapper_4_io_in = $signed(_T_474) < $signed(32'sh6); // @[package.scala 94:16:@27484.4]
  assign RetimeWrapper_5_clock = clock; // @[:@27491.4]
  assign RetimeWrapper_5_reset = reset; // @[:@27492.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27494.4]
  assign RetimeWrapper_5_io_in = $signed(_T_474) < $signed(32'sh3); // @[package.scala 94:16:@27493.4]
  assign RetimeWrapper_6_clock = clock; // @[:@27500.4]
  assign RetimeWrapper_6_reset = reset; // @[:@27501.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27503.4]
  assign RetimeWrapper_6_io_in = x489_sum_1_io_result; // @[package.scala 94:16:@27502.4]
  assign x496_sum_1_clock = clock; // @[:@27531.4]
  assign x496_sum_1_reset = reset; // @[:@27532.4]
  assign x496_sum_1_io_a = _T_516[31:0]; // @[Math.scala 151:17:@27533.4]
  assign x496_sum_1_io_b = _T_520[31:0]; // @[Math.scala 152:17:@27534.4]
  assign x496_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@27535.4]
  assign x323_div_1_clock = clock; // @[:@27543.4]
  assign x323_div_1_reset = reset; // @[:@27544.4]
  assign x323_div_1_io_a = __1_io_result; // @[Math.scala 328:17:@27545.4]
  assign x323_div_1_io_flow = io_in_x279_TREADY; // @[Math.scala 330:20:@27547.4]
  assign RetimeWrapper_7_clock = clock; // @[:@27553.4]
  assign RetimeWrapper_7_reset = reset; // @[:@27554.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27556.4]
  assign RetimeWrapper_7_io_in = x496_sum_1_io_result; // @[package.scala 94:16:@27555.4]
  assign x324_sum_1_clock = clock; // @[:@27562.4]
  assign x324_sum_1_reset = reset; // @[:@27563.4]
  assign x324_sum_1_io_a = RetimeWrapper_7_io_out; // @[Math.scala 151:17:@27564.4]
  assign x324_sum_1_io_b = x323_div_1_io_result; // @[Math.scala 152:17:@27565.4]
  assign x324_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@27566.4]
  assign RetimeWrapper_8_clock = clock; // @[:@27572.4]
  assign RetimeWrapper_8_reset = reset; // @[:@27573.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27575.4]
  assign RetimeWrapper_8_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@27574.4]
  assign RetimeWrapper_9_clock = clock; // @[:@27581.4]
  assign RetimeWrapper_9_reset = reset; // @[:@27582.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27584.4]
  assign RetimeWrapper_9_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@27583.4]
  assign RetimeWrapper_10_clock = clock; // @[:@27590.4]
  assign RetimeWrapper_10_reset = reset; // @[:@27591.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27593.4]
  assign RetimeWrapper_10_io_in = x564_x490_D1 ? x565_x489_sum_D1_number : x492_sub_number; // @[package.scala 94:16:@27592.4]
  assign RetimeWrapper_11_clock = clock; // @[:@27599.4]
  assign RetimeWrapper_11_reset = reset; // @[:@27600.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27602.4]
  assign RetimeWrapper_11_io_in = $unsigned(_T_311); // @[package.scala 94:16:@27601.4]
  assign RetimeWrapper_12_clock = clock; // @[:@27608.4]
  assign RetimeWrapper_12_reset = reset; // @[:@27609.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27611.4]
  assign RetimeWrapper_12_io_in = RetimeWrapper_io_out; // @[package.scala 94:16:@27610.4]
  assign RetimeWrapper_13_clock = clock; // @[:@27619.4]
  assign RetimeWrapper_13_reset = reset; // @[:@27620.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27622.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27621.4]
  assign RetimeWrapper_14_clock = clock; // @[:@27640.4]
  assign RetimeWrapper_14_reset = reset; // @[:@27641.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27643.4]
  assign RetimeWrapper_14_io_in = __io_result; // @[package.scala 94:16:@27642.4]
  assign RetimeWrapper_15_clock = clock; // @[:@27658.4]
  assign RetimeWrapper_15_reset = reset; // @[:@27659.4]
  assign RetimeWrapper_15_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@27662.4]
  assign RetimeWrapper_15_io_in = $unsigned(_T_581); // @[package.scala 94:16:@27661.4]
  assign RetimeWrapper_16_clock = clock; // @[:@27676.4]
  assign RetimeWrapper_16_reset = reset; // @[:@27677.4]
  assign RetimeWrapper_16_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@27679.4]
  assign RetimeWrapper_16_io_in = $signed(_T_578) < $signed(32'sh0); // @[package.scala 94:16:@27678.4]
  assign RetimeWrapper_17_clock = clock; // @[:@27685.4]
  assign RetimeWrapper_17_reset = reset; // @[:@27686.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27688.4]
  assign RetimeWrapper_17_io_in = __1_io_result; // @[package.scala 94:16:@27687.4]
  assign RetimeWrapper_18_clock = clock; // @[:@27699.4]
  assign RetimeWrapper_18_reset = reset; // @[:@27700.4]
  assign RetimeWrapper_18_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@27702.4]
  assign RetimeWrapper_18_io_in = $signed(_T_605) < $signed(32'sh0); // @[package.scala 94:16:@27701.4]
  assign x501_sum_1_clock = clock; // @[:@27744.4]
  assign x501_sum_1_reset = reset; // @[:@27745.4]
  assign x501_sum_1_io_a = _T_639[31:0]; // @[Math.scala 151:17:@27746.4]
  assign x501_sum_1_io_b = _T_643[31:0]; // @[Math.scala 152:17:@27747.4]
  assign x501_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@27748.4]
  assign RetimeWrapper_19_clock = clock; // @[:@27754.4]
  assign RetimeWrapper_19_reset = reset; // @[:@27755.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27757.4]
  assign RetimeWrapper_19_io_in = x501_sum_1_io_result; // @[package.scala 94:16:@27756.4]
  assign RetimeWrapper_20_clock = clock; // @[:@27763.4]
  assign RetimeWrapper_20_reset = reset; // @[:@27764.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27766.4]
  assign RetimeWrapper_20_io_in = x323_div_1_io_result; // @[package.scala 94:16:@27765.4]
  assign x335_sum_1_clock = clock; // @[:@27772.4]
  assign x335_sum_1_reset = reset; // @[:@27773.4]
  assign x335_sum_1_io_a = RetimeWrapper_19_io_out; // @[Math.scala 151:17:@27774.4]
  assign x335_sum_1_io_b = RetimeWrapper_20_io_out; // @[Math.scala 152:17:@27775.4]
  assign x335_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@27776.4]
  assign RetimeWrapper_21_clock = clock; // @[:@27782.4]
  assign RetimeWrapper_21_reset = reset; // @[:@27783.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27785.4]
  assign RetimeWrapper_21_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@27784.4]
  assign RetimeWrapper_22_clock = clock; // @[:@27791.4]
  assign RetimeWrapper_22_reset = reset; // @[:@27792.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27794.4]
  assign RetimeWrapper_22_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@27793.4]
  assign RetimeWrapper_23_clock = clock; // @[:@27800.4]
  assign RetimeWrapper_23_reset = reset; // @[:@27801.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27803.4]
  assign RetimeWrapper_23_io_in = x564_x490_D1 ? x565_x489_sum_D1_number : x492_sub_number; // @[package.scala 94:16:@27802.4]
  assign RetimeWrapper_24_clock = clock; // @[:@27809.4]
  assign RetimeWrapper_24_reset = reset; // @[:@27810.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27812.4]
  assign RetimeWrapper_24_io_in = $unsigned(_T_624); // @[package.scala 94:16:@27811.4]
  assign RetimeWrapper_25_clock = clock; // @[:@27818.4]
  assign RetimeWrapper_25_reset = reset; // @[:@27819.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27821.4]
  assign RetimeWrapper_25_io_in = x335_sum_1_io_result; // @[package.scala 94:16:@27820.4]
  assign RetimeWrapper_26_clock = clock; // @[:@27827.4]
  assign RetimeWrapper_26_reset = reset; // @[:@27828.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27830.4]
  assign RetimeWrapper_26_io_in = ~ x330; // @[package.scala 94:16:@27829.4]
  assign RetimeWrapper_27_clock = clock; // @[:@27839.4]
  assign RetimeWrapper_27_reset = reset; // @[:@27840.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27842.4]
  assign RetimeWrapper_27_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27841.4]
  assign x338_rdcol_1_clock = clock; // @[:@27862.4]
  assign x338_rdcol_1_reset = reset; // @[:@27863.4]
  assign x338_rdcol_1_io_a = RetimeWrapper_17_io_out; // @[Math.scala 192:17:@27864.4]
  assign x338_rdcol_1_io_b = 32'h1; // @[Math.scala 193:17:@27865.4]
  assign x338_rdcol_1_io_flow = io_in_x279_TREADY; // @[Math.scala 194:20:@27866.4]
  assign RetimeWrapper_28_clock = clock; // @[:@27877.4]
  assign RetimeWrapper_28_reset = reset; // @[:@27878.4]
  assign RetimeWrapper_28_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@27880.4]
  assign RetimeWrapper_28_io_in = $signed(_T_705) < $signed(32'sh0); // @[package.scala 94:16:@27879.4]
  assign RetimeWrapper_29_clock = clock; // @[:@27886.4]
  assign RetimeWrapper_29_reset = reset; // @[:@27887.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27889.4]
  assign RetimeWrapper_29_io_in = RetimeWrapper_16_io_out; // @[package.scala 94:16:@27888.4]
  assign RetimeWrapper_30_clock = clock; // @[:@27907.4]
  assign RetimeWrapper_30_reset = reset; // @[:@27908.4]
  assign RetimeWrapper_30_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@27910.4]
  assign RetimeWrapper_30_io_in = {_T_724,_T_725}; // @[package.scala 94:16:@27909.4]
  assign RetimeWrapper_31_clock = clock; // @[:@27924.4]
  assign RetimeWrapper_31_reset = reset; // @[:@27925.4]
  assign RetimeWrapper_31_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@27928.4]
  assign RetimeWrapper_31_io_in = $unsigned(_T_739); // @[package.scala 94:16:@27927.4]
  assign x504_sum_1_clock = clock; // @[:@27937.4]
  assign x504_sum_1_reset = reset; // @[:@27938.4]
  assign x504_sum_1_io_a = RetimeWrapper_30_io_out; // @[Math.scala 151:17:@27939.4]
  assign x504_sum_1_io_b = $unsigned(_T_743); // @[Math.scala 152:17:@27940.4]
  assign x504_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@27941.4]
  assign x507_sum_1_clock = clock; // @[:@27967.4]
  assign x507_sum_1_reset = reset; // @[:@27968.4]
  assign x507_sum_1_io_a = {_T_755,_T_756}; // @[Math.scala 151:17:@27969.4]
  assign x507_sum_1_io_b = $unsigned(_T_768); // @[Math.scala 152:17:@27970.4]
  assign x507_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@27971.4]
  assign x510_sum_1_clock = clock; // @[:@27997.4]
  assign x510_sum_1_reset = reset; // @[:@27998.4]
  assign x510_sum_1_io_a = {_T_780,_T_781}; // @[Math.scala 151:17:@27999.4]
  assign x510_sum_1_io_b = $unsigned(_T_793); // @[Math.scala 152:17:@28000.4]
  assign x510_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@28001.4]
  assign x513_sum_1_clock = clock; // @[:@28027.4]
  assign x513_sum_1_reset = reset; // @[:@28028.4]
  assign x513_sum_1_io_a = {_T_805,_T_806}; // @[Math.scala 151:17:@28029.4]
  assign x513_sum_1_io_b = $unsigned(_T_818); // @[Math.scala 152:17:@28030.4]
  assign x513_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@28031.4]
  assign x516_sum_1_clock = clock; // @[:@28057.4]
  assign x516_sum_1_reset = reset; // @[:@28058.4]
  assign x516_sum_1_io_a = {_T_830,_T_831}; // @[Math.scala 151:17:@28059.4]
  assign x516_sum_1_io_b = $unsigned(_T_843); // @[Math.scala 152:17:@28060.4]
  assign x516_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@28061.4]
  assign RetimeWrapper_32_clock = clock; // @[:@28073.4]
  assign RetimeWrapper_32_reset = reset; // @[:@28074.4]
  assign RetimeWrapper_32_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@28076.4]
  assign RetimeWrapper_32_io_in = {_T_855,_T_856}; // @[package.scala 94:16:@28075.4]
  assign RetimeWrapper_33_clock = clock; // @[:@28090.4]
  assign RetimeWrapper_33_reset = reset; // @[:@28091.4]
  assign RetimeWrapper_33_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@28094.4]
  assign RetimeWrapper_33_io_in = $unsigned(_T_870); // @[package.scala 94:16:@28093.4]
  assign x519_sum_1_clock = clock; // @[:@28103.4]
  assign x519_sum_1_reset = reset; // @[:@28104.4]
  assign x519_sum_1_io_a = RetimeWrapper_32_io_out; // @[Math.scala 151:17:@28105.4]
  assign x519_sum_1_io_b = $unsigned(_T_874); // @[Math.scala 152:17:@28106.4]
  assign x519_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@28107.4]
  assign x522_sub_1_clock = clock; // @[:@28131.4]
  assign x522_sub_1_reset = reset; // @[:@28132.4]
  assign x522_sub_1_io_a = x519_sum_1_io_result; // @[Math.scala 192:17:@28133.4]
  assign x522_sub_1_io_b = 32'h3; // @[Math.scala 193:17:@28134.4]
  assign x522_sub_1_io_flow = io_in_x279_TREADY; // @[Math.scala 194:20:@28135.4]
  assign RetimeWrapper_34_clock = clock; // @[:@28141.4]
  assign RetimeWrapper_34_reset = reset; // @[:@28142.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28144.4]
  assign RetimeWrapper_34_io_in = $signed(_T_886) < $signed(32'sh6); // @[package.scala 94:16:@28143.4]
  assign RetimeWrapper_35_clock = clock; // @[:@28150.4]
  assign RetimeWrapper_35_reset = reset; // @[:@28151.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28153.4]
  assign RetimeWrapper_35_io_in = $signed(_T_886) < $signed(32'sh3); // @[package.scala 94:16:@28152.4]
  assign RetimeWrapper_36_clock = clock; // @[:@28159.4]
  assign RetimeWrapper_36_reset = reset; // @[:@28160.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28162.4]
  assign RetimeWrapper_36_io_in = x519_sum_1_io_result; // @[package.scala 94:16:@28161.4]
  assign x343_div_1_clock = clock; // @[:@28173.4]
  assign x343_div_1_reset = reset; // @[:@28174.4]
  assign x343_div_1_io_a = x338_rdcol_1_io_result; // @[Math.scala 328:17:@28175.4]
  assign x343_div_1_io_flow = io_in_x279_TREADY; // @[Math.scala 330:20:@28177.4]
  assign RetimeWrapper_37_clock = clock; // @[:@28183.4]
  assign RetimeWrapper_37_reset = reset; // @[:@28184.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28186.4]
  assign RetimeWrapper_37_io_in = x501_sum_1_io_result; // @[package.scala 94:16:@28185.4]
  assign x344_sum_1_clock = clock; // @[:@28192.4]
  assign x344_sum_1_reset = reset; // @[:@28193.4]
  assign x344_sum_1_io_a = RetimeWrapper_37_io_out; // @[Math.scala 151:17:@28194.4]
  assign x344_sum_1_io_b = x343_div_1_io_result; // @[Math.scala 152:17:@28195.4]
  assign x344_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@28196.4]
  assign RetimeWrapper_38_clock = clock; // @[:@28202.4]
  assign RetimeWrapper_38_reset = reset; // @[:@28203.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28205.4]
  assign RetimeWrapper_38_io_in = x584_x520_D1 ? x585_x519_sum_D1_number : x522_sub_number; // @[package.scala 94:16:@28204.4]
  assign RetimeWrapper_39_clock = clock; // @[:@28211.4]
  assign RetimeWrapper_39_reset = reset; // @[:@28212.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28214.4]
  assign RetimeWrapper_39_io_in = ~ x340; // @[package.scala 94:16:@28213.4]
  assign RetimeWrapper_40_clock = clock; // @[:@28223.4]
  assign RetimeWrapper_40_reset = reset; // @[:@28224.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28226.4]
  assign RetimeWrapper_40_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28225.4]
  assign x347_rdcol_1_clock = clock; // @[:@28246.4]
  assign x347_rdcol_1_reset = reset; // @[:@28247.4]
  assign x347_rdcol_1_io_a = RetimeWrapper_17_io_out; // @[Math.scala 192:17:@28248.4]
  assign x347_rdcol_1_io_b = 32'h2; // @[Math.scala 193:17:@28249.4]
  assign x347_rdcol_1_io_flow = io_in_x279_TREADY; // @[Math.scala 194:20:@28250.4]
  assign RetimeWrapper_41_clock = clock; // @[:@28261.4]
  assign RetimeWrapper_41_reset = reset; // @[:@28262.4]
  assign RetimeWrapper_41_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@28264.4]
  assign RetimeWrapper_41_io_in = $signed(_T_965) < $signed(32'sh0); // @[package.scala 94:16:@28263.4]
  assign RetimeWrapper_42_clock = clock; // @[:@28282.4]
  assign RetimeWrapper_42_reset = reset; // @[:@28283.4]
  assign RetimeWrapper_42_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@28285.4]
  assign RetimeWrapper_42_io_in = {_T_981,_T_982}; // @[package.scala 94:16:@28284.4]
  assign RetimeWrapper_43_clock = clock; // @[:@28299.4]
  assign RetimeWrapper_43_reset = reset; // @[:@28300.4]
  assign RetimeWrapper_43_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@28303.4]
  assign RetimeWrapper_43_io_in = $unsigned(_T_996); // @[package.scala 94:16:@28302.4]
  assign x526_sum_1_clock = clock; // @[:@28312.4]
  assign x526_sum_1_reset = reset; // @[:@28313.4]
  assign x526_sum_1_io_a = RetimeWrapper_42_io_out; // @[Math.scala 151:17:@28314.4]
  assign x526_sum_1_io_b = $unsigned(_T_1000); // @[Math.scala 152:17:@28315.4]
  assign x526_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@28316.4]
  assign x529_sum_1_clock = clock; // @[:@28342.4]
  assign x529_sum_1_reset = reset; // @[:@28343.4]
  assign x529_sum_1_io_a = {_T_1012,_T_1013}; // @[Math.scala 151:17:@28344.4]
  assign x529_sum_1_io_b = $unsigned(_T_1025); // @[Math.scala 152:17:@28345.4]
  assign x529_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@28346.4]
  assign x532_sum_1_clock = clock; // @[:@28372.4]
  assign x532_sum_1_reset = reset; // @[:@28373.4]
  assign x532_sum_1_io_a = {_T_1037,_T_1038}; // @[Math.scala 151:17:@28374.4]
  assign x532_sum_1_io_b = $unsigned(_T_1050); // @[Math.scala 152:17:@28375.4]
  assign x532_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@28376.4]
  assign x535_sum_1_clock = clock; // @[:@28402.4]
  assign x535_sum_1_reset = reset; // @[:@28403.4]
  assign x535_sum_1_io_a = {_T_1062,_T_1063}; // @[Math.scala 151:17:@28404.4]
  assign x535_sum_1_io_b = $unsigned(_T_1075); // @[Math.scala 152:17:@28405.4]
  assign x535_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@28406.4]
  assign x538_sum_1_clock = clock; // @[:@28432.4]
  assign x538_sum_1_reset = reset; // @[:@28433.4]
  assign x538_sum_1_io_a = {_T_1087,_T_1088}; // @[Math.scala 151:17:@28434.4]
  assign x538_sum_1_io_b = $unsigned(_T_1100); // @[Math.scala 152:17:@28435.4]
  assign x538_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@28436.4]
  assign RetimeWrapper_44_clock = clock; // @[:@28448.4]
  assign RetimeWrapper_44_reset = reset; // @[:@28449.4]
  assign RetimeWrapper_44_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@28451.4]
  assign RetimeWrapper_44_io_in = {_T_1112,_T_1113}; // @[package.scala 94:16:@28450.4]
  assign RetimeWrapper_45_clock = clock; // @[:@28465.4]
  assign RetimeWrapper_45_reset = reset; // @[:@28466.4]
  assign RetimeWrapper_45_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@28469.4]
  assign RetimeWrapper_45_io_in = $unsigned(_T_1127); // @[package.scala 94:16:@28468.4]
  assign x541_sum_1_clock = clock; // @[:@28478.4]
  assign x541_sum_1_reset = reset; // @[:@28479.4]
  assign x541_sum_1_io_a = RetimeWrapper_44_io_out; // @[Math.scala 151:17:@28480.4]
  assign x541_sum_1_io_b = $unsigned(_T_1131); // @[Math.scala 152:17:@28481.4]
  assign x541_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@28482.4]
  assign x544_sub_1_clock = clock; // @[:@28504.4]
  assign x544_sub_1_reset = reset; // @[:@28505.4]
  assign x544_sub_1_io_a = x541_sum_1_io_result; // @[Math.scala 192:17:@28506.4]
  assign x544_sub_1_io_b = 32'h3; // @[Math.scala 193:17:@28507.4]
  assign x544_sub_1_io_flow = io_in_x279_TREADY; // @[Math.scala 194:20:@28508.4]
  assign RetimeWrapper_46_clock = clock; // @[:@28514.4]
  assign RetimeWrapper_46_reset = reset; // @[:@28515.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28517.4]
  assign RetimeWrapper_46_io_in = $signed(_T_1141) < $signed(32'sh6); // @[package.scala 94:16:@28516.4]
  assign RetimeWrapper_47_clock = clock; // @[:@28523.4]
  assign RetimeWrapper_47_reset = reset; // @[:@28524.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28526.4]
  assign RetimeWrapper_47_io_in = x541_sum_1_io_result; // @[package.scala 94:16:@28525.4]
  assign RetimeWrapper_48_clock = clock; // @[:@28532.4]
  assign RetimeWrapper_48_reset = reset; // @[:@28533.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28535.4]
  assign RetimeWrapper_48_io_in = $signed(_T_1141) < $signed(32'sh3); // @[package.scala 94:16:@28534.4]
  assign x352_div_1_clock = clock; // @[:@28546.4]
  assign x352_div_1_reset = reset; // @[:@28547.4]
  assign x352_div_1_io_a = x347_rdcol_1_io_result; // @[Math.scala 328:17:@28548.4]
  assign x352_div_1_io_flow = io_in_x279_TREADY; // @[Math.scala 330:20:@28550.4]
  assign x353_sum_1_clock = clock; // @[:@28556.4]
  assign x353_sum_1_reset = reset; // @[:@28557.4]
  assign x353_sum_1_io_a = RetimeWrapper_37_io_out; // @[Math.scala 151:17:@28558.4]
  assign x353_sum_1_io_b = x352_div_1_io_result; // @[Math.scala 152:17:@28559.4]
  assign x353_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@28560.4]
  assign RetimeWrapper_49_clock = clock; // @[:@28566.4]
  assign RetimeWrapper_49_reset = reset; // @[:@28567.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28569.4]
  assign RetimeWrapper_49_io_in = x591_x542_D1 ? x590_x541_sum_D1_number : x544_sub_number; // @[package.scala 94:16:@28568.4]
  assign RetimeWrapper_50_clock = clock; // @[:@28575.4]
  assign RetimeWrapper_50_reset = reset; // @[:@28576.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28578.4]
  assign RetimeWrapper_50_io_in = ~ x349; // @[package.scala 94:16:@28577.4]
  assign RetimeWrapper_51_clock = clock; // @[:@28587.4]
  assign RetimeWrapper_51_reset = reset; // @[:@28588.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28590.4]
  assign RetimeWrapper_51_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28589.4]
  assign x356_rdrow_1_clock = clock; // @[:@28612.4]
  assign x356_rdrow_1_reset = reset; // @[:@28613.4]
  assign x356_rdrow_1_io_a = RetimeWrapper_14_io_out; // @[Math.scala 192:17:@28614.4]
  assign x356_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@28615.4]
  assign x356_rdrow_1_io_flow = io_in_x279_TREADY; // @[Math.scala 194:20:@28616.4]
  assign RetimeWrapper_52_clock = clock; // @[:@28629.4]
  assign RetimeWrapper_52_reset = reset; // @[:@28630.4]
  assign RetimeWrapper_52_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@28633.4]
  assign RetimeWrapper_52_io_in = $unsigned(_T_1224); // @[package.scala 94:16:@28632.4]
  assign RetimeWrapper_53_clock = clock; // @[:@28647.4]
  assign RetimeWrapper_53_reset = reset; // @[:@28648.4]
  assign RetimeWrapper_53_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@28650.4]
  assign RetimeWrapper_53_io_in = $signed(_T_1221) < $signed(32'sh0); // @[package.scala 94:16:@28649.4]
  assign RetimeWrapper_54_clock = clock; // @[:@28656.4]
  assign RetimeWrapper_54_reset = reset; // @[:@28657.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28659.4]
  assign RetimeWrapper_54_io_in = RetimeWrapper_18_io_out; // @[package.scala 94:16:@28658.4]
  assign x550_sum_1_clock = clock; // @[:@28701.4]
  assign x550_sum_1_reset = reset; // @[:@28702.4]
  assign x550_sum_1_io_a = _T_1272[31:0]; // @[Math.scala 151:17:@28703.4]
  assign x550_sum_1_io_b = _T_1276[31:0]; // @[Math.scala 152:17:@28704.4]
  assign x550_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@28705.4]
  assign RetimeWrapper_55_clock = clock; // @[:@28711.4]
  assign RetimeWrapper_55_reset = reset; // @[:@28712.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28714.4]
  assign RetimeWrapper_55_io_in = x550_sum_1_io_result; // @[package.scala 94:16:@28713.4]
  assign x364_sum_1_clock = clock; // @[:@28720.4]
  assign x364_sum_1_reset = reset; // @[:@28721.4]
  assign x364_sum_1_io_a = RetimeWrapper_55_io_out; // @[Math.scala 151:17:@28722.4]
  assign x364_sum_1_io_b = RetimeWrapper_20_io_out; // @[Math.scala 152:17:@28723.4]
  assign x364_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@28724.4]
  assign RetimeWrapper_56_clock = clock; // @[:@28730.4]
  assign RetimeWrapper_56_reset = reset; // @[:@28731.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28733.4]
  assign RetimeWrapper_56_io_in = $unsigned(_T_1257); // @[package.scala 94:16:@28732.4]
  assign RetimeWrapper_57_clock = clock; // @[:@28739.4]
  assign RetimeWrapper_57_reset = reset; // @[:@28740.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28742.4]
  assign RetimeWrapper_57_io_in = ~ x359; // @[package.scala 94:16:@28741.4]
  assign RetimeWrapper_58_clock = clock; // @[:@28748.4]
  assign RetimeWrapper_58_reset = reset; // @[:@28749.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28751.4]
  assign RetimeWrapper_58_io_in = x364_sum_1_io_result; // @[package.scala 94:16:@28750.4]
  assign RetimeWrapper_59_clock = clock; // @[:@28760.4]
  assign RetimeWrapper_59_reset = reset; // @[:@28761.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28763.4]
  assign RetimeWrapper_59_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28762.4]
  assign RetimeWrapper_60_clock = clock; // @[:@28787.4]
  assign RetimeWrapper_60_reset = reset; // @[:@28788.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28790.4]
  assign RetimeWrapper_60_io_in = x550_sum_1_io_result; // @[package.scala 94:16:@28789.4]
  assign x369_sum_1_clock = clock; // @[:@28796.4]
  assign x369_sum_1_reset = reset; // @[:@28797.4]
  assign x369_sum_1_io_a = RetimeWrapper_60_io_out; // @[Math.scala 151:17:@28798.4]
  assign x369_sum_1_io_b = x343_div_1_io_result; // @[Math.scala 152:17:@28799.4]
  assign x369_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@28800.4]
  assign RetimeWrapper_61_clock = clock; // @[:@28806.4]
  assign RetimeWrapper_61_reset = reset; // @[:@28807.4]
  assign RetimeWrapper_61_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28809.4]
  assign RetimeWrapper_61_io_in = ~ x367; // @[package.scala 94:16:@28808.4]
  assign RetimeWrapper_62_clock = clock; // @[:@28818.4]
  assign RetimeWrapper_62_reset = reset; // @[:@28819.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28821.4]
  assign RetimeWrapper_62_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28820.4]
  assign x374_sum_1_clock = clock; // @[:@28845.4]
  assign x374_sum_1_reset = reset; // @[:@28846.4]
  assign x374_sum_1_io_a = RetimeWrapper_60_io_out; // @[Math.scala 151:17:@28847.4]
  assign x374_sum_1_io_b = x352_div_1_io_result; // @[Math.scala 152:17:@28848.4]
  assign x374_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@28849.4]
  assign RetimeWrapper_63_clock = clock; // @[:@28855.4]
  assign RetimeWrapper_63_reset = reset; // @[:@28856.4]
  assign RetimeWrapper_63_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28858.4]
  assign RetimeWrapper_63_io_in = ~ x372; // @[package.scala 94:16:@28857.4]
  assign RetimeWrapper_64_clock = clock; // @[:@28867.4]
  assign RetimeWrapper_64_reset = reset; // @[:@28868.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28870.4]
  assign RetimeWrapper_64_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@28869.4]
  assign x377_rdrow_1_clock = clock; // @[:@28890.4]
  assign x377_rdrow_1_reset = reset; // @[:@28891.4]
  assign x377_rdrow_1_io_a = RetimeWrapper_14_io_out; // @[Math.scala 192:17:@28892.4]
  assign x377_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@28893.4]
  assign x377_rdrow_1_io_flow = io_in_x279_TREADY; // @[Math.scala 194:20:@28894.4]
  assign RetimeWrapper_65_clock = clock; // @[:@28907.4]
  assign RetimeWrapper_65_reset = reset; // @[:@28908.4]
  assign RetimeWrapper_65_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@28911.4]
  assign RetimeWrapper_65_io_in = $unsigned(_T_1392); // @[package.scala 94:16:@28910.4]
  assign RetimeWrapper_66_clock = clock; // @[:@28925.4]
  assign RetimeWrapper_66_reset = reset; // @[:@28926.4]
  assign RetimeWrapper_66_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@28928.4]
  assign RetimeWrapper_66_io_in = $signed(_T_1389) < $signed(32'sh0); // @[package.scala 94:16:@28927.4]
  assign x555_sum_1_clock = clock; // @[:@28970.4]
  assign x555_sum_1_reset = reset; // @[:@28971.4]
  assign x555_sum_1_io_a = _T_1437[31:0]; // @[Math.scala 151:17:@28972.4]
  assign x555_sum_1_io_b = _T_1441[31:0]; // @[Math.scala 152:17:@28973.4]
  assign x555_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@28974.4]
  assign RetimeWrapper_67_clock = clock; // @[:@28980.4]
  assign RetimeWrapper_67_reset = reset; // @[:@28981.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@28983.4]
  assign RetimeWrapper_67_io_in = x555_sum_1_io_result; // @[package.scala 94:16:@28982.4]
  assign x385_sum_1_clock = clock; // @[:@28989.4]
  assign x385_sum_1_reset = reset; // @[:@28990.4]
  assign x385_sum_1_io_a = RetimeWrapper_67_io_out; // @[Math.scala 151:17:@28991.4]
  assign x385_sum_1_io_b = RetimeWrapper_20_io_out; // @[Math.scala 152:17:@28992.4]
  assign x385_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@28993.4]
  assign RetimeWrapper_68_clock = clock; // @[:@28999.4]
  assign RetimeWrapper_68_reset = reset; // @[:@29000.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29002.4]
  assign RetimeWrapper_68_io_in = x385_sum_1_io_result; // @[package.scala 94:16:@29001.4]
  assign RetimeWrapper_69_clock = clock; // @[:@29008.4]
  assign RetimeWrapper_69_reset = reset; // @[:@29009.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29011.4]
  assign RetimeWrapper_69_io_in = ~ x380; // @[package.scala 94:16:@29010.4]
  assign RetimeWrapper_70_clock = clock; // @[:@29017.4]
  assign RetimeWrapper_70_reset = reset; // @[:@29018.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29020.4]
  assign RetimeWrapper_70_io_in = $unsigned(_T_1422); // @[package.scala 94:16:@29019.4]
  assign RetimeWrapper_71_clock = clock; // @[:@29029.4]
  assign RetimeWrapper_71_reset = reset; // @[:@29030.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29032.4]
  assign RetimeWrapper_71_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@29031.4]
  assign RetimeWrapper_72_clock = clock; // @[:@29056.4]
  assign RetimeWrapper_72_reset = reset; // @[:@29057.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29059.4]
  assign RetimeWrapper_72_io_in = x555_sum_1_io_result; // @[package.scala 94:16:@29058.4]
  assign x390_sum_1_clock = clock; // @[:@29067.4]
  assign x390_sum_1_reset = reset; // @[:@29068.4]
  assign x390_sum_1_io_a = RetimeWrapper_72_io_out; // @[Math.scala 151:17:@29069.4]
  assign x390_sum_1_io_b = x343_div_1_io_result; // @[Math.scala 152:17:@29070.4]
  assign x390_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@29071.4]
  assign RetimeWrapper_73_clock = clock; // @[:@29077.4]
  assign RetimeWrapper_73_reset = reset; // @[:@29078.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29080.4]
  assign RetimeWrapper_73_io_in = ~ x388; // @[package.scala 94:16:@29079.4]
  assign RetimeWrapper_74_clock = clock; // @[:@29089.4]
  assign RetimeWrapper_74_reset = reset; // @[:@29090.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29092.4]
  assign RetimeWrapper_74_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@29091.4]
  assign x395_sum_1_clock = clock; // @[:@29116.4]
  assign x395_sum_1_reset = reset; // @[:@29117.4]
  assign x395_sum_1_io_a = RetimeWrapper_72_io_out; // @[Math.scala 151:17:@29118.4]
  assign x395_sum_1_io_b = x352_div_1_io_result; // @[Math.scala 152:17:@29119.4]
  assign x395_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@29120.4]
  assign RetimeWrapper_75_clock = clock; // @[:@29126.4]
  assign RetimeWrapper_75_reset = reset; // @[:@29127.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29129.4]
  assign RetimeWrapper_75_io_in = ~ x393; // @[package.scala 94:16:@29128.4]
  assign RetimeWrapper_76_clock = clock; // @[:@29138.4]
  assign RetimeWrapper_76_reset = reset; // @[:@29139.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29141.4]
  assign RetimeWrapper_76_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@29140.4]
  assign RetimeWrapper_77_clock = clock; // @[:@29161.4]
  assign RetimeWrapper_77_reset = reset; // @[:@29162.4]
  assign RetimeWrapper_77_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@29164.4]
  assign RetimeWrapper_77_io_in = _GEN_8 << 1; // @[package.scala 94:16:@29163.4]
  assign RetimeWrapper_78_clock = clock; // @[:@29173.4]
  assign RetimeWrapper_78_reset = reset; // @[:@29174.4]
  assign RetimeWrapper_78_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@29176.4]
  assign RetimeWrapper_78_io_in = _GEN_9 << 1; // @[package.scala 94:16:@29175.4]
  assign RetimeWrapper_79_clock = clock; // @[:@29185.4]
  assign RetimeWrapper_79_reset = reset; // @[:@29186.4]
  assign RetimeWrapper_79_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@29188.4]
  assign RetimeWrapper_79_io_in = _GEN_10 << 2; // @[package.scala 94:16:@29187.4]
  assign RetimeWrapper_80_clock = clock; // @[:@29197.4]
  assign RetimeWrapper_80_reset = reset; // @[:@29198.4]
  assign RetimeWrapper_80_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@29200.4]
  assign RetimeWrapper_80_io_in = _GEN_11 << 1; // @[package.scala 94:16:@29199.4]
  assign RetimeWrapper_81_clock = clock; // @[:@29209.4]
  assign RetimeWrapper_81_reset = reset; // @[:@29210.4]
  assign RetimeWrapper_81_io_flow = io_in_x279_TREADY; // @[package.scala 95:18:@29212.4]
  assign RetimeWrapper_81_io_in = _GEN_12 << 1; // @[package.scala 94:16:@29211.4]
  assign RetimeWrapper_82_clock = clock; // @[:@29219.4]
  assign RetimeWrapper_82_reset = reset; // @[:@29220.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29222.4]
  assign RetimeWrapper_82_io_in = x311_lb_0_io_rPort_6_output_0; // @[package.scala 94:16:@29221.4]
  assign x403_x15_1_io_a = RetimeWrapper_82_io_out; // @[Math.scala 151:17:@29230.4]
  assign x403_x15_1_io_b = _T_1547[7:0]; // @[Math.scala 152:17:@29231.4]
  assign RetimeWrapper_83_clock = clock; // @[:@29238.4]
  assign RetimeWrapper_83_reset = reset; // @[:@29239.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29241.4]
  assign RetimeWrapper_83_io_in = x311_lb_0_io_rPort_8_output_0; // @[package.scala 94:16:@29240.4]
  assign x404_x16_1_io_a = RetimeWrapper_83_io_out; // @[Math.scala 151:17:@29249.4]
  assign x404_x16_1_io_b = _T_1553[7:0]; // @[Math.scala 152:17:@29250.4]
  assign x405_x15_1_io_a = _T_1559[7:0]; // @[Math.scala 151:17:@29259.4]
  assign x405_x15_1_io_b = _T_1565[7:0]; // @[Math.scala 152:17:@29260.4]
  assign RetimeWrapper_84_clock = clock; // @[:@29267.4]
  assign RetimeWrapper_84_reset = reset; // @[:@29268.4]
  assign RetimeWrapper_84_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29270.4]
  assign RetimeWrapper_84_io_in = x311_lb_0_io_rPort_7_output_0; // @[package.scala 94:16:@29269.4]
  assign x406_x16_1_io_a = RetimeWrapper_84_io_out; // @[Math.scala 151:17:@29278.4]
  assign x406_x16_1_io_b = _T_1571[7:0]; // @[Math.scala 152:17:@29279.4]
  assign x407_x15_1_io_a = x403_x15_1_io_result; // @[Math.scala 151:17:@29288.4]
  assign x407_x15_1_io_b = x404_x16_1_io_result; // @[Math.scala 152:17:@29289.4]
  assign x408_x16_1_io_a = x405_x15_1_io_result; // @[Math.scala 151:17:@29298.4]
  assign x408_x16_1_io_b = x406_x16_1_io_result; // @[Math.scala 152:17:@29299.4]
  assign x409_x15_1_io_a = x407_x15_1_io_result; // @[Math.scala 151:17:@29308.4]
  assign x409_x15_1_io_b = x408_x16_1_io_result; // @[Math.scala 152:17:@29309.4]
  assign RetimeWrapper_85_clock = clock; // @[:@29316.4]
  assign RetimeWrapper_85_reset = reset; // @[:@29317.4]
  assign RetimeWrapper_85_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29319.4]
  assign RetimeWrapper_85_io_in = x311_lb_0_io_rPort_1_output_0; // @[package.scala 94:16:@29318.4]
  assign x410_sum_1_clock = clock; // @[:@29325.4]
  assign x410_sum_1_reset = reset; // @[:@29326.4]
  assign x410_sum_1_io_a = x409_x15_1_io_result; // @[Math.scala 151:17:@29327.4]
  assign x410_sum_1_io_b = RetimeWrapper_85_io_out; // @[Math.scala 152:17:@29328.4]
  assign x410_sum_1_io_flow = io_in_x279_TREADY; // @[Math.scala 153:20:@29329.4]
  assign RetimeWrapper_86_clock = clock; // @[:@29346.4]
  assign RetimeWrapper_86_reset = reset; // @[:@29347.4]
  assign RetimeWrapper_86_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29349.4]
  assign RetimeWrapper_86_io_in = {4'h0,_T_1616}; // @[package.scala 94:16:@29348.4]
  assign RetimeWrapper_87_clock = clock; // @[:@29355.4]
  assign RetimeWrapper_87_reset = reset; // @[:@29356.4]
  assign RetimeWrapper_87_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29358.4]
  assign RetimeWrapper_87_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@29357.4]
  assign RetimeWrapper_88_clock = clock; // @[:@29364.4]
  assign RetimeWrapper_88_reset = reset; // @[:@29365.4]
  assign RetimeWrapper_88_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29367.4]
  assign RetimeWrapper_88_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@29366.4]
  assign RetimeWrapper_89_clock = clock; // @[:@29373.4]
  assign RetimeWrapper_89_reset = reset; // @[:@29374.4]
  assign RetimeWrapper_89_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@29376.4]
  assign RetimeWrapper_89_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@29375.4]
endmodule
module x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1( // @[:@29394.2]
  input          clock, // @[:@29395.4]
  input          reset, // @[:@29396.4]
  output         io_in_x279_TVALID, // @[:@29397.4]
  input          io_in_x279_TREADY, // @[:@29397.4]
  output [255:0] io_in_x279_TDATA, // @[:@29397.4]
  input          io_in_x278_TVALID, // @[:@29397.4]
  output         io_in_x278_TREADY, // @[:@29397.4]
  input  [255:0] io_in_x278_TDATA, // @[:@29397.4]
  input  [7:0]   io_in_x278_TID, // @[:@29397.4]
  input  [7:0]   io_in_x278_TDEST, // @[:@29397.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@29397.4]
  input          io_sigsIn_smChildAcks_0, // @[:@29397.4]
  output         io_sigsOut_smDoneIn_0, // @[:@29397.4]
  input          io_rr // @[:@29397.4]
);
  wire  x304_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@29431.4]
  wire  x304_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@29431.4]
  wire  x304_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@29431.4]
  wire  x304_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@29431.4]
  wire [12:0] x304_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@29431.4]
  wire [12:0] x304_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@29431.4]
  wire  x304_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@29431.4]
  wire  x304_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@29431.4]
  wire  x304_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@29431.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 32:18:@29491.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 32:18:@29491.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 32:18:@29491.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 32:18:@29491.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 32:18:@29491.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 32:18:@29491.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 32:18:@29491.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 32:18:@29491.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 32:18:@29491.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 32:18:@29491.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 32:18:@29491.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 32:18:@29491.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@29519.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@29519.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@29519.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@29519.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@29519.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@29561.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@29561.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@29561.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@29561.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@29561.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@29569.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@29569.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@29569.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@29569.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@29569.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 604:24:@29603.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 604:24:@29603.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x279_TVALID; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 604:24:@29603.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x279_TREADY; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 604:24:@29603.4]
  wire [255:0] x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x279_TDATA; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 604:24:@29603.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x278_TREADY; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 604:24:@29603.4]
  wire [255:0] x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x278_TDATA; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 604:24:@29603.4]
  wire [7:0] x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x278_TID; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 604:24:@29603.4]
  wire [7:0] x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x278_TDEST; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 604:24:@29603.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 604:24:@29603.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 604:24:@29603.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 604:24:@29603.4]
  wire [31:0] x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 604:24:@29603.4]
  wire [31:0] x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 604:24:@29603.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 604:24:@29603.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 604:24:@29603.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 604:24:@29603.4]
  wire  _T_240; // @[package.scala 96:25:@29524.4 package.scala 96:25:@29525.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x417_outr_UnitPipe.scala 69:66:@29530.4]
  wire  _T_253; // @[package.scala 96:25:@29566.4 package.scala 96:25:@29567.4]
  wire  _T_259; // @[package.scala 96:25:@29574.4 package.scala 96:25:@29575.4]
  wire  _T_262; // @[SpatialBlocks.scala 138:93:@29577.4]
  wire  x416_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@29578.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:36:@29586.4]
  wire  _T_265; // @[SpatialBlocks.scala 157:78:@29587.4]
  wire  _T_272; // @[SpatialBlocks.scala 159:58:@29599.4]
  x286_ctrchain x304_ctrchain ( // @[SpatialBlocks.scala 37:22:@29431.4]
    .clock(x304_ctrchain_clock),
    .reset(x304_ctrchain_reset),
    .io_input_reset(x304_ctrchain_io_input_reset),
    .io_input_enable(x304_ctrchain_io_input_enable),
    .io_output_counts_1(x304_ctrchain_io_output_counts_1),
    .io_output_counts_0(x304_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x304_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x304_ctrchain_io_output_oobs_1),
    .io_output_done(x304_ctrchain_io_output_done)
  );
  x416_inr_Foreach_SAMPLER_BOX_sm x416_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 32:18:@29491.4]
    .clock(x416_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x416_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x416_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x416_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x416_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x416_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x416_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x416_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x416_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x416_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x416_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x416_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@29519.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@29561.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@29569.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1 x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 604:24:@29603.4]
    .clock(x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x279_TVALID(x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x279_TVALID),
    .io_in_x279_TREADY(x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x279_TREADY),
    .io_in_x279_TDATA(x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x279_TDATA),
    .io_in_x278_TREADY(x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x278_TREADY),
    .io_in_x278_TDATA(x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x278_TDATA),
    .io_in_x278_TID(x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x278_TID),
    .io_in_x278_TDEST(x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x278_TDEST),
    .io_sigsIn_backpressure(x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_240 = RetimeWrapper_io_out; // @[package.scala 96:25:@29524.4 package.scala 96:25:@29525.4]
  assign x416_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x278_TVALID | x416_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x417_outr_UnitPipe.scala 69:66:@29530.4]
  assign _T_253 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@29566.4 package.scala 96:25:@29567.4]
  assign _T_259 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@29574.4 package.scala 96:25:@29575.4]
  assign _T_262 = ~ _T_259; // @[SpatialBlocks.scala 138:93:@29577.4]
  assign x416_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_253 & _T_262; // @[SpatialBlocks.scala 138:90:@29578.4]
  assign _T_264 = x416_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@29586.4]
  assign _T_265 = ~ x416_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@29587.4]
  assign _T_272 = x416_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@29599.4]
  assign io_in_x279_TVALID = x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x279_TVALID; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 48:23:@29662.4]
  assign io_in_x279_TDATA = x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x279_TDATA; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 48:23:@29660.4]
  assign io_in_x278_TREADY = x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x278_TREADY; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 49:23:@29670.4]
  assign io_sigsOut_smDoneIn_0 = x416_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@29584.4]
  assign x304_ctrchain_clock = clock; // @[:@29432.4]
  assign x304_ctrchain_reset = reset; // @[:@29433.4]
  assign x304_ctrchain_io_input_reset = x416_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@29602.4]
  assign x304_ctrchain_io_input_enable = _T_272 & x416_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@29554.4 SpatialBlocks.scala 159:42:@29601.4]
  assign x416_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@29492.4]
  assign x416_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@29493.4]
  assign x416_inr_Foreach_SAMPLER_BOX_sm_io_enable = x416_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x416_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@29581.4]
  assign x416_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_240 : 1'h0; // @[sm_x417_outr_UnitPipe.scala 67:50:@29527.4]
  assign x416_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@29583.4]
  assign x416_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x279_TREADY | x416_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@29555.4]
  assign x416_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x417_outr_UnitPipe.scala 71:48:@29533.4]
  assign RetimeWrapper_clock = clock; // @[:@29520.4]
  assign RetimeWrapper_reset = reset; // @[:@29521.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@29523.4]
  assign RetimeWrapper_io_in = x304_ctrchain_io_output_done; // @[package.scala 94:16:@29522.4]
  assign RetimeWrapper_1_clock = clock; // @[:@29562.4]
  assign RetimeWrapper_1_reset = reset; // @[:@29563.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@29565.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@29564.4]
  assign RetimeWrapper_2_clock = clock; // @[:@29570.4]
  assign RetimeWrapper_2_reset = reset; // @[:@29571.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@29573.4]
  assign RetimeWrapper_2_io_in = x416_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@29572.4]
  assign x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@29604.4]
  assign x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@29605.4]
  assign x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x279_TREADY = io_in_x279_TREADY; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 48:23:@29661.4]
  assign x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x278_TDATA = io_in_x278_TDATA; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 49:23:@29669.4]
  assign x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x278_TID = io_in_x278_TID; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 49:23:@29665.4]
  assign x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x278_TDEST = io_in_x278_TDEST; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 49:23:@29664.4]
  assign x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x279_TREADY | x416_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 609:22:@29688.4]
  assign x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_264 & _T_265; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 609:22:@29686.4]
  assign x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x416_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 609:22:@29684.4]
  assign x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x304_ctrchain_io_output_counts_1[12]}},x304_ctrchain_io_output_counts_1}; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 609:22:@29679.4]
  assign x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x304_ctrchain_io_output_counts_0[12]}},x304_ctrchain_io_output_counts_0}; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 609:22:@29678.4]
  assign x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x304_ctrchain_io_output_oobs_0; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 609:22:@29676.4]
  assign x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x304_ctrchain_io_output_oobs_1; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 609:22:@29677.4]
  assign x416_inr_Foreach_SAMPLER_BOX_kernelx416_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x416_inr_Foreach_SAMPLER_BOX.scala 608:18:@29672.4]
endmodule
module x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1( // @[:@29702.2]
  input          clock, // @[:@29703.4]
  input          reset, // @[:@29704.4]
  output         io_in_x279_TVALID, // @[:@29705.4]
  input          io_in_x279_TREADY, // @[:@29705.4]
  output [255:0] io_in_x279_TDATA, // @[:@29705.4]
  input          io_in_x278_TVALID, // @[:@29705.4]
  output         io_in_x278_TREADY, // @[:@29705.4]
  input  [255:0] io_in_x278_TDATA, // @[:@29705.4]
  input  [7:0]   io_in_x278_TID, // @[:@29705.4]
  input  [7:0]   io_in_x278_TDEST, // @[:@29705.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@29705.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@29705.4]
  input          io_sigsIn_smChildAcks_0, // @[:@29705.4]
  input          io_sigsIn_smChildAcks_1, // @[:@29705.4]
  output         io_sigsOut_smDoneIn_0, // @[:@29705.4]
  output         io_sigsOut_smDoneIn_1, // @[:@29705.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@29705.4]
  output         io_sigsOut_smCtrCopyDone_1, // @[:@29705.4]
  input          io_rr // @[:@29705.4]
);
  wire  x281_fifoinraw_0_clock; // @[m_x281_fifoinraw_0.scala 27:17:@29719.4]
  wire  x281_fifoinraw_0_reset; // @[m_x281_fifoinraw_0.scala 27:17:@29719.4]
  wire  x282_fifoinpacked_0_clock; // @[m_x282_fifoinpacked_0.scala 27:17:@29743.4]
  wire  x282_fifoinpacked_0_reset; // @[m_x282_fifoinpacked_0.scala 27:17:@29743.4]
  wire  x282_fifoinpacked_0_io_wPort_0_en_0; // @[m_x282_fifoinpacked_0.scala 27:17:@29743.4]
  wire  x282_fifoinpacked_0_io_full; // @[m_x282_fifoinpacked_0.scala 27:17:@29743.4]
  wire  x282_fifoinpacked_0_io_active_0_in; // @[m_x282_fifoinpacked_0.scala 27:17:@29743.4]
  wire  x282_fifoinpacked_0_io_active_0_out; // @[m_x282_fifoinpacked_0.scala 27:17:@29743.4]
  wire  x283_fifooutraw_0_clock; // @[m_x283_fifooutraw_0.scala 27:17:@29767.4]
  wire  x283_fifooutraw_0_reset; // @[m_x283_fifooutraw_0.scala 27:17:@29767.4]
  wire  x286_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@29791.4]
  wire  x286_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@29791.4]
  wire  x286_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@29791.4]
  wire  x286_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@29791.4]
  wire [12:0] x286_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@29791.4]
  wire [12:0] x286_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@29791.4]
  wire  x286_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@29791.4]
  wire  x286_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@29791.4]
  wire  x286_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@29791.4]
  wire  x300_inr_Foreach_sm_clock; // @[sm_x300_inr_Foreach.scala 32:18:@29851.4]
  wire  x300_inr_Foreach_sm_reset; // @[sm_x300_inr_Foreach.scala 32:18:@29851.4]
  wire  x300_inr_Foreach_sm_io_enable; // @[sm_x300_inr_Foreach.scala 32:18:@29851.4]
  wire  x300_inr_Foreach_sm_io_done; // @[sm_x300_inr_Foreach.scala 32:18:@29851.4]
  wire  x300_inr_Foreach_sm_io_doneLatch; // @[sm_x300_inr_Foreach.scala 32:18:@29851.4]
  wire  x300_inr_Foreach_sm_io_ctrDone; // @[sm_x300_inr_Foreach.scala 32:18:@29851.4]
  wire  x300_inr_Foreach_sm_io_datapathEn; // @[sm_x300_inr_Foreach.scala 32:18:@29851.4]
  wire  x300_inr_Foreach_sm_io_ctrInc; // @[sm_x300_inr_Foreach.scala 32:18:@29851.4]
  wire  x300_inr_Foreach_sm_io_ctrRst; // @[sm_x300_inr_Foreach.scala 32:18:@29851.4]
  wire  x300_inr_Foreach_sm_io_parentAck; // @[sm_x300_inr_Foreach.scala 32:18:@29851.4]
  wire  x300_inr_Foreach_sm_io_backpressure; // @[sm_x300_inr_Foreach.scala 32:18:@29851.4]
  wire  x300_inr_Foreach_sm_io_break; // @[sm_x300_inr_Foreach.scala 32:18:@29851.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@29879.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@29879.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@29879.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@29879.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@29879.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@29925.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@29925.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@29925.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@29925.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@29925.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@29933.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@29933.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@29933.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@29933.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@29933.4]
  wire  x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_clock; // @[sm_x300_inr_Foreach.scala 96:24:@29968.4]
  wire  x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_reset; // @[sm_x300_inr_Foreach.scala 96:24:@29968.4]
  wire  x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_in_x282_fifoinpacked_0_wPort_0_en_0; // @[sm_x300_inr_Foreach.scala 96:24:@29968.4]
  wire  x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_in_x282_fifoinpacked_0_full; // @[sm_x300_inr_Foreach.scala 96:24:@29968.4]
  wire  x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_in_x282_fifoinpacked_0_active_0_in; // @[sm_x300_inr_Foreach.scala 96:24:@29968.4]
  wire  x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_in_x282_fifoinpacked_0_active_0_out; // @[sm_x300_inr_Foreach.scala 96:24:@29968.4]
  wire  x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x300_inr_Foreach.scala 96:24:@29968.4]
  wire  x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x300_inr_Foreach.scala 96:24:@29968.4]
  wire  x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x300_inr_Foreach.scala 96:24:@29968.4]
  wire [31:0] x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x300_inr_Foreach.scala 96:24:@29968.4]
  wire [31:0] x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x300_inr_Foreach.scala 96:24:@29968.4]
  wire  x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x300_inr_Foreach.scala 96:24:@29968.4]
  wire  x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x300_inr_Foreach.scala 96:24:@29968.4]
  wire  x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_rr; // @[sm_x300_inr_Foreach.scala 96:24:@29968.4]
  wire  x417_outr_UnitPipe_sm_clock; // @[sm_x417_outr_UnitPipe.scala 32:18:@30100.4]
  wire  x417_outr_UnitPipe_sm_reset; // @[sm_x417_outr_UnitPipe.scala 32:18:@30100.4]
  wire  x417_outr_UnitPipe_sm_io_enable; // @[sm_x417_outr_UnitPipe.scala 32:18:@30100.4]
  wire  x417_outr_UnitPipe_sm_io_done; // @[sm_x417_outr_UnitPipe.scala 32:18:@30100.4]
  wire  x417_outr_UnitPipe_sm_io_rst; // @[sm_x417_outr_UnitPipe.scala 32:18:@30100.4]
  wire  x417_outr_UnitPipe_sm_io_ctrDone; // @[sm_x417_outr_UnitPipe.scala 32:18:@30100.4]
  wire  x417_outr_UnitPipe_sm_io_ctrInc; // @[sm_x417_outr_UnitPipe.scala 32:18:@30100.4]
  wire  x417_outr_UnitPipe_sm_io_parentAck; // @[sm_x417_outr_UnitPipe.scala 32:18:@30100.4]
  wire  x417_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x417_outr_UnitPipe.scala 32:18:@30100.4]
  wire  x417_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x417_outr_UnitPipe.scala 32:18:@30100.4]
  wire  x417_outr_UnitPipe_sm_io_childAck_0; // @[sm_x417_outr_UnitPipe.scala 32:18:@30100.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@30157.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@30157.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@30157.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@30157.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@30157.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@30165.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@30165.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@30165.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@30165.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@30165.4]
  wire  x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_clock; // @[sm_x417_outr_UnitPipe.scala 76:24:@30195.4]
  wire  x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_reset; // @[sm_x417_outr_UnitPipe.scala 76:24:@30195.4]
  wire  x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x279_TVALID; // @[sm_x417_outr_UnitPipe.scala 76:24:@30195.4]
  wire  x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x279_TREADY; // @[sm_x417_outr_UnitPipe.scala 76:24:@30195.4]
  wire [255:0] x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x279_TDATA; // @[sm_x417_outr_UnitPipe.scala 76:24:@30195.4]
  wire  x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x278_TVALID; // @[sm_x417_outr_UnitPipe.scala 76:24:@30195.4]
  wire  x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x278_TREADY; // @[sm_x417_outr_UnitPipe.scala 76:24:@30195.4]
  wire [255:0] x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x278_TDATA; // @[sm_x417_outr_UnitPipe.scala 76:24:@30195.4]
  wire [7:0] x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x278_TID; // @[sm_x417_outr_UnitPipe.scala 76:24:@30195.4]
  wire [7:0] x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x278_TDEST; // @[sm_x417_outr_UnitPipe.scala 76:24:@30195.4]
  wire  x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x417_outr_UnitPipe.scala 76:24:@30195.4]
  wire  x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x417_outr_UnitPipe.scala 76:24:@30195.4]
  wire  x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x417_outr_UnitPipe.scala 76:24:@30195.4]
  wire  x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_rr; // @[sm_x417_outr_UnitPipe.scala 76:24:@30195.4]
  wire  _T_254; // @[package.scala 96:25:@29884.4 package.scala 96:25:@29885.4]
  wire  _T_260; // @[implicits.scala 47:10:@29888.4]
  wire  _T_261; // @[sm_x418_outr_UnitPipe.scala 70:41:@29889.4]
  wire  _T_262; // @[sm_x418_outr_UnitPipe.scala 70:78:@29890.4]
  wire  _T_263; // @[sm_x418_outr_UnitPipe.scala 70:76:@29891.4]
  wire  _T_275; // @[package.scala 96:25:@29930.4 package.scala 96:25:@29931.4]
  wire  _T_281; // @[package.scala 96:25:@29938.4 package.scala 96:25:@29939.4]
  wire  _T_284; // @[SpatialBlocks.scala 138:93:@29941.4]
  wire  _T_286; // @[SpatialBlocks.scala 157:36:@29950.4]
  wire  _T_287; // @[SpatialBlocks.scala 157:78:@29951.4]
  wire  _T_354; // @[package.scala 100:49:@30128.4]
  reg  _T_357; // @[package.scala 48:56:@30129.4]
  reg [31:0] _RAND_0;
  wire  _T_371; // @[package.scala 96:25:@30162.4 package.scala 96:25:@30163.4]
  wire  _T_377; // @[package.scala 96:25:@30170.4 package.scala 96:25:@30171.4]
  wire  _T_380; // @[SpatialBlocks.scala 138:93:@30173.4]
  x281_fifoinraw_0 x281_fifoinraw_0 ( // @[m_x281_fifoinraw_0.scala 27:17:@29719.4]
    .clock(x281_fifoinraw_0_clock),
    .reset(x281_fifoinraw_0_reset)
  );
  x282_fifoinpacked_0 x282_fifoinpacked_0 ( // @[m_x282_fifoinpacked_0.scala 27:17:@29743.4]
    .clock(x282_fifoinpacked_0_clock),
    .reset(x282_fifoinpacked_0_reset),
    .io_wPort_0_en_0(x282_fifoinpacked_0_io_wPort_0_en_0),
    .io_full(x282_fifoinpacked_0_io_full),
    .io_active_0_in(x282_fifoinpacked_0_io_active_0_in),
    .io_active_0_out(x282_fifoinpacked_0_io_active_0_out)
  );
  x281_fifoinraw_0 x283_fifooutraw_0 ( // @[m_x283_fifooutraw_0.scala 27:17:@29767.4]
    .clock(x283_fifooutraw_0_clock),
    .reset(x283_fifooutraw_0_reset)
  );
  x286_ctrchain x286_ctrchain ( // @[SpatialBlocks.scala 37:22:@29791.4]
    .clock(x286_ctrchain_clock),
    .reset(x286_ctrchain_reset),
    .io_input_reset(x286_ctrchain_io_input_reset),
    .io_input_enable(x286_ctrchain_io_input_enable),
    .io_output_counts_1(x286_ctrchain_io_output_counts_1),
    .io_output_counts_0(x286_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x286_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x286_ctrchain_io_output_oobs_1),
    .io_output_done(x286_ctrchain_io_output_done)
  );
  x300_inr_Foreach_sm x300_inr_Foreach_sm ( // @[sm_x300_inr_Foreach.scala 32:18:@29851.4]
    .clock(x300_inr_Foreach_sm_clock),
    .reset(x300_inr_Foreach_sm_reset),
    .io_enable(x300_inr_Foreach_sm_io_enable),
    .io_done(x300_inr_Foreach_sm_io_done),
    .io_doneLatch(x300_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x300_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x300_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x300_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x300_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x300_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x300_inr_Foreach_sm_io_backpressure),
    .io_break(x300_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@29879.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@29925.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@29933.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x300_inr_Foreach_kernelx300_inr_Foreach_concrete1 x300_inr_Foreach_kernelx300_inr_Foreach_concrete1 ( // @[sm_x300_inr_Foreach.scala 96:24:@29968.4]
    .clock(x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_clock),
    .reset(x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_reset),
    .io_in_x282_fifoinpacked_0_wPort_0_en_0(x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_in_x282_fifoinpacked_0_wPort_0_en_0),
    .io_in_x282_fifoinpacked_0_full(x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_in_x282_fifoinpacked_0_full),
    .io_in_x282_fifoinpacked_0_active_0_in(x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_in_x282_fifoinpacked_0_active_0_in),
    .io_in_x282_fifoinpacked_0_active_0_out(x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_in_x282_fifoinpacked_0_active_0_out),
    .io_sigsIn_backpressure(x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_rr)
  );
  RootController_sm x417_outr_UnitPipe_sm ( // @[sm_x417_outr_UnitPipe.scala 32:18:@30100.4]
    .clock(x417_outr_UnitPipe_sm_clock),
    .reset(x417_outr_UnitPipe_sm_reset),
    .io_enable(x417_outr_UnitPipe_sm_io_enable),
    .io_done(x417_outr_UnitPipe_sm_io_done),
    .io_rst(x417_outr_UnitPipe_sm_io_rst),
    .io_ctrDone(x417_outr_UnitPipe_sm_io_ctrDone),
    .io_ctrInc(x417_outr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x417_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x417_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x417_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x417_outr_UnitPipe_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@30157.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@30165.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1 x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1 ( // @[sm_x417_outr_UnitPipe.scala 76:24:@30195.4]
    .clock(x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_clock),
    .reset(x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_reset),
    .io_in_x279_TVALID(x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x279_TVALID),
    .io_in_x279_TREADY(x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x279_TREADY),
    .io_in_x279_TDATA(x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x279_TDATA),
    .io_in_x278_TVALID(x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x278_TVALID),
    .io_in_x278_TREADY(x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x278_TREADY),
    .io_in_x278_TDATA(x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x278_TDATA),
    .io_in_x278_TID(x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x278_TID),
    .io_in_x278_TDEST(x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x278_TDEST),
    .io_sigsIn_smEnableOuts_0(x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_254 = RetimeWrapper_io_out; // @[package.scala 96:25:@29884.4 package.scala 96:25:@29885.4]
  assign _T_260 = x282_fifoinpacked_0_io_full; // @[implicits.scala 47:10:@29888.4]
  assign _T_261 = ~ _T_260; // @[sm_x418_outr_UnitPipe.scala 70:41:@29889.4]
  assign _T_262 = ~ x282_fifoinpacked_0_io_active_0_out; // @[sm_x418_outr_UnitPipe.scala 70:78:@29890.4]
  assign _T_263 = _T_261 | _T_262; // @[sm_x418_outr_UnitPipe.scala 70:76:@29891.4]
  assign _T_275 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@29930.4 package.scala 96:25:@29931.4]
  assign _T_281 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@29938.4 package.scala 96:25:@29939.4]
  assign _T_284 = ~ _T_281; // @[SpatialBlocks.scala 138:93:@29941.4]
  assign _T_286 = x300_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@29950.4]
  assign _T_287 = ~ x300_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@29951.4]
  assign _T_354 = x417_outr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@30128.4]
  assign _T_371 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@30162.4 package.scala 96:25:@30163.4]
  assign _T_377 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@30170.4 package.scala 96:25:@30171.4]
  assign _T_380 = ~ _T_377; // @[SpatialBlocks.scala 138:93:@30173.4]
  assign io_in_x279_TVALID = x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x279_TVALID; // @[sm_x417_outr_UnitPipe.scala 48:23:@30252.4]
  assign io_in_x279_TDATA = x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x279_TDATA; // @[sm_x417_outr_UnitPipe.scala 48:23:@30250.4]
  assign io_in_x278_TREADY = x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x278_TREADY; // @[sm_x417_outr_UnitPipe.scala 49:23:@30260.4]
  assign io_sigsOut_smDoneIn_0 = x300_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@29948.4]
  assign io_sigsOut_smDoneIn_1 = x417_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@30180.4]
  assign io_sigsOut_smCtrCopyDone_0 = x300_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@29967.4]
  assign io_sigsOut_smCtrCopyDone_1 = x417_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@30194.4]
  assign x281_fifoinraw_0_clock = clock; // @[:@29720.4]
  assign x281_fifoinraw_0_reset = reset; // @[:@29721.4]
  assign x282_fifoinpacked_0_clock = clock; // @[:@29744.4]
  assign x282_fifoinpacked_0_reset = reset; // @[:@29745.4]
  assign x282_fifoinpacked_0_io_wPort_0_en_0 = x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_in_x282_fifoinpacked_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@30028.4]
  assign x282_fifoinpacked_0_io_active_0_in = x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_in_x282_fifoinpacked_0_active_0_in; // @[MemInterfaceType.scala 167:86:@30027.4]
  assign x283_fifooutraw_0_clock = clock; // @[:@29768.4]
  assign x283_fifooutraw_0_reset = reset; // @[:@29769.4]
  assign x286_ctrchain_clock = clock; // @[:@29792.4]
  assign x286_ctrchain_reset = reset; // @[:@29793.4]
  assign x286_ctrchain_io_input_reset = x300_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@29966.4]
  assign x286_ctrchain_io_input_enable = x300_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@29918.4 SpatialBlocks.scala 159:42:@29965.4]
  assign x300_inr_Foreach_sm_clock = clock; // @[:@29852.4]
  assign x300_inr_Foreach_sm_reset = reset; // @[:@29853.4]
  assign x300_inr_Foreach_sm_io_enable = _T_275 & _T_284; // @[SpatialBlocks.scala 140:18:@29945.4]
  assign x300_inr_Foreach_sm_io_ctrDone = io_rr ? _T_254 : 1'h0; // @[sm_x418_outr_UnitPipe.scala 69:38:@29887.4]
  assign x300_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@29947.4]
  assign x300_inr_Foreach_sm_io_backpressure = _T_263 | x300_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@29919.4]
  assign x300_inr_Foreach_sm_io_break = 1'h0; // @[sm_x418_outr_UnitPipe.scala 73:36:@29897.4]
  assign RetimeWrapper_clock = clock; // @[:@29880.4]
  assign RetimeWrapper_reset = reset; // @[:@29881.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@29883.4]
  assign RetimeWrapper_io_in = x286_ctrchain_io_output_done; // @[package.scala 94:16:@29882.4]
  assign RetimeWrapper_1_clock = clock; // @[:@29926.4]
  assign RetimeWrapper_1_reset = reset; // @[:@29927.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@29929.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@29928.4]
  assign RetimeWrapper_2_clock = clock; // @[:@29934.4]
  assign RetimeWrapper_2_reset = reset; // @[:@29935.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@29937.4]
  assign RetimeWrapper_2_io_in = x300_inr_Foreach_sm_io_done; // @[package.scala 94:16:@29936.4]
  assign x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_clock = clock; // @[:@29969.4]
  assign x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_reset = reset; // @[:@29970.4]
  assign x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_in_x282_fifoinpacked_0_full = x282_fifoinpacked_0_io_full; // @[MemInterfaceType.scala 159:15:@30022.4]
  assign x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_in_x282_fifoinpacked_0_active_0_out = x282_fifoinpacked_0_io_active_0_out; // @[MemInterfaceType.scala 158:75:@30021.4]
  assign x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_263 | x300_inr_Foreach_sm_io_doneLatch; // @[sm_x300_inr_Foreach.scala 101:22:@30051.4]
  assign x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_286 & _T_287; // @[sm_x300_inr_Foreach.scala 101:22:@30049.4]
  assign x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_break = x300_inr_Foreach_sm_io_break; // @[sm_x300_inr_Foreach.scala 101:22:@30047.4]
  assign x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x286_ctrchain_io_output_counts_1[12]}},x286_ctrchain_io_output_counts_1}; // @[sm_x300_inr_Foreach.scala 101:22:@30042.4]
  assign x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x286_ctrchain_io_output_counts_0[12]}},x286_ctrchain_io_output_counts_0}; // @[sm_x300_inr_Foreach.scala 101:22:@30041.4]
  assign x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x286_ctrchain_io_output_oobs_0; // @[sm_x300_inr_Foreach.scala 101:22:@30039.4]
  assign x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x286_ctrchain_io_output_oobs_1; // @[sm_x300_inr_Foreach.scala 101:22:@30040.4]
  assign x300_inr_Foreach_kernelx300_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x300_inr_Foreach.scala 100:18:@30035.4]
  assign x417_outr_UnitPipe_sm_clock = clock; // @[:@30101.4]
  assign x417_outr_UnitPipe_sm_reset = reset; // @[:@30102.4]
  assign x417_outr_UnitPipe_sm_io_enable = _T_371 & _T_380; // @[SpatialBlocks.scala 140:18:@30177.4]
  assign x417_outr_UnitPipe_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 134:15:@30152.4]
  assign x417_outr_UnitPipe_sm_io_ctrDone = x417_outr_UnitPipe_sm_io_ctrInc & _T_357; // @[sm_x418_outr_UnitPipe.scala 78:40:@30132.4]
  assign x417_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@30179.4]
  assign x417_outr_UnitPipe_sm_io_doneIn_0 = x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@30149.4]
  assign RetimeWrapper_3_clock = clock; // @[:@30158.4]
  assign RetimeWrapper_3_reset = reset; // @[:@30159.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@30161.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@30160.4]
  assign RetimeWrapper_4_clock = clock; // @[:@30166.4]
  assign RetimeWrapper_4_reset = reset; // @[:@30167.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@30169.4]
  assign RetimeWrapper_4_io_in = x417_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@30168.4]
  assign x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_clock = clock; // @[:@30196.4]
  assign x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_reset = reset; // @[:@30197.4]
  assign x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x279_TREADY = io_in_x279_TREADY; // @[sm_x417_outr_UnitPipe.scala 48:23:@30251.4]
  assign x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x278_TVALID = io_in_x278_TVALID; // @[sm_x417_outr_UnitPipe.scala 49:23:@30261.4]
  assign x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x278_TDATA = io_in_x278_TDATA; // @[sm_x417_outr_UnitPipe.scala 49:23:@30259.4]
  assign x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x278_TID = io_in_x278_TID; // @[sm_x417_outr_UnitPipe.scala 49:23:@30255.4]
  assign x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_in_x278_TDEST = io_in_x278_TDEST; // @[sm_x417_outr_UnitPipe.scala 49:23:@30254.4]
  assign x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x417_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x417_outr_UnitPipe.scala 81:22:@30270.4]
  assign x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x417_outr_UnitPipe_sm_io_childAck_0; // @[sm_x417_outr_UnitPipe.scala 81:22:@30268.4]
  assign x417_outr_UnitPipe_kernelx417_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x417_outr_UnitPipe.scala 80:18:@30262.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_357 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_357 <= 1'h0;
    end else begin
      _T_357 <= _T_354;
    end
  end
endmodule
module x440_outr_UnitPipe_sm( // @[:@30759.2]
  input   clock, // @[:@30760.4]
  input   reset, // @[:@30761.4]
  input   io_enable, // @[:@30762.4]
  output  io_done, // @[:@30762.4]
  input   io_parentAck, // @[:@30762.4]
  input   io_doneIn_0, // @[:@30762.4]
  input   io_doneIn_1, // @[:@30762.4]
  input   io_doneIn_2, // @[:@30762.4]
  output  io_enableOut_0, // @[:@30762.4]
  output  io_enableOut_1, // @[:@30762.4]
  output  io_enableOut_2, // @[:@30762.4]
  output  io_childAck_0, // @[:@30762.4]
  output  io_childAck_1, // @[:@30762.4]
  output  io_childAck_2, // @[:@30762.4]
  input   io_ctrCopyDone_0, // @[:@30762.4]
  input   io_ctrCopyDone_1, // @[:@30762.4]
  input   io_ctrCopyDone_2 // @[:@30762.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@30765.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@30765.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@30765.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@30765.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@30765.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@30765.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@30768.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@30768.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@30768.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@30768.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@30768.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@30768.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@30771.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@30771.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@30771.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@30771.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@30771.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@30771.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@30774.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@30774.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@30774.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@30774.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@30774.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@30774.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@30777.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@30777.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@30777.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@30777.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@30777.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@30777.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@30780.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@30780.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@30780.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@30780.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@30780.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@30780.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@30821.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@30821.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@30821.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@30821.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@30821.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@30821.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@30824.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@30824.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@30824.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@30824.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@30824.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@30824.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@30827.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@30827.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@30827.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@30827.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@30827.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@30827.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@30878.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@30878.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@30878.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@30878.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@30878.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@30892.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@30892.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@30892.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@30892.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@30892.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@30910.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@30910.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@30910.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@30910.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@30910.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@30947.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@30947.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@30947.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@30947.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@30947.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@30961.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@30961.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@30961.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@30961.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@30961.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@30979.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@30979.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@30979.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@30979.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@30979.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@31016.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@31016.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@31016.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@31016.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@31016.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@31030.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@31030.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@31030.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@31030.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@31030.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@31048.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@31048.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@31048.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@31048.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@31048.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@31105.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@31105.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@31105.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@31105.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@31105.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@31122.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@31122.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@31122.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@31122.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@31122.4]
  wire  _T_77; // @[Controllers.scala 80:47:@30783.4]
  wire  allDone; // @[Controllers.scala 80:47:@30784.4]
  wire  _T_151; // @[Controllers.scala 165:35:@30862.4]
  wire  _T_153; // @[Controllers.scala 165:60:@30863.4]
  wire  _T_154; // @[Controllers.scala 165:58:@30864.4]
  wire  _T_156; // @[Controllers.scala 165:76:@30865.4]
  wire  _T_157; // @[Controllers.scala 165:74:@30866.4]
  wire  _T_161; // @[Controllers.scala 165:109:@30869.4]
  wire  _T_164; // @[Controllers.scala 165:141:@30871.4]
  wire  _T_172; // @[package.scala 96:25:@30883.4 package.scala 96:25:@30884.4]
  wire  _T_176; // @[Controllers.scala 167:54:@30886.4]
  wire  _T_177; // @[Controllers.scala 167:52:@30887.4]
  wire  _T_184; // @[package.scala 96:25:@30897.4 package.scala 96:25:@30898.4]
  wire  _T_202; // @[package.scala 96:25:@30915.4 package.scala 96:25:@30916.4]
  wire  _T_206; // @[Controllers.scala 169:67:@30918.4]
  wire  _T_207; // @[Controllers.scala 169:86:@30919.4]
  wire  _T_219; // @[Controllers.scala 165:35:@30931.4]
  wire  _T_221; // @[Controllers.scala 165:60:@30932.4]
  wire  _T_222; // @[Controllers.scala 165:58:@30933.4]
  wire  _T_224; // @[Controllers.scala 165:76:@30934.4]
  wire  _T_225; // @[Controllers.scala 165:74:@30935.4]
  wire  _T_229; // @[Controllers.scala 165:109:@30938.4]
  wire  _T_232; // @[Controllers.scala 165:141:@30940.4]
  wire  _T_240; // @[package.scala 96:25:@30952.4 package.scala 96:25:@30953.4]
  wire  _T_244; // @[Controllers.scala 167:54:@30955.4]
  wire  _T_245; // @[Controllers.scala 167:52:@30956.4]
  wire  _T_252; // @[package.scala 96:25:@30966.4 package.scala 96:25:@30967.4]
  wire  _T_270; // @[package.scala 96:25:@30984.4 package.scala 96:25:@30985.4]
  wire  _T_274; // @[Controllers.scala 169:67:@30987.4]
  wire  _T_275; // @[Controllers.scala 169:86:@30988.4]
  wire  _T_287; // @[Controllers.scala 165:35:@31000.4]
  wire  _T_289; // @[Controllers.scala 165:60:@31001.4]
  wire  _T_290; // @[Controllers.scala 165:58:@31002.4]
  wire  _T_292; // @[Controllers.scala 165:76:@31003.4]
  wire  _T_293; // @[Controllers.scala 165:74:@31004.4]
  wire  _T_297; // @[Controllers.scala 165:109:@31007.4]
  wire  _T_300; // @[Controllers.scala 165:141:@31009.4]
  wire  _T_308; // @[package.scala 96:25:@31021.4 package.scala 96:25:@31022.4]
  wire  _T_312; // @[Controllers.scala 167:54:@31024.4]
  wire  _T_313; // @[Controllers.scala 167:52:@31025.4]
  wire  _T_320; // @[package.scala 96:25:@31035.4 package.scala 96:25:@31036.4]
  wire  _T_338; // @[package.scala 96:25:@31053.4 package.scala 96:25:@31054.4]
  wire  _T_342; // @[Controllers.scala 169:67:@31056.4]
  wire  _T_343; // @[Controllers.scala 169:86:@31057.4]
  wire  _T_358; // @[Controllers.scala 213:68:@31075.4]
  wire  _T_360; // @[Controllers.scala 213:90:@31077.4]
  wire  _T_362; // @[Controllers.scala 213:132:@31079.4]
  wire  _T_366; // @[Controllers.scala 213:68:@31084.4]
  wire  _T_368; // @[Controllers.scala 213:90:@31086.4]
  wire  _T_374; // @[Controllers.scala 213:68:@31092.4]
  wire  _T_376; // @[Controllers.scala 213:90:@31094.4]
  wire  _T_383; // @[package.scala 100:49:@31100.4]
  reg  _T_386; // @[package.scala 48:56:@31101.4]
  reg [31:0] _RAND_0;
  wire  _T_387; // @[package.scala 100:41:@31103.4]
  reg  _T_400; // @[package.scala 48:56:@31119.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@30765.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@30768.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@30771.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@30774.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@30777.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@30780.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@30821.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@30824.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@30827.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@30878.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@30892.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@30910.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@30947.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@30961.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@30979.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@31016.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@31030.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@31048.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@31105.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@31122.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@30783.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@30784.4]
  assign _T_151 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@30862.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@30863.4]
  assign _T_154 = _T_151 & _T_153; // @[Controllers.scala 165:58:@30864.4]
  assign _T_156 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@30865.4]
  assign _T_157 = _T_154 & _T_156; // @[Controllers.scala 165:74:@30866.4]
  assign _T_161 = _T_157 & io_enable; // @[Controllers.scala 165:109:@30869.4]
  assign _T_164 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@30871.4]
  assign _T_172 = RetimeWrapper_io_out; // @[package.scala 96:25:@30883.4 package.scala 96:25:@30884.4]
  assign _T_176 = _T_172 == 1'h0; // @[Controllers.scala 167:54:@30886.4]
  assign _T_177 = io_doneIn_0 | _T_176; // @[Controllers.scala 167:52:@30887.4]
  assign _T_184 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@30897.4 package.scala 96:25:@30898.4]
  assign _T_202 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@30915.4 package.scala 96:25:@30916.4]
  assign _T_206 = _T_202 == 1'h0; // @[Controllers.scala 169:67:@30918.4]
  assign _T_207 = _T_206 & io_enable; // @[Controllers.scala 169:86:@30919.4]
  assign _T_219 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@30931.4]
  assign _T_221 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@30932.4]
  assign _T_222 = _T_219 & _T_221; // @[Controllers.scala 165:58:@30933.4]
  assign _T_224 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@30934.4]
  assign _T_225 = _T_222 & _T_224; // @[Controllers.scala 165:74:@30935.4]
  assign _T_229 = _T_225 & io_enable; // @[Controllers.scala 165:109:@30938.4]
  assign _T_232 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@30940.4]
  assign _T_240 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@30952.4 package.scala 96:25:@30953.4]
  assign _T_244 = _T_240 == 1'h0; // @[Controllers.scala 167:54:@30955.4]
  assign _T_245 = io_doneIn_1 | _T_244; // @[Controllers.scala 167:52:@30956.4]
  assign _T_252 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@30966.4 package.scala 96:25:@30967.4]
  assign _T_270 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@30984.4 package.scala 96:25:@30985.4]
  assign _T_274 = _T_270 == 1'h0; // @[Controllers.scala 169:67:@30987.4]
  assign _T_275 = _T_274 & io_enable; // @[Controllers.scala 169:86:@30988.4]
  assign _T_287 = ~ iterDone_2_io_output; // @[Controllers.scala 165:35:@31000.4]
  assign _T_289 = io_doneIn_2 == 1'h0; // @[Controllers.scala 165:60:@31001.4]
  assign _T_290 = _T_287 & _T_289; // @[Controllers.scala 165:58:@31002.4]
  assign _T_292 = done_2_io_output == 1'h0; // @[Controllers.scala 165:76:@31003.4]
  assign _T_293 = _T_290 & _T_292; // @[Controllers.scala 165:74:@31004.4]
  assign _T_297 = _T_293 & io_enable; // @[Controllers.scala 165:109:@31007.4]
  assign _T_300 = io_ctrCopyDone_2 == 1'h0; // @[Controllers.scala 165:141:@31009.4]
  assign _T_308 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@31021.4 package.scala 96:25:@31022.4]
  assign _T_312 = _T_308 == 1'h0; // @[Controllers.scala 167:54:@31024.4]
  assign _T_313 = io_doneIn_2 | _T_312; // @[Controllers.scala 167:52:@31025.4]
  assign _T_320 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@31035.4 package.scala 96:25:@31036.4]
  assign _T_338 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@31053.4 package.scala 96:25:@31054.4]
  assign _T_342 = _T_338 == 1'h0; // @[Controllers.scala 169:67:@31056.4]
  assign _T_343 = _T_342 & io_enable; // @[Controllers.scala 169:86:@31057.4]
  assign _T_358 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@31075.4]
  assign _T_360 = _T_358 & _T_151; // @[Controllers.scala 213:90:@31077.4]
  assign _T_362 = ~ allDone; // @[Controllers.scala 213:132:@31079.4]
  assign _T_366 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@31084.4]
  assign _T_368 = _T_366 & _T_219; // @[Controllers.scala 213:90:@31086.4]
  assign _T_374 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@31092.4]
  assign _T_376 = _T_374 & _T_287; // @[Controllers.scala 213:90:@31094.4]
  assign _T_383 = allDone == 1'h0; // @[package.scala 100:49:@31100.4]
  assign _T_387 = allDone & _T_386; // @[package.scala 100:41:@31103.4]
  assign io_done = RetimeWrapper_10_io_out; // @[Controllers.scala 245:13:@31129.4]
  assign io_enableOut_0 = _T_360 & _T_362; // @[Controllers.scala 213:55:@31083.4]
  assign io_enableOut_1 = _T_368 & _T_362; // @[Controllers.scala 213:55:@31091.4]
  assign io_enableOut_2 = _T_376 & _T_362; // @[Controllers.scala 213:55:@31099.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@31070.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@31072.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@31074.4]
  assign active_0_clock = clock; // @[:@30766.4]
  assign active_0_reset = reset; // @[:@30767.4]
  assign active_0_io_input_set = _T_161 & _T_164; // @[Controllers.scala 165:32:@30873.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@30877.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@30787.4]
  assign active_1_clock = clock; // @[:@30769.4]
  assign active_1_reset = reset; // @[:@30770.4]
  assign active_1_io_input_set = _T_229 & _T_232; // @[Controllers.scala 165:32:@30942.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@30946.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@30788.4]
  assign active_2_clock = clock; // @[:@30772.4]
  assign active_2_reset = reset; // @[:@30773.4]
  assign active_2_io_input_set = _T_297 & _T_300; // @[Controllers.scala 165:32:@31011.4]
  assign active_2_io_input_reset = io_ctrCopyDone_2 | io_parentAck; // @[Controllers.scala 166:34:@31015.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@30789.4]
  assign done_0_clock = clock; // @[:@30775.4]
  assign done_0_reset = reset; // @[:@30776.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_207; // @[Controllers.scala 169:30:@30923.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@30801.4 Controllers.scala 170:32:@30930.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@30790.4]
  assign done_1_clock = clock; // @[:@30778.4]
  assign done_1_reset = reset; // @[:@30779.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_275; // @[Controllers.scala 169:30:@30992.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@30810.4 Controllers.scala 170:32:@30999.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@30791.4]
  assign done_2_clock = clock; // @[:@30781.4]
  assign done_2_reset = reset; // @[:@30782.4]
  assign done_2_io_input_set = io_ctrCopyDone_2 | _T_343; // @[Controllers.scala 169:30:@31061.4]
  assign done_2_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@30819.4 Controllers.scala 170:32:@31068.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@30792.4]
  assign iterDone_0_clock = clock; // @[:@30822.4]
  assign iterDone_0_reset = reset; // @[:@30823.4]
  assign iterDone_0_io_input_set = _T_177 & io_enable; // @[Controllers.scala 167:34:@30891.4]
  assign iterDone_0_io_input_reset = _T_184 | io_parentAck; // @[Controllers.scala 92:37:@30841.4 Controllers.scala 168:36:@30907.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@30830.4]
  assign iterDone_1_clock = clock; // @[:@30825.4]
  assign iterDone_1_reset = reset; // @[:@30826.4]
  assign iterDone_1_io_input_set = _T_245 & io_enable; // @[Controllers.scala 167:34:@30960.4]
  assign iterDone_1_io_input_reset = _T_252 | io_parentAck; // @[Controllers.scala 92:37:@30850.4 Controllers.scala 168:36:@30976.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@30831.4]
  assign iterDone_2_clock = clock; // @[:@30828.4]
  assign iterDone_2_reset = reset; // @[:@30829.4]
  assign iterDone_2_io_input_set = _T_313 & io_enable; // @[Controllers.scala 167:34:@31029.4]
  assign iterDone_2_io_input_reset = _T_320 | io_parentAck; // @[Controllers.scala 92:37:@30859.4 Controllers.scala 168:36:@31045.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@30832.4]
  assign RetimeWrapper_clock = clock; // @[:@30879.4]
  assign RetimeWrapper_reset = reset; // @[:@30880.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@30882.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@30881.4]
  assign RetimeWrapper_1_clock = clock; // @[:@30893.4]
  assign RetimeWrapper_1_reset = reset; // @[:@30894.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@30896.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@30895.4]
  assign RetimeWrapper_2_clock = clock; // @[:@30911.4]
  assign RetimeWrapper_2_reset = reset; // @[:@30912.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@30914.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@30913.4]
  assign RetimeWrapper_3_clock = clock; // @[:@30948.4]
  assign RetimeWrapper_3_reset = reset; // @[:@30949.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@30951.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@30950.4]
  assign RetimeWrapper_4_clock = clock; // @[:@30962.4]
  assign RetimeWrapper_4_reset = reset; // @[:@30963.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@30965.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@30964.4]
  assign RetimeWrapper_5_clock = clock; // @[:@30980.4]
  assign RetimeWrapper_5_reset = reset; // @[:@30981.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@30983.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@30982.4]
  assign RetimeWrapper_6_clock = clock; // @[:@31017.4]
  assign RetimeWrapper_6_reset = reset; // @[:@31018.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@31020.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@31019.4]
  assign RetimeWrapper_7_clock = clock; // @[:@31031.4]
  assign RetimeWrapper_7_reset = reset; // @[:@31032.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@31034.4]
  assign RetimeWrapper_7_io_in = io_doneIn_2; // @[package.scala 94:16:@31033.4]
  assign RetimeWrapper_8_clock = clock; // @[:@31049.4]
  assign RetimeWrapper_8_reset = reset; // @[:@31050.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@31052.4]
  assign RetimeWrapper_8_io_in = 1'h1; // @[package.scala 94:16:@31051.4]
  assign RetimeWrapper_9_clock = clock; // @[:@31106.4]
  assign RetimeWrapper_9_reset = reset; // @[:@31107.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@31109.4]
  assign RetimeWrapper_9_io_in = _T_387 | io_parentAck; // @[package.scala 94:16:@31108.4]
  assign RetimeWrapper_10_clock = clock; // @[:@31123.4]
  assign RetimeWrapper_10_reset = reset; // @[:@31124.4]
  assign RetimeWrapper_10_io_flow = io_enable; // @[package.scala 95:18:@31126.4]
  assign RetimeWrapper_10_io_in = allDone & _T_400; // @[package.scala 94:16:@31125.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_386 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_400 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_386 <= 1'h0;
    end else begin
      _T_386 <= _T_383;
    end
    if (reset) begin
      _T_400 <= 1'h0;
    end else begin
      _T_400 <= _T_383;
    end
  end
endmodule
module x426_inr_UnitPipe_sm( // @[:@31302.2]
  input   clock, // @[:@31303.4]
  input   reset, // @[:@31304.4]
  input   io_enable, // @[:@31305.4]
  output  io_done, // @[:@31305.4]
  output  io_doneLatch, // @[:@31305.4]
  input   io_ctrDone, // @[:@31305.4]
  output  io_datapathEn, // @[:@31305.4]
  output  io_ctrInc, // @[:@31305.4]
  input   io_parentAck, // @[:@31305.4]
  input   io_backpressure // @[:@31305.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@31307.4]
  wire  active_reset; // @[Controllers.scala 261:22:@31307.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@31307.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@31307.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@31307.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@31307.4]
  wire  done_clock; // @[Controllers.scala 262:20:@31310.4]
  wire  done_reset; // @[Controllers.scala 262:20:@31310.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@31310.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@31310.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@31310.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@31310.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@31364.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@31364.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@31364.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@31364.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@31364.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@31372.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@31372.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@31372.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@31372.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@31372.4]
  wire  _T_80; // @[Controllers.scala 264:48:@31315.4]
  wire  _T_81; // @[Controllers.scala 264:46:@31316.4]
  wire  _T_82; // @[Controllers.scala 264:62:@31317.4]
  wire  _T_83; // @[Controllers.scala 264:60:@31318.4]
  wire  _T_100; // @[package.scala 100:49:@31335.4]
  reg  _T_103; // @[package.scala 48:56:@31336.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 100:49:@31344.4]
  wire  _T_116; // @[Controllers.scala 283:41:@31352.4]
  wire  _T_117; // @[Controllers.scala 283:59:@31353.4]
  wire  _T_119; // @[Controllers.scala 284:37:@31356.4]
  reg  _T_125; // @[package.scala 48:56:@31360.4]
  reg [31:0] _RAND_1;
  reg  _T_142; // @[Controllers.scala 291:31:@31382.4]
  reg [31:0] _RAND_2;
  reg  _T_149; // @[package.scala 48:56:@31385.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:41:@31387.4]
  wire  _T_152; // @[Controllers.scala 292:61:@31388.4]
  wire  _T_153; // @[Controllers.scala 292:24:@31389.4]
  SRFF active ( // @[Controllers.scala 261:22:@31307.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@31310.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@31364.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@31372.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@31315.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@31316.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@31317.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@31318.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@31335.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 100:49:@31344.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@31352.4]
  assign _T_117 = _T_116 & io_enable; // @[Controllers.scala 283:59:@31353.4]
  assign _T_119 = active_io_output & io_enable; // @[Controllers.scala 284:37:@31356.4]
  assign _T_150 = done_io_output & _T_149; // @[package.scala 100:41:@31387.4]
  assign _T_152 = _T_150 ? 1'h1 : _T_142; // @[Controllers.scala 292:61:@31388.4]
  assign _T_153 = io_parentAck ? 1'h0 : _T_152; // @[Controllers.scala 292:24:@31389.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@31363.4]
  assign io_doneLatch = _T_142; // @[Controllers.scala 293:18:@31391.4]
  assign io_datapathEn = _T_117 & io_backpressure; // @[Controllers.scala 283:21:@31355.4]
  assign io_ctrInc = _T_119 & io_backpressure; // @[Controllers.scala 284:17:@31358.4]
  assign active_clock = clock; // @[:@31308.4]
  assign active_reset = reset; // @[:@31309.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@31320.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@31324.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@31325.4]
  assign done_clock = clock; // @[:@31311.4]
  assign done_reset = reset; // @[:@31312.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@31340.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@31333.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@31334.4]
  assign RetimeWrapper_clock = clock; // @[:@31365.4]
  assign RetimeWrapper_reset = reset; // @[:@31366.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@31368.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@31367.4]
  assign RetimeWrapper_1_clock = clock; // @[:@31373.4]
  assign RetimeWrapper_1_reset = reset; // @[:@31374.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@31376.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 94:16:@31375.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_125 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_142 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_149 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_142 <= 1'h0;
      end else begin
        if (_T_150) begin
          _T_142 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_108;
    end
  end
endmodule
module x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1( // @[:@31466.2]
  input  [63:0] io_in_x276_outdram_number, // @[:@31469.4]
  output        io_in_x419_valid, // @[:@31469.4]
  output [63:0] io_in_x419_bits_addr, // @[:@31469.4]
  output [31:0] io_in_x419_bits_size, // @[:@31469.4]
  input         io_sigsIn_backpressure, // @[:@31469.4]
  input         io_sigsIn_datapathEn, // @[:@31469.4]
  input         io_rr // @[:@31469.4]
);
  wire [96:0] x423_tuple; // @[Cat.scala 30:58:@31483.4]
  wire  _T_135; // @[implicits.scala 55:10:@31486.4]
  assign x423_tuple = {33'h1fa400,io_in_x276_outdram_number}; // @[Cat.scala 30:58:@31483.4]
  assign _T_135 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@31486.4]
  assign io_in_x419_valid = _T_135 & io_sigsIn_backpressure; // @[sm_x426_inr_UnitPipe.scala 65:18:@31489.4]
  assign io_in_x419_bits_addr = x423_tuple[63:0]; // @[sm_x426_inr_UnitPipe.scala 66:22:@31491.4]
  assign io_in_x419_bits_size = x423_tuple[95:64]; // @[sm_x426_inr_UnitPipe.scala 67:22:@31493.4]
endmodule
module FF_13( // @[:@31495.2]
  input         clock, // @[:@31496.4]
  input         reset, // @[:@31497.4]
  output [22:0] io_rPort_0_output_0, // @[:@31498.4]
  input  [22:0] io_wPort_0_data_0, // @[:@31498.4]
  input         io_wPort_0_reset, // @[:@31498.4]
  input         io_wPort_0_en_0 // @[:@31498.4]
);
  reg [22:0] ff; // @[MemPrimitives.scala 311:19:@31513.4]
  reg [31:0] _RAND_0;
  wire [22:0] _T_68; // @[MemPrimitives.scala 315:32:@31515.4]
  wire [22:0] _T_69; // @[MemPrimitives.scala 315:12:@31516.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 315:32:@31515.4]
  assign _T_69 = io_wPort_0_reset ? 23'h0 : _T_68; // @[MemPrimitives.scala 315:12:@31516.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 316:34:@31518.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[22:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 23'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 23'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_5( // @[:@31533.2]
  input         clock, // @[:@31534.4]
  input         reset, // @[:@31535.4]
  input         io_input_reset, // @[:@31536.4]
  input         io_input_enable, // @[:@31536.4]
  output [22:0] io_output_count_0, // @[:@31536.4]
  output        io_output_oobs_0, // @[:@31536.4]
  output        io_output_done // @[:@31536.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@31549.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@31549.4]
  wire [22:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@31549.4]
  wire [22:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@31549.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@31549.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@31549.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@31565.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@31565.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@31565.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@31565.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@31565.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@31565.4]
  wire  _T_36; // @[Counter.scala 264:45:@31568.4]
  wire [22:0] _T_48; // @[Counter.scala 287:52:@31593.4]
  wire [23:0] _T_50; // @[Counter.scala 291:33:@31594.4]
  wire [22:0] _T_51; // @[Counter.scala 291:33:@31595.4]
  wire [22:0] _T_52; // @[Counter.scala 291:33:@31596.4]
  wire  _T_57; // @[Counter.scala 293:18:@31598.4]
  wire [22:0] _T_68; // @[Counter.scala 299:115:@31606.4]
  wire [22:0] _T_71; // @[Counter.scala 299:152:@31609.4]
  wire [22:0] _T_72; // @[Counter.scala 299:74:@31610.4]
  wire  _T_75; // @[Counter.scala 322:102:@31614.4]
  wire  _T_77; // @[Counter.scala 322:130:@31615.4]
  FF_13 bases_0 ( // @[Counter.scala 261:53:@31549.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@31565.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@31568.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@31593.4]
  assign _T_50 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@31594.4]
  assign _T_51 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@31595.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@31596.4]
  assign _T_57 = $signed(_T_52) >= $signed(23'sh1fa400); // @[Counter.scala 293:18:@31598.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@31606.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@31609.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@31610.4]
  assign _T_75 = $signed(_T_48) < $signed(23'sh0); // @[Counter.scala 322:102:@31614.4]
  assign _T_77 = $signed(_T_48) >= $signed(23'sh1fa400); // @[Counter.scala 322:130:@31615.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@31613.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@31617.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@31619.4]
  assign bases_0_clock = clock; // @[:@31550.4]
  assign bases_0_reset = reset; // @[:@31551.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 23'h0 : _T_72; // @[Counter.scala 299:31:@31612.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@31591.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@31592.4]
  assign SRFF_clock = clock; // @[:@31566.4]
  assign SRFF_reset = reset; // @[:@31567.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@31570.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@31572.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@31573.4]
endmodule
module x428_ctrchain( // @[:@31624.2]
  input         clock, // @[:@31625.4]
  input         reset, // @[:@31626.4]
  input         io_input_reset, // @[:@31627.4]
  input         io_input_enable, // @[:@31627.4]
  output [22:0] io_output_counts_0, // @[:@31627.4]
  output        io_output_oobs_0, // @[:@31627.4]
  output        io_output_done // @[:@31627.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@31629.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@31629.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@31629.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@31629.4]
  wire [22:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@31629.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@31629.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@31629.4]
  reg  wasDone; // @[Counter.scala 542:24:@31638.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 546:69:@31644.4]
  wire  _T_47; // @[Counter.scala 546:80:@31645.4]
  reg  doneLatch; // @[Counter.scala 550:26:@31650.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 551:48:@31651.4]
  wire  _T_55; // @[Counter.scala 551:19:@31652.4]
  SingleCounter_5 ctrs_0 ( // @[Counter.scala 513:46:@31629.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 546:69:@31644.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 546:80:@31645.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@31651.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 551:19:@31652.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@31654.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@31656.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 546:18:@31647.4]
  assign ctrs_0_clock = clock; // @[:@31630.4]
  assign ctrs_0_reset = reset; // @[:@31631.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@31635.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@31636.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x435_inr_Foreach_sm( // @[:@31844.2]
  input   clock, // @[:@31845.4]
  input   reset, // @[:@31846.4]
  input   io_enable, // @[:@31847.4]
  output  io_done, // @[:@31847.4]
  output  io_doneLatch, // @[:@31847.4]
  input   io_ctrDone, // @[:@31847.4]
  output  io_datapathEn, // @[:@31847.4]
  output  io_ctrInc, // @[:@31847.4]
  output  io_ctrRst, // @[:@31847.4]
  input   io_parentAck, // @[:@31847.4]
  input   io_backpressure, // @[:@31847.4]
  input   io_break // @[:@31847.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@31849.4]
  wire  active_reset; // @[Controllers.scala 261:22:@31849.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@31849.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@31849.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@31849.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@31849.4]
  wire  done_clock; // @[Controllers.scala 262:20:@31852.4]
  wire  done_reset; // @[Controllers.scala 262:20:@31852.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@31852.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@31852.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@31852.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@31852.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@31886.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@31886.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@31886.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@31886.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@31886.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@31908.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@31908.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@31908.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@31908.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@31908.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@31920.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@31920.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@31920.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@31920.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@31920.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@31928.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@31928.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@31928.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@31928.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@31928.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@31944.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@31944.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@31944.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@31944.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@31944.4]
  wire  _T_80; // @[Controllers.scala 264:48:@31857.4]
  wire  _T_81; // @[Controllers.scala 264:46:@31858.4]
  wire  _T_82; // @[Controllers.scala 264:62:@31859.4]
  wire  _T_83; // @[Controllers.scala 264:60:@31860.4]
  wire  _T_100; // @[package.scala 100:49:@31877.4]
  reg  _T_103; // @[package.scala 48:56:@31878.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@31891.4 package.scala 96:25:@31892.4]
  wire  _T_110; // @[package.scala 100:49:@31893.4]
  reg  _T_113; // @[package.scala 48:56:@31894.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@31896.4]
  wire  _T_118; // @[Controllers.scala 283:41:@31901.4]
  wire  _T_119; // @[Controllers.scala 283:59:@31902.4]
  wire  _T_121; // @[Controllers.scala 284:37:@31905.4]
  wire  _T_124; // @[package.scala 96:25:@31913.4 package.scala 96:25:@31914.4]
  wire  _T_126; // @[package.scala 100:49:@31915.4]
  reg  _T_129; // @[package.scala 48:56:@31916.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@31938.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@31940.4]
  reg  _T_153; // @[package.scala 48:56:@31941.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@31949.4 package.scala 96:25:@31950.4]
  wire  _T_158; // @[Controllers.scala 292:61:@31951.4]
  wire  _T_159; // @[Controllers.scala 292:24:@31952.4]
  SRFF active ( // @[Controllers.scala 261:22:@31849.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@31852.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@31886.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@31908.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@31920.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@31928.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@31944.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@31857.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@31858.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@31859.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@31860.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@31877.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@31891.4 package.scala 96:25:@31892.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@31893.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@31896.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@31901.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@31902.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@31905.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@31913.4 package.scala 96:25:@31914.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@31915.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@31940.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@31949.4 package.scala 96:25:@31950.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@31951.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@31952.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@31919.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@31954.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@31904.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@31907.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@31899.4]
  assign active_clock = clock; // @[:@31850.4]
  assign active_reset = reset; // @[:@31851.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@31862.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@31866.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@31867.4]
  assign done_clock = clock; // @[:@31853.4]
  assign done_reset = reset; // @[:@31854.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@31882.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@31875.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@31876.4]
  assign RetimeWrapper_clock = clock; // @[:@31887.4]
  assign RetimeWrapper_reset = reset; // @[:@31888.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@31890.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@31889.4]
  assign RetimeWrapper_1_clock = clock; // @[:@31909.4]
  assign RetimeWrapper_1_reset = reset; // @[:@31910.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@31912.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@31911.4]
  assign RetimeWrapper_2_clock = clock; // @[:@31921.4]
  assign RetimeWrapper_2_reset = reset; // @[:@31922.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@31924.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@31923.4]
  assign RetimeWrapper_3_clock = clock; // @[:@31929.4]
  assign RetimeWrapper_3_reset = reset; // @[:@31930.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@31932.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@31931.4]
  assign RetimeWrapper_4_clock = clock; // @[:@31945.4]
  assign RetimeWrapper_4_reset = reset; // @[:@31946.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@31948.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@31947.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x435_inr_Foreach_kernelx435_inr_Foreach_concrete1( // @[:@32166.2]
  input         clock, // @[:@32167.4]
  input         reset, // @[:@32168.4]
  output [20:0] io_in_x280_outbuf_0_rPort_0_ofs_0, // @[:@32169.4]
  output        io_in_x280_outbuf_0_rPort_0_en_0, // @[:@32169.4]
  output        io_in_x280_outbuf_0_rPort_0_backpressure, // @[:@32169.4]
  input  [7:0]  io_in_x280_outbuf_0_rPort_0_output_0, // @[:@32169.4]
  output        io_in_x420_valid, // @[:@32169.4]
  output [7:0]  io_in_x420_bits_wdata_0, // @[:@32169.4]
  output        io_in_x420_bits_wstrb, // @[:@32169.4]
  input         io_sigsIn_backpressure, // @[:@32169.4]
  input         io_sigsIn_datapathEn, // @[:@32169.4]
  input         io_sigsIn_break, // @[:@32169.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@32169.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@32169.4]
  input         io_rr // @[:@32169.4]
);
  wire [31:0] __io_b; // @[Math.scala 709:24:@32196.4]
  wire [31:0] __io_result; // @[Math.scala 709:24:@32196.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@32225.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@32225.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@32225.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@32225.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@32225.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32234.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32234.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32234.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@32234.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@32234.4]
  wire  b430; // @[sm_x435_inr_Foreach.scala 62:18:@32204.4]
  wire  _T_274; // @[sm_x435_inr_Foreach.scala 67:129:@32208.4]
  wire  _T_278; // @[implicits.scala 55:10:@32211.4]
  wire  _T_279; // @[sm_x435_inr_Foreach.scala 67:146:@32212.4]
  wire [8:0] x433_tuple; // @[Cat.scala 30:58:@32222.4]
  wire  _T_290; // @[package.scala 96:25:@32239.4 package.scala 96:25:@32240.4]
  wire  _T_292; // @[implicits.scala 55:10:@32241.4]
  wire  x615_b430_D2; // @[package.scala 96:25:@32230.4 package.scala 96:25:@32231.4]
  wire  _T_293; // @[sm_x435_inr_Foreach.scala 74:112:@32242.4]
  wire [31:0] b429_number; // @[Math.scala 712:22:@32201.4 Math.scala 713:14:@32202.4]
  _ _ ( // @[Math.scala 709:24:@32196.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@32225.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@32234.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign b430 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x435_inr_Foreach.scala 62:18:@32204.4]
  assign _T_274 = ~ io_sigsIn_break; // @[sm_x435_inr_Foreach.scala 67:129:@32208.4]
  assign _T_278 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@32211.4]
  assign _T_279 = _T_274 & _T_278; // @[sm_x435_inr_Foreach.scala 67:146:@32212.4]
  assign x433_tuple = {1'h1,io_in_x280_outbuf_0_rPort_0_output_0}; // @[Cat.scala 30:58:@32222.4]
  assign _T_290 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@32239.4 package.scala 96:25:@32240.4]
  assign _T_292 = io_rr ? _T_290 : 1'h0; // @[implicits.scala 55:10:@32241.4]
  assign x615_b430_D2 = RetimeWrapper_io_out; // @[package.scala 96:25:@32230.4 package.scala 96:25:@32231.4]
  assign _T_293 = _T_292 & x615_b430_D2; // @[sm_x435_inr_Foreach.scala 74:112:@32242.4]
  assign b429_number = __io_result; // @[Math.scala 712:22:@32201.4 Math.scala 713:14:@32202.4]
  assign io_in_x280_outbuf_0_rPort_0_ofs_0 = b429_number[20:0]; // @[MemInterfaceType.scala 107:54:@32215.4]
  assign io_in_x280_outbuf_0_rPort_0_en_0 = _T_279 & b430; // @[MemInterfaceType.scala 110:79:@32217.4]
  assign io_in_x280_outbuf_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@32216.4]
  assign io_in_x420_valid = _T_293 & io_sigsIn_backpressure; // @[sm_x435_inr_Foreach.scala 74:18:@32244.4]
  assign io_in_x420_bits_wdata_0 = x433_tuple[7:0]; // @[sm_x435_inr_Foreach.scala 75:26:@32246.4]
  assign io_in_x420_bits_wstrb = x433_tuple[8]; // @[sm_x435_inr_Foreach.scala 76:23:@32248.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 710:17:@32199.4]
  assign RetimeWrapper_clock = clock; // @[:@32226.4]
  assign RetimeWrapper_reset = reset; // @[:@32227.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32229.4]
  assign RetimeWrapper_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@32228.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32235.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32236.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@32238.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@32237.4]
endmodule
module x439_inr_UnitPipe_sm( // @[:@32404.2]
  input   clock, // @[:@32405.4]
  input   reset, // @[:@32406.4]
  input   io_enable, // @[:@32407.4]
  output  io_done, // @[:@32407.4]
  output  io_doneLatch, // @[:@32407.4]
  input   io_ctrDone, // @[:@32407.4]
  output  io_datapathEn, // @[:@32407.4]
  output  io_ctrInc, // @[:@32407.4]
  input   io_parentAck // @[:@32407.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@32409.4]
  wire  active_reset; // @[Controllers.scala 261:22:@32409.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@32409.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@32409.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@32409.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@32409.4]
  wire  done_clock; // @[Controllers.scala 262:20:@32412.4]
  wire  done_reset; // @[Controllers.scala 262:20:@32412.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@32412.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@32412.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@32412.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@32412.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@32446.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@32446.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@32446.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@32446.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@32446.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32468.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32468.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32468.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@32468.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@32468.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@32480.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@32480.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@32480.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@32480.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@32480.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@32488.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@32488.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@32488.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@32488.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@32488.4]
  wire  _T_80; // @[Controllers.scala 264:48:@32417.4]
  wire  _T_81; // @[Controllers.scala 264:46:@32418.4]
  wire  _T_82; // @[Controllers.scala 264:62:@32419.4]
  wire  _T_100; // @[package.scala 100:49:@32437.4]
  reg  _T_103; // @[package.scala 48:56:@32438.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@32461.4]
  wire  _T_124; // @[package.scala 96:25:@32473.4 package.scala 96:25:@32474.4]
  wire  _T_126; // @[package.scala 100:49:@32475.4]
  reg  _T_129; // @[package.scala 48:56:@32476.4]
  reg [31:0] _RAND_1;
  reg  _T_146; // @[Controllers.scala 291:31:@32498.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@32500.4]
  reg  _T_153; // @[package.scala 48:56:@32501.4]
  reg [31:0] _RAND_3;
  wire  _T_154; // @[package.scala 100:41:@32503.4]
  wire  _T_156; // @[Controllers.scala 292:61:@32504.4]
  wire  _T_157; // @[Controllers.scala 292:24:@32505.4]
  SRFF active ( // @[Controllers.scala 261:22:@32409.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@32412.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@32446.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@32468.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@32480.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@32488.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@32417.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@32418.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@32419.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@32437.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@32461.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@32473.4 package.scala 96:25:@32474.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@32475.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@32500.4]
  assign _T_154 = done_io_output & _T_153; // @[package.scala 100:41:@32503.4]
  assign _T_156 = _T_154 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@32504.4]
  assign _T_157 = io_parentAck ? 1'h0 : _T_156; // @[Controllers.scala 292:24:@32505.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@32479.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@32507.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@32464.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@32467.4]
  assign active_clock = clock; // @[:@32410.4]
  assign active_reset = reset; // @[:@32411.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@32422.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@32426.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@32427.4]
  assign done_clock = clock; // @[:@32413.4]
  assign done_reset = reset; // @[:@32414.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@32442.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@32435.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@32436.4]
  assign RetimeWrapper_clock = clock; // @[:@32447.4]
  assign RetimeWrapper_reset = reset; // @[:@32448.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@32450.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@32449.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32469.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32470.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@32472.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@32471.4]
  assign RetimeWrapper_2_clock = clock; // @[:@32481.4]
  assign RetimeWrapper_2_reset = reset; // @[:@32482.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@32484.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@32483.4]
  assign RetimeWrapper_3_clock = clock; // @[:@32489.4]
  assign RetimeWrapper_3_reset = reset; // @[:@32490.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@32492.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@32491.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_154) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x439_inr_UnitPipe_kernelx439_inr_UnitPipe_concrete1( // @[:@32582.2]
  output  io_in_x421_ready, // @[:@32585.4]
  input   io_sigsIn_datapathEn // @[:@32585.4]
);
  assign io_in_x421_ready = io_sigsIn_datapathEn; // @[sm_x439_inr_UnitPipe.scala 57:18:@32597.4]
endmodule
module x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1( // @[:@32600.2]
  input         clock, // @[:@32601.4]
  input         reset, // @[:@32602.4]
  input  [63:0] io_in_x276_outdram_number, // @[:@32603.4]
  output        io_in_x421_ready, // @[:@32603.4]
  input         io_in_x421_valid, // @[:@32603.4]
  output [20:0] io_in_x280_outbuf_0_rPort_0_ofs_0, // @[:@32603.4]
  output        io_in_x280_outbuf_0_rPort_0_en_0, // @[:@32603.4]
  output        io_in_x280_outbuf_0_rPort_0_backpressure, // @[:@32603.4]
  input  [7:0]  io_in_x280_outbuf_0_rPort_0_output_0, // @[:@32603.4]
  input         io_in_x420_ready, // @[:@32603.4]
  output        io_in_x420_valid, // @[:@32603.4]
  output [7:0]  io_in_x420_bits_wdata_0, // @[:@32603.4]
  output        io_in_x420_bits_wstrb, // @[:@32603.4]
  input         io_in_x419_ready, // @[:@32603.4]
  output        io_in_x419_valid, // @[:@32603.4]
  output [63:0] io_in_x419_bits_addr, // @[:@32603.4]
  output [31:0] io_in_x419_bits_size, // @[:@32603.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@32603.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@32603.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@32603.4]
  input         io_sigsIn_smChildAcks_0, // @[:@32603.4]
  input         io_sigsIn_smChildAcks_1, // @[:@32603.4]
  input         io_sigsIn_smChildAcks_2, // @[:@32603.4]
  output        io_sigsOut_smDoneIn_0, // @[:@32603.4]
  output        io_sigsOut_smDoneIn_1, // @[:@32603.4]
  output        io_sigsOut_smDoneIn_2, // @[:@32603.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@32603.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@32603.4]
  output        io_sigsOut_smCtrCopyDone_2, // @[:@32603.4]
  input         io_rr // @[:@32603.4]
);
  wire  x426_inr_UnitPipe_sm_clock; // @[sm_x426_inr_UnitPipe.scala 33:18:@32670.4]
  wire  x426_inr_UnitPipe_sm_reset; // @[sm_x426_inr_UnitPipe.scala 33:18:@32670.4]
  wire  x426_inr_UnitPipe_sm_io_enable; // @[sm_x426_inr_UnitPipe.scala 33:18:@32670.4]
  wire  x426_inr_UnitPipe_sm_io_done; // @[sm_x426_inr_UnitPipe.scala 33:18:@32670.4]
  wire  x426_inr_UnitPipe_sm_io_doneLatch; // @[sm_x426_inr_UnitPipe.scala 33:18:@32670.4]
  wire  x426_inr_UnitPipe_sm_io_ctrDone; // @[sm_x426_inr_UnitPipe.scala 33:18:@32670.4]
  wire  x426_inr_UnitPipe_sm_io_datapathEn; // @[sm_x426_inr_UnitPipe.scala 33:18:@32670.4]
  wire  x426_inr_UnitPipe_sm_io_ctrInc; // @[sm_x426_inr_UnitPipe.scala 33:18:@32670.4]
  wire  x426_inr_UnitPipe_sm_io_parentAck; // @[sm_x426_inr_UnitPipe.scala 33:18:@32670.4]
  wire  x426_inr_UnitPipe_sm_io_backpressure; // @[sm_x426_inr_UnitPipe.scala 33:18:@32670.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@32727.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@32727.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@32727.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@32727.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@32727.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32735.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32735.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32735.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@32735.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@32735.4]
  wire [63:0] x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_in_x276_outdram_number; // @[sm_x426_inr_UnitPipe.scala 69:24:@32765.4]
  wire  x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_in_x419_valid; // @[sm_x426_inr_UnitPipe.scala 69:24:@32765.4]
  wire [63:0] x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_in_x419_bits_addr; // @[sm_x426_inr_UnitPipe.scala 69:24:@32765.4]
  wire [31:0] x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_in_x419_bits_size; // @[sm_x426_inr_UnitPipe.scala 69:24:@32765.4]
  wire  x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x426_inr_UnitPipe.scala 69:24:@32765.4]
  wire  x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x426_inr_UnitPipe.scala 69:24:@32765.4]
  wire  x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_rr; // @[sm_x426_inr_UnitPipe.scala 69:24:@32765.4]
  wire  x428_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@32833.4]
  wire  x428_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@32833.4]
  wire  x428_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@32833.4]
  wire  x428_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@32833.4]
  wire [22:0] x428_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@32833.4]
  wire  x428_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@32833.4]
  wire  x428_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@32833.4]
  wire  x435_inr_Foreach_sm_clock; // @[sm_x435_inr_Foreach.scala 33:18:@32886.4]
  wire  x435_inr_Foreach_sm_reset; // @[sm_x435_inr_Foreach.scala 33:18:@32886.4]
  wire  x435_inr_Foreach_sm_io_enable; // @[sm_x435_inr_Foreach.scala 33:18:@32886.4]
  wire  x435_inr_Foreach_sm_io_done; // @[sm_x435_inr_Foreach.scala 33:18:@32886.4]
  wire  x435_inr_Foreach_sm_io_doneLatch; // @[sm_x435_inr_Foreach.scala 33:18:@32886.4]
  wire  x435_inr_Foreach_sm_io_ctrDone; // @[sm_x435_inr_Foreach.scala 33:18:@32886.4]
  wire  x435_inr_Foreach_sm_io_datapathEn; // @[sm_x435_inr_Foreach.scala 33:18:@32886.4]
  wire  x435_inr_Foreach_sm_io_ctrInc; // @[sm_x435_inr_Foreach.scala 33:18:@32886.4]
  wire  x435_inr_Foreach_sm_io_ctrRst; // @[sm_x435_inr_Foreach.scala 33:18:@32886.4]
  wire  x435_inr_Foreach_sm_io_parentAck; // @[sm_x435_inr_Foreach.scala 33:18:@32886.4]
  wire  x435_inr_Foreach_sm_io_backpressure; // @[sm_x435_inr_Foreach.scala 33:18:@32886.4]
  wire  x435_inr_Foreach_sm_io_break; // @[sm_x435_inr_Foreach.scala 33:18:@32886.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@32914.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@32914.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@32914.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@32914.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@32914.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@32954.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@32954.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@32954.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@32954.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@32954.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@32962.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@32962.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@32962.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@32962.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@32962.4]
  wire  x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_clock; // @[sm_x435_inr_Foreach.scala 78:24:@32997.4]
  wire  x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_reset; // @[sm_x435_inr_Foreach.scala 78:24:@32997.4]
  wire [20:0] x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x280_outbuf_0_rPort_0_ofs_0; // @[sm_x435_inr_Foreach.scala 78:24:@32997.4]
  wire  x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x280_outbuf_0_rPort_0_en_0; // @[sm_x435_inr_Foreach.scala 78:24:@32997.4]
  wire  x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x280_outbuf_0_rPort_0_backpressure; // @[sm_x435_inr_Foreach.scala 78:24:@32997.4]
  wire [7:0] x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x280_outbuf_0_rPort_0_output_0; // @[sm_x435_inr_Foreach.scala 78:24:@32997.4]
  wire  x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x420_valid; // @[sm_x435_inr_Foreach.scala 78:24:@32997.4]
  wire [7:0] x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x420_bits_wdata_0; // @[sm_x435_inr_Foreach.scala 78:24:@32997.4]
  wire  x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x420_bits_wstrb; // @[sm_x435_inr_Foreach.scala 78:24:@32997.4]
  wire  x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x435_inr_Foreach.scala 78:24:@32997.4]
  wire  x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x435_inr_Foreach.scala 78:24:@32997.4]
  wire  x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x435_inr_Foreach.scala 78:24:@32997.4]
  wire [31:0] x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x435_inr_Foreach.scala 78:24:@32997.4]
  wire  x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x435_inr_Foreach.scala 78:24:@32997.4]
  wire  x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_rr; // @[sm_x435_inr_Foreach.scala 78:24:@32997.4]
  wire  x439_inr_UnitPipe_sm_clock; // @[sm_x439_inr_UnitPipe.scala 32:18:@33117.4]
  wire  x439_inr_UnitPipe_sm_reset; // @[sm_x439_inr_UnitPipe.scala 32:18:@33117.4]
  wire  x439_inr_UnitPipe_sm_io_enable; // @[sm_x439_inr_UnitPipe.scala 32:18:@33117.4]
  wire  x439_inr_UnitPipe_sm_io_done; // @[sm_x439_inr_UnitPipe.scala 32:18:@33117.4]
  wire  x439_inr_UnitPipe_sm_io_doneLatch; // @[sm_x439_inr_UnitPipe.scala 32:18:@33117.4]
  wire  x439_inr_UnitPipe_sm_io_ctrDone; // @[sm_x439_inr_UnitPipe.scala 32:18:@33117.4]
  wire  x439_inr_UnitPipe_sm_io_datapathEn; // @[sm_x439_inr_UnitPipe.scala 32:18:@33117.4]
  wire  x439_inr_UnitPipe_sm_io_ctrInc; // @[sm_x439_inr_UnitPipe.scala 32:18:@33117.4]
  wire  x439_inr_UnitPipe_sm_io_parentAck; // @[sm_x439_inr_UnitPipe.scala 32:18:@33117.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@33174.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@33174.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@33174.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@33174.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@33174.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@33182.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@33182.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@33182.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@33182.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@33182.4]
  wire  x439_inr_UnitPipe_kernelx439_inr_UnitPipe_concrete1_io_in_x421_ready; // @[sm_x439_inr_UnitPipe.scala 60:24:@33212.4]
  wire  x439_inr_UnitPipe_kernelx439_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x439_inr_UnitPipe.scala 60:24:@33212.4]
  wire  _T_359; // @[package.scala 100:49:@32698.4]
  reg  _T_362; // @[package.scala 48:56:@32699.4]
  reg [31:0] _RAND_0;
  wire  _T_375; // @[package.scala 96:25:@32732.4 package.scala 96:25:@32733.4]
  wire  _T_381; // @[package.scala 96:25:@32740.4 package.scala 96:25:@32741.4]
  wire  _T_384; // @[SpatialBlocks.scala 138:93:@32743.4]
  wire  _T_454; // @[package.scala 96:25:@32919.4 package.scala 96:25:@32920.4]
  wire  _T_468; // @[package.scala 96:25:@32959.4 package.scala 96:25:@32960.4]
  wire  _T_474; // @[package.scala 96:25:@32967.4 package.scala 96:25:@32968.4]
  wire  _T_477; // @[SpatialBlocks.scala 138:93:@32970.4]
  wire  _T_479; // @[SpatialBlocks.scala 157:36:@32979.4]
  wire  _T_480; // @[SpatialBlocks.scala 157:78:@32980.4]
  wire  _T_547; // @[package.scala 100:49:@33145.4]
  reg  _T_550; // @[package.scala 48:56:@33146.4]
  reg [31:0] _RAND_1;
  wire  x439_inr_UnitPipe_sigsIn_forwardpressure; // @[sm_x440_outr_UnitPipe.scala 101:55:@33152.4]
  wire  _T_563; // @[package.scala 96:25:@33179.4 package.scala 96:25:@33180.4]
  wire  _T_569; // @[package.scala 96:25:@33187.4 package.scala 96:25:@33188.4]
  wire  _T_572; // @[SpatialBlocks.scala 138:93:@33190.4]
  wire  x439_inr_UnitPipe_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@33191.4]
  x426_inr_UnitPipe_sm x426_inr_UnitPipe_sm ( // @[sm_x426_inr_UnitPipe.scala 33:18:@32670.4]
    .clock(x426_inr_UnitPipe_sm_clock),
    .reset(x426_inr_UnitPipe_sm_reset),
    .io_enable(x426_inr_UnitPipe_sm_io_enable),
    .io_done(x426_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x426_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x426_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x426_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x426_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x426_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x426_inr_UnitPipe_sm_io_backpressure)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@32727.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@32735.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1 x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1 ( // @[sm_x426_inr_UnitPipe.scala 69:24:@32765.4]
    .io_in_x276_outdram_number(x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_in_x276_outdram_number),
    .io_in_x419_valid(x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_in_x419_valid),
    .io_in_x419_bits_addr(x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_in_x419_bits_addr),
    .io_in_x419_bits_size(x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_in_x419_bits_size),
    .io_sigsIn_backpressure(x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_rr(x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_rr)
  );
  x428_ctrchain x428_ctrchain ( // @[SpatialBlocks.scala 37:22:@32833.4]
    .clock(x428_ctrchain_clock),
    .reset(x428_ctrchain_reset),
    .io_input_reset(x428_ctrchain_io_input_reset),
    .io_input_enable(x428_ctrchain_io_input_enable),
    .io_output_counts_0(x428_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x428_ctrchain_io_output_oobs_0),
    .io_output_done(x428_ctrchain_io_output_done)
  );
  x435_inr_Foreach_sm x435_inr_Foreach_sm ( // @[sm_x435_inr_Foreach.scala 33:18:@32886.4]
    .clock(x435_inr_Foreach_sm_clock),
    .reset(x435_inr_Foreach_sm_reset),
    .io_enable(x435_inr_Foreach_sm_io_enable),
    .io_done(x435_inr_Foreach_sm_io_done),
    .io_doneLatch(x435_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x435_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x435_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x435_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x435_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x435_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x435_inr_Foreach_sm_io_backpressure),
    .io_break(x435_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@32914.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@32954.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@32962.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x435_inr_Foreach_kernelx435_inr_Foreach_concrete1 x435_inr_Foreach_kernelx435_inr_Foreach_concrete1 ( // @[sm_x435_inr_Foreach.scala 78:24:@32997.4]
    .clock(x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_clock),
    .reset(x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_reset),
    .io_in_x280_outbuf_0_rPort_0_ofs_0(x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x280_outbuf_0_rPort_0_ofs_0),
    .io_in_x280_outbuf_0_rPort_0_en_0(x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x280_outbuf_0_rPort_0_en_0),
    .io_in_x280_outbuf_0_rPort_0_backpressure(x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x280_outbuf_0_rPort_0_backpressure),
    .io_in_x280_outbuf_0_rPort_0_output_0(x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x280_outbuf_0_rPort_0_output_0),
    .io_in_x420_valid(x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x420_valid),
    .io_in_x420_bits_wdata_0(x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x420_bits_wdata_0),
    .io_in_x420_bits_wstrb(x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x420_bits_wstrb),
    .io_sigsIn_backpressure(x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_rr)
  );
  x439_inr_UnitPipe_sm x439_inr_UnitPipe_sm ( // @[sm_x439_inr_UnitPipe.scala 32:18:@33117.4]
    .clock(x439_inr_UnitPipe_sm_clock),
    .reset(x439_inr_UnitPipe_sm_reset),
    .io_enable(x439_inr_UnitPipe_sm_io_enable),
    .io_done(x439_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x439_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x439_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x439_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x439_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x439_inr_UnitPipe_sm_io_parentAck)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@33174.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@33182.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x439_inr_UnitPipe_kernelx439_inr_UnitPipe_concrete1 x439_inr_UnitPipe_kernelx439_inr_UnitPipe_concrete1 ( // @[sm_x439_inr_UnitPipe.scala 60:24:@33212.4]
    .io_in_x421_ready(x439_inr_UnitPipe_kernelx439_inr_UnitPipe_concrete1_io_in_x421_ready),
    .io_sigsIn_datapathEn(x439_inr_UnitPipe_kernelx439_inr_UnitPipe_concrete1_io_sigsIn_datapathEn)
  );
  assign _T_359 = x426_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@32698.4]
  assign _T_375 = RetimeWrapper_io_out; // @[package.scala 96:25:@32732.4 package.scala 96:25:@32733.4]
  assign _T_381 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@32740.4 package.scala 96:25:@32741.4]
  assign _T_384 = ~ _T_381; // @[SpatialBlocks.scala 138:93:@32743.4]
  assign _T_454 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@32919.4 package.scala 96:25:@32920.4]
  assign _T_468 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@32959.4 package.scala 96:25:@32960.4]
  assign _T_474 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@32967.4 package.scala 96:25:@32968.4]
  assign _T_477 = ~ _T_474; // @[SpatialBlocks.scala 138:93:@32970.4]
  assign _T_479 = x435_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@32979.4]
  assign _T_480 = ~ x435_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@32980.4]
  assign _T_547 = x439_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@33145.4]
  assign x439_inr_UnitPipe_sigsIn_forwardpressure = io_in_x421_valid | x439_inr_UnitPipe_sm_io_doneLatch; // @[sm_x440_outr_UnitPipe.scala 101:55:@33152.4]
  assign _T_563 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@33179.4 package.scala 96:25:@33180.4]
  assign _T_569 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@33187.4 package.scala 96:25:@33188.4]
  assign _T_572 = ~ _T_569; // @[SpatialBlocks.scala 138:93:@33190.4]
  assign x439_inr_UnitPipe_sigsIn_baseEn = _T_563 & _T_572; // @[SpatialBlocks.scala 138:90:@33191.4]
  assign io_in_x421_ready = x439_inr_UnitPipe_kernelx439_inr_UnitPipe_concrete1_io_in_x421_ready; // @[sm_x439_inr_UnitPipe.scala 46:23:@33248.4]
  assign io_in_x280_outbuf_0_rPort_0_ofs_0 = x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x280_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@33048.4]
  assign io_in_x280_outbuf_0_rPort_0_en_0 = x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x280_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@33047.4]
  assign io_in_x280_outbuf_0_rPort_0_backpressure = x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x280_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@33046.4]
  assign io_in_x420_valid = x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x420_valid; // @[sm_x435_inr_Foreach.scala 50:23:@33052.4]
  assign io_in_x420_bits_wdata_0 = x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x420_bits_wdata_0; // @[sm_x435_inr_Foreach.scala 50:23:@33051.4]
  assign io_in_x420_bits_wstrb = x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x420_bits_wstrb; // @[sm_x435_inr_Foreach.scala 50:23:@33050.4]
  assign io_in_x419_valid = x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_in_x419_valid; // @[sm_x426_inr_UnitPipe.scala 50:23:@32804.4]
  assign io_in_x419_bits_addr = x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_in_x419_bits_addr; // @[sm_x426_inr_UnitPipe.scala 50:23:@32803.4]
  assign io_in_x419_bits_size = x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_in_x419_bits_size; // @[sm_x426_inr_UnitPipe.scala 50:23:@32802.4]
  assign io_sigsOut_smDoneIn_0 = x426_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@32750.4]
  assign io_sigsOut_smDoneIn_1 = x435_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@32977.4]
  assign io_sigsOut_smDoneIn_2 = x439_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@33197.4]
  assign io_sigsOut_smCtrCopyDone_0 = x426_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@32764.4]
  assign io_sigsOut_smCtrCopyDone_1 = x435_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@32996.4]
  assign io_sigsOut_smCtrCopyDone_2 = x439_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@33211.4]
  assign x426_inr_UnitPipe_sm_clock = clock; // @[:@32671.4]
  assign x426_inr_UnitPipe_sm_reset = reset; // @[:@32672.4]
  assign x426_inr_UnitPipe_sm_io_enable = _T_375 & _T_384; // @[SpatialBlocks.scala 140:18:@32747.4]
  assign x426_inr_UnitPipe_sm_io_ctrDone = x426_inr_UnitPipe_sm_io_ctrInc & _T_362; // @[sm_x440_outr_UnitPipe.scala 77:39:@32702.4]
  assign x426_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@32749.4]
  assign x426_inr_UnitPipe_sm_io_backpressure = io_in_x419_ready | x426_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@32721.4]
  assign RetimeWrapper_clock = clock; // @[:@32728.4]
  assign RetimeWrapper_reset = reset; // @[:@32729.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@32731.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@32730.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32736.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32737.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@32739.4]
  assign RetimeWrapper_1_io_in = x426_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@32738.4]
  assign x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_in_x276_outdram_number = io_in_x276_outdram_number; // @[sm_x426_inr_UnitPipe.scala 49:31:@32801.4]
  assign x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x419_ready | x426_inr_UnitPipe_sm_io_doneLatch; // @[sm_x426_inr_UnitPipe.scala 74:22:@32820.4]
  assign x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x426_inr_UnitPipe_sm_io_datapathEn; // @[sm_x426_inr_UnitPipe.scala 74:22:@32818.4]
  assign x426_inr_UnitPipe_kernelx426_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x426_inr_UnitPipe.scala 73:18:@32806.4]
  assign x428_ctrchain_clock = clock; // @[:@32834.4]
  assign x428_ctrchain_reset = reset; // @[:@32835.4]
  assign x428_ctrchain_io_input_reset = x435_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@32995.4]
  assign x428_ctrchain_io_input_enable = x435_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@32947.4 SpatialBlocks.scala 159:42:@32994.4]
  assign x435_inr_Foreach_sm_clock = clock; // @[:@32887.4]
  assign x435_inr_Foreach_sm_reset = reset; // @[:@32888.4]
  assign x435_inr_Foreach_sm_io_enable = _T_468 & _T_477; // @[SpatialBlocks.scala 140:18:@32974.4]
  assign x435_inr_Foreach_sm_io_ctrDone = io_rr ? _T_454 : 1'h0; // @[sm_x440_outr_UnitPipe.scala 90:38:@32922.4]
  assign x435_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@32976.4]
  assign x435_inr_Foreach_sm_io_backpressure = io_in_x420_ready | x435_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@32948.4]
  assign x435_inr_Foreach_sm_io_break = 1'h0; // @[sm_x440_outr_UnitPipe.scala 94:36:@32928.4]
  assign RetimeWrapper_2_clock = clock; // @[:@32915.4]
  assign RetimeWrapper_2_reset = reset; // @[:@32916.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@32918.4]
  assign RetimeWrapper_2_io_in = x428_ctrchain_io_output_done; // @[package.scala 94:16:@32917.4]
  assign RetimeWrapper_3_clock = clock; // @[:@32955.4]
  assign RetimeWrapper_3_reset = reset; // @[:@32956.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@32958.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@32957.4]
  assign RetimeWrapper_4_clock = clock; // @[:@32963.4]
  assign RetimeWrapper_4_reset = reset; // @[:@32964.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@32966.4]
  assign RetimeWrapper_4_io_in = x435_inr_Foreach_sm_io_done; // @[package.scala 94:16:@32965.4]
  assign x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_clock = clock; // @[:@32998.4]
  assign x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_reset = reset; // @[:@32999.4]
  assign x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_in_x280_outbuf_0_rPort_0_output_0 = io_in_x280_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@33045.4]
  assign x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x420_ready | x435_inr_Foreach_sm_io_doneLatch; // @[sm_x435_inr_Foreach.scala 83:22:@33068.4]
  assign x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_479 & _T_480; // @[sm_x435_inr_Foreach.scala 83:22:@33066.4]
  assign x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_sigsIn_break = x435_inr_Foreach_sm_io_break; // @[sm_x435_inr_Foreach.scala 83:22:@33064.4]
  assign x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{9{x428_ctrchain_io_output_counts_0[22]}},x428_ctrchain_io_output_counts_0}; // @[sm_x435_inr_Foreach.scala 83:22:@33059.4]
  assign x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x428_ctrchain_io_output_oobs_0; // @[sm_x435_inr_Foreach.scala 83:22:@33058.4]
  assign x435_inr_Foreach_kernelx435_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x435_inr_Foreach.scala 82:18:@33054.4]
  assign x439_inr_UnitPipe_sm_clock = clock; // @[:@33118.4]
  assign x439_inr_UnitPipe_sm_reset = reset; // @[:@33119.4]
  assign x439_inr_UnitPipe_sm_io_enable = x439_inr_UnitPipe_sigsIn_baseEn & x439_inr_UnitPipe_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@33194.4]
  assign x439_inr_UnitPipe_sm_io_ctrDone = x439_inr_UnitPipe_sm_io_ctrInc & _T_550; // @[sm_x440_outr_UnitPipe.scala 99:39:@33149.4]
  assign x439_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 142:21:@33196.4]
  assign RetimeWrapper_5_clock = clock; // @[:@33175.4]
  assign RetimeWrapper_5_reset = reset; // @[:@33176.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@33178.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@33177.4]
  assign RetimeWrapper_6_clock = clock; // @[:@33183.4]
  assign RetimeWrapper_6_reset = reset; // @[:@33184.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@33186.4]
  assign RetimeWrapper_6_io_in = x439_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@33185.4]
  assign x439_inr_UnitPipe_kernelx439_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x439_inr_UnitPipe_sm_io_datapathEn; // @[sm_x439_inr_UnitPipe.scala 65:22:@33261.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_362 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_550 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_362 <= 1'h0;
    end else begin
      _T_362 <= _T_359;
    end
    if (reset) begin
      _T_550 <= 1'h0;
    end else begin
      _T_550 <= _T_547;
    end
  end
endmodule
module x556_kernelx556_concrete1( // @[:@33277.2]
  input          clock, // @[:@33278.4]
  input          reset, // @[:@33279.4]
  input  [63:0]  io_in_x276_outdram_number, // @[:@33280.4]
  output         io_in_x421_ready, // @[:@33280.4]
  input          io_in_x421_valid, // @[:@33280.4]
  output [20:0]  io_in_x280_outbuf_0_rPort_0_ofs_0, // @[:@33280.4]
  output         io_in_x280_outbuf_0_rPort_0_en_0, // @[:@33280.4]
  output         io_in_x280_outbuf_0_rPort_0_backpressure, // @[:@33280.4]
  input  [7:0]   io_in_x280_outbuf_0_rPort_0_output_0, // @[:@33280.4]
  input          io_in_x420_ready, // @[:@33280.4]
  output         io_in_x420_valid, // @[:@33280.4]
  output [7:0]   io_in_x420_bits_wdata_0, // @[:@33280.4]
  output         io_in_x420_bits_wstrb, // @[:@33280.4]
  output         io_in_x279_TVALID, // @[:@33280.4]
  input          io_in_x279_TREADY, // @[:@33280.4]
  output [255:0] io_in_x279_TDATA, // @[:@33280.4]
  input          io_in_x419_ready, // @[:@33280.4]
  output         io_in_x419_valid, // @[:@33280.4]
  output [63:0]  io_in_x419_bits_addr, // @[:@33280.4]
  output [31:0]  io_in_x419_bits_size, // @[:@33280.4]
  input          io_in_x278_TVALID, // @[:@33280.4]
  output         io_in_x278_TREADY, // @[:@33280.4]
  input  [255:0] io_in_x278_TDATA, // @[:@33280.4]
  input  [7:0]   io_in_x278_TID, // @[:@33280.4]
  input  [7:0]   io_in_x278_TDEST, // @[:@33280.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@33280.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@33280.4]
  input          io_sigsIn_smChildAcks_0, // @[:@33280.4]
  input          io_sigsIn_smChildAcks_1, // @[:@33280.4]
  output         io_sigsOut_smDoneIn_0, // @[:@33280.4]
  output         io_sigsOut_smDoneIn_1, // @[:@33280.4]
  input          io_rr // @[:@33280.4]
);
  wire  x418_outr_UnitPipe_sm_clock; // @[sm_x418_outr_UnitPipe.scala 32:18:@33353.4]
  wire  x418_outr_UnitPipe_sm_reset; // @[sm_x418_outr_UnitPipe.scala 32:18:@33353.4]
  wire  x418_outr_UnitPipe_sm_io_enable; // @[sm_x418_outr_UnitPipe.scala 32:18:@33353.4]
  wire  x418_outr_UnitPipe_sm_io_done; // @[sm_x418_outr_UnitPipe.scala 32:18:@33353.4]
  wire  x418_outr_UnitPipe_sm_io_parentAck; // @[sm_x418_outr_UnitPipe.scala 32:18:@33353.4]
  wire  x418_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x418_outr_UnitPipe.scala 32:18:@33353.4]
  wire  x418_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x418_outr_UnitPipe.scala 32:18:@33353.4]
  wire  x418_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x418_outr_UnitPipe.scala 32:18:@33353.4]
  wire  x418_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x418_outr_UnitPipe.scala 32:18:@33353.4]
  wire  x418_outr_UnitPipe_sm_io_childAck_0; // @[sm_x418_outr_UnitPipe.scala 32:18:@33353.4]
  wire  x418_outr_UnitPipe_sm_io_childAck_1; // @[sm_x418_outr_UnitPipe.scala 32:18:@33353.4]
  wire  x418_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x418_outr_UnitPipe.scala 32:18:@33353.4]
  wire  x418_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x418_outr_UnitPipe.scala 32:18:@33353.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@33415.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@33415.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@33415.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@33415.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@33415.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@33423.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@33423.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@33423.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@33423.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@33423.4]
  wire  x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_clock; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire  x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_reset; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire  x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x279_TVALID; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire  x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x279_TREADY; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire [255:0] x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x279_TDATA; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire  x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x278_TVALID; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire  x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x278_TREADY; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire [255:0] x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x278_TDATA; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire [7:0] x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x278_TID; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire [7:0] x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x278_TDEST; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire  x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire  x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire  x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire  x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire  x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire  x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire  x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire  x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire  x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_rr; // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
  wire  x440_outr_UnitPipe_sm_clock; // @[sm_x440_outr_UnitPipe.scala 36:18:@33632.4]
  wire  x440_outr_UnitPipe_sm_reset; // @[sm_x440_outr_UnitPipe.scala 36:18:@33632.4]
  wire  x440_outr_UnitPipe_sm_io_enable; // @[sm_x440_outr_UnitPipe.scala 36:18:@33632.4]
  wire  x440_outr_UnitPipe_sm_io_done; // @[sm_x440_outr_UnitPipe.scala 36:18:@33632.4]
  wire  x440_outr_UnitPipe_sm_io_parentAck; // @[sm_x440_outr_UnitPipe.scala 36:18:@33632.4]
  wire  x440_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x440_outr_UnitPipe.scala 36:18:@33632.4]
  wire  x440_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x440_outr_UnitPipe.scala 36:18:@33632.4]
  wire  x440_outr_UnitPipe_sm_io_doneIn_2; // @[sm_x440_outr_UnitPipe.scala 36:18:@33632.4]
  wire  x440_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x440_outr_UnitPipe.scala 36:18:@33632.4]
  wire  x440_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x440_outr_UnitPipe.scala 36:18:@33632.4]
  wire  x440_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x440_outr_UnitPipe.scala 36:18:@33632.4]
  wire  x440_outr_UnitPipe_sm_io_childAck_0; // @[sm_x440_outr_UnitPipe.scala 36:18:@33632.4]
  wire  x440_outr_UnitPipe_sm_io_childAck_1; // @[sm_x440_outr_UnitPipe.scala 36:18:@33632.4]
  wire  x440_outr_UnitPipe_sm_io_childAck_2; // @[sm_x440_outr_UnitPipe.scala 36:18:@33632.4]
  wire  x440_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x440_outr_UnitPipe.scala 36:18:@33632.4]
  wire  x440_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x440_outr_UnitPipe.scala 36:18:@33632.4]
  wire  x440_outr_UnitPipe_sm_io_ctrCopyDone_2; // @[sm_x440_outr_UnitPipe.scala 36:18:@33632.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@33704.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@33704.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@33704.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@33704.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@33704.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@33712.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@33712.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@33712.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@33712.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@33712.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_clock; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_reset; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire [63:0] x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x276_outdram_number; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x421_ready; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x421_valid; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire [20:0] x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x280_outbuf_0_rPort_0_ofs_0; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x280_outbuf_0_rPort_0_en_0; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x280_outbuf_0_rPort_0_backpressure; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire [7:0] x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x280_outbuf_0_rPort_0_output_0; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x420_ready; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x420_valid; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire [7:0] x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x420_bits_wdata_0; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x420_bits_wstrb; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x419_ready; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x419_valid; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire [63:0] x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x419_bits_addr; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire [31:0] x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x419_bits_size; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_rr; // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
  wire  _T_408; // @[package.scala 96:25:@33420.4 package.scala 96:25:@33421.4]
  wire  _T_414; // @[package.scala 96:25:@33428.4 package.scala 96:25:@33429.4]
  wire  _T_417; // @[SpatialBlocks.scala 138:93:@33431.4]
  wire  _T_508; // @[package.scala 96:25:@33709.4 package.scala 96:25:@33710.4]
  wire  _T_514; // @[package.scala 96:25:@33717.4 package.scala 96:25:@33718.4]
  wire  _T_517; // @[SpatialBlocks.scala 138:93:@33720.4]
  x418_outr_UnitPipe_sm x418_outr_UnitPipe_sm ( // @[sm_x418_outr_UnitPipe.scala 32:18:@33353.4]
    .clock(x418_outr_UnitPipe_sm_clock),
    .reset(x418_outr_UnitPipe_sm_reset),
    .io_enable(x418_outr_UnitPipe_sm_io_enable),
    .io_done(x418_outr_UnitPipe_sm_io_done),
    .io_parentAck(x418_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x418_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x418_outr_UnitPipe_sm_io_doneIn_1),
    .io_enableOut_0(x418_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x418_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x418_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x418_outr_UnitPipe_sm_io_childAck_1),
    .io_ctrCopyDone_0(x418_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x418_outr_UnitPipe_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@33415.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@33423.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1 x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1 ( // @[sm_x418_outr_UnitPipe.scala 87:24:@33454.4]
    .clock(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_clock),
    .reset(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_reset),
    .io_in_x279_TVALID(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x279_TVALID),
    .io_in_x279_TREADY(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x279_TREADY),
    .io_in_x279_TDATA(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x279_TDATA),
    .io_in_x278_TVALID(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x278_TVALID),
    .io_in_x278_TREADY(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x278_TREADY),
    .io_in_x278_TDATA(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x278_TDATA),
    .io_in_x278_TID(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x278_TID),
    .io_in_x278_TDEST(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x278_TDEST),
    .io_sigsIn_smEnableOuts_0(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_rr)
  );
  x440_outr_UnitPipe_sm x440_outr_UnitPipe_sm ( // @[sm_x440_outr_UnitPipe.scala 36:18:@33632.4]
    .clock(x440_outr_UnitPipe_sm_clock),
    .reset(x440_outr_UnitPipe_sm_reset),
    .io_enable(x440_outr_UnitPipe_sm_io_enable),
    .io_done(x440_outr_UnitPipe_sm_io_done),
    .io_parentAck(x440_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x440_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x440_outr_UnitPipe_sm_io_doneIn_1),
    .io_doneIn_2(x440_outr_UnitPipe_sm_io_doneIn_2),
    .io_enableOut_0(x440_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x440_outr_UnitPipe_sm_io_enableOut_1),
    .io_enableOut_2(x440_outr_UnitPipe_sm_io_enableOut_2),
    .io_childAck_0(x440_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x440_outr_UnitPipe_sm_io_childAck_1),
    .io_childAck_2(x440_outr_UnitPipe_sm_io_childAck_2),
    .io_ctrCopyDone_0(x440_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x440_outr_UnitPipe_sm_io_ctrCopyDone_1),
    .io_ctrCopyDone_2(x440_outr_UnitPipe_sm_io_ctrCopyDone_2)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@33704.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@33712.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1 x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1 ( // @[sm_x440_outr_UnitPipe.scala 108:24:@33744.4]
    .clock(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_clock),
    .reset(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_reset),
    .io_in_x276_outdram_number(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x276_outdram_number),
    .io_in_x421_ready(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x421_ready),
    .io_in_x421_valid(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x421_valid),
    .io_in_x280_outbuf_0_rPort_0_ofs_0(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x280_outbuf_0_rPort_0_ofs_0),
    .io_in_x280_outbuf_0_rPort_0_en_0(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x280_outbuf_0_rPort_0_en_0),
    .io_in_x280_outbuf_0_rPort_0_backpressure(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x280_outbuf_0_rPort_0_backpressure),
    .io_in_x280_outbuf_0_rPort_0_output_0(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x280_outbuf_0_rPort_0_output_0),
    .io_in_x420_ready(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x420_ready),
    .io_in_x420_valid(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x420_valid),
    .io_in_x420_bits_wdata_0(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x420_bits_wdata_0),
    .io_in_x420_bits_wstrb(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x420_bits_wstrb),
    .io_in_x419_ready(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x419_ready),
    .io_in_x419_valid(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x419_valid),
    .io_in_x419_bits_addr(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x419_bits_addr),
    .io_in_x419_bits_size(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x419_bits_size),
    .io_sigsIn_smEnableOuts_0(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smCtrCopyDone_0(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_sigsOut_smCtrCopyDone_2(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2),
    .io_rr(x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_408 = RetimeWrapper_io_out; // @[package.scala 96:25:@33420.4 package.scala 96:25:@33421.4]
  assign _T_414 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@33428.4 package.scala 96:25:@33429.4]
  assign _T_417 = ~ _T_414; // @[SpatialBlocks.scala 138:93:@33431.4]
  assign _T_508 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@33709.4 package.scala 96:25:@33710.4]
  assign _T_514 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@33717.4 package.scala 96:25:@33718.4]
  assign _T_517 = ~ _T_514; // @[SpatialBlocks.scala 138:93:@33720.4]
  assign io_in_x421_ready = x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x421_ready; // @[sm_x440_outr_UnitPipe.scala 59:23:@33827.4]
  assign io_in_x280_outbuf_0_rPort_0_ofs_0 = x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x280_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@33831.4]
  assign io_in_x280_outbuf_0_rPort_0_en_0 = x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x280_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@33830.4]
  assign io_in_x280_outbuf_0_rPort_0_backpressure = x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x280_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@33829.4]
  assign io_in_x420_valid = x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x420_valid; // @[sm_x440_outr_UnitPipe.scala 61:23:@33835.4]
  assign io_in_x420_bits_wdata_0 = x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x420_bits_wdata_0; // @[sm_x440_outr_UnitPipe.scala 61:23:@33834.4]
  assign io_in_x420_bits_wstrb = x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x420_bits_wstrb; // @[sm_x440_outr_UnitPipe.scala 61:23:@33833.4]
  assign io_in_x279_TVALID = x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x279_TVALID; // @[sm_x418_outr_UnitPipe.scala 48:23:@33523.4]
  assign io_in_x279_TDATA = x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x279_TDATA; // @[sm_x418_outr_UnitPipe.scala 48:23:@33521.4]
  assign io_in_x419_valid = x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x419_valid; // @[sm_x440_outr_UnitPipe.scala 62:23:@33839.4]
  assign io_in_x419_bits_addr = x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x419_bits_addr; // @[sm_x440_outr_UnitPipe.scala 62:23:@33838.4]
  assign io_in_x419_bits_size = x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x419_bits_size; // @[sm_x440_outr_UnitPipe.scala 62:23:@33837.4]
  assign io_in_x278_TREADY = x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x278_TREADY; // @[sm_x418_outr_UnitPipe.scala 49:23:@33531.4]
  assign io_sigsOut_smDoneIn_0 = x418_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@33438.4]
  assign io_sigsOut_smDoneIn_1 = x440_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@33727.4]
  assign x418_outr_UnitPipe_sm_clock = clock; // @[:@33354.4]
  assign x418_outr_UnitPipe_sm_reset = reset; // @[:@33355.4]
  assign x418_outr_UnitPipe_sm_io_enable = _T_408 & _T_417; // @[SpatialBlocks.scala 140:18:@33435.4]
  assign x418_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@33437.4]
  assign x418_outr_UnitPipe_sm_io_doneIn_0 = x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@33405.4]
  assign x418_outr_UnitPipe_sm_io_doneIn_1 = x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@33406.4]
  assign x418_outr_UnitPipe_sm_io_ctrCopyDone_0 = x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@33452.4]
  assign x418_outr_UnitPipe_sm_io_ctrCopyDone_1 = x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@33453.4]
  assign RetimeWrapper_clock = clock; // @[:@33416.4]
  assign RetimeWrapper_reset = reset; // @[:@33417.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@33419.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@33418.4]
  assign RetimeWrapper_1_clock = clock; // @[:@33424.4]
  assign RetimeWrapper_1_reset = reset; // @[:@33425.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@33427.4]
  assign RetimeWrapper_1_io_in = x418_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@33426.4]
  assign x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_clock = clock; // @[:@33455.4]
  assign x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_reset = reset; // @[:@33456.4]
  assign x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x279_TREADY = io_in_x279_TREADY; // @[sm_x418_outr_UnitPipe.scala 48:23:@33522.4]
  assign x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x278_TVALID = io_in_x278_TVALID; // @[sm_x418_outr_UnitPipe.scala 49:23:@33532.4]
  assign x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x278_TDATA = io_in_x278_TDATA; // @[sm_x418_outr_UnitPipe.scala 49:23:@33530.4]
  assign x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x278_TID = io_in_x278_TID; // @[sm_x418_outr_UnitPipe.scala 49:23:@33526.4]
  assign x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_in_x278_TDEST = io_in_x278_TDEST; // @[sm_x418_outr_UnitPipe.scala 49:23:@33525.4]
  assign x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x418_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x418_outr_UnitPipe.scala 92:22:@33548.4]
  assign x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x418_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x418_outr_UnitPipe.scala 92:22:@33549.4]
  assign x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x418_outr_UnitPipe_sm_io_childAck_0; // @[sm_x418_outr_UnitPipe.scala 92:22:@33544.4]
  assign x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x418_outr_UnitPipe_sm_io_childAck_1; // @[sm_x418_outr_UnitPipe.scala 92:22:@33545.4]
  assign x418_outr_UnitPipe_kernelx418_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x418_outr_UnitPipe.scala 91:18:@33533.4]
  assign x440_outr_UnitPipe_sm_clock = clock; // @[:@33633.4]
  assign x440_outr_UnitPipe_sm_reset = reset; // @[:@33634.4]
  assign x440_outr_UnitPipe_sm_io_enable = _T_508 & _T_517; // @[SpatialBlocks.scala 140:18:@33724.4]
  assign x440_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@33726.4]
  assign x440_outr_UnitPipe_sm_io_doneIn_0 = x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@33692.4]
  assign x440_outr_UnitPipe_sm_io_doneIn_1 = x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@33693.4]
  assign x440_outr_UnitPipe_sm_io_doneIn_2 = x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:67:@33694.4]
  assign x440_outr_UnitPipe_sm_io_ctrCopyDone_0 = x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@33741.4]
  assign x440_outr_UnitPipe_sm_io_ctrCopyDone_1 = x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@33742.4]
  assign x440_outr_UnitPipe_sm_io_ctrCopyDone_2 = x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[SpatialBlocks.scala 161:90:@33743.4]
  assign RetimeWrapper_2_clock = clock; // @[:@33705.4]
  assign RetimeWrapper_2_reset = reset; // @[:@33706.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@33708.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@33707.4]
  assign RetimeWrapper_3_clock = clock; // @[:@33713.4]
  assign RetimeWrapper_3_reset = reset; // @[:@33714.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@33716.4]
  assign RetimeWrapper_3_io_in = x440_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@33715.4]
  assign x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_clock = clock; // @[:@33745.4]
  assign x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_reset = reset; // @[:@33746.4]
  assign x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x276_outdram_number = io_in_x276_outdram_number; // @[sm_x440_outr_UnitPipe.scala 58:31:@33824.4]
  assign x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x421_valid = io_in_x421_valid; // @[sm_x440_outr_UnitPipe.scala 59:23:@33826.4]
  assign x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x280_outbuf_0_rPort_0_output_0 = io_in_x280_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@33828.4]
  assign x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x420_ready = io_in_x420_ready; // @[sm_x440_outr_UnitPipe.scala 61:23:@33836.4]
  assign x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_in_x419_ready = io_in_x419_ready; // @[sm_x440_outr_UnitPipe.scala 62:23:@33840.4]
  assign x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x440_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x440_outr_UnitPipe.scala 113:22:@33863.4]
  assign x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x440_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x440_outr_UnitPipe.scala 113:22:@33864.4]
  assign x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2 = x440_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x440_outr_UnitPipe.scala 113:22:@33865.4]
  assign x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x440_outr_UnitPipe_sm_io_childAck_0; // @[sm_x440_outr_UnitPipe.scala 113:22:@33857.4]
  assign x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x440_outr_UnitPipe_sm_io_childAck_1; // @[sm_x440_outr_UnitPipe.scala 113:22:@33858.4]
  assign x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2 = x440_outr_UnitPipe_sm_io_childAck_2; // @[sm_x440_outr_UnitPipe.scala 113:22:@33859.4]
  assign x440_outr_UnitPipe_kernelx440_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x440_outr_UnitPipe.scala 112:18:@33841.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@33893.2]
  input          clock, // @[:@33894.4]
  input          reset, // @[:@33895.4]
  input  [63:0]  io_in_x276_outdram_number, // @[:@33896.4]
  output         io_in_x421_ready, // @[:@33896.4]
  input          io_in_x421_valid, // @[:@33896.4]
  input          io_in_x420_ready, // @[:@33896.4]
  output         io_in_x420_valid, // @[:@33896.4]
  output [7:0]   io_in_x420_bits_wdata_0, // @[:@33896.4]
  output         io_in_x420_bits_wstrb, // @[:@33896.4]
  output         io_in_x279_TVALID, // @[:@33896.4]
  input          io_in_x279_TREADY, // @[:@33896.4]
  output [255:0] io_in_x279_TDATA, // @[:@33896.4]
  input          io_in_x419_ready, // @[:@33896.4]
  output         io_in_x419_valid, // @[:@33896.4]
  output [63:0]  io_in_x419_bits_addr, // @[:@33896.4]
  output [31:0]  io_in_x419_bits_size, // @[:@33896.4]
  input          io_in_x278_TVALID, // @[:@33896.4]
  output         io_in_x278_TREADY, // @[:@33896.4]
  input  [255:0] io_in_x278_TDATA, // @[:@33896.4]
  input  [7:0]   io_in_x278_TID, // @[:@33896.4]
  input  [7:0]   io_in_x278_TDEST, // @[:@33896.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@33896.4]
  input          io_sigsIn_smChildAcks_0, // @[:@33896.4]
  output         io_sigsOut_smDoneIn_0, // @[:@33896.4]
  input          io_rr // @[:@33896.4]
);
  wire  x280_outbuf_0_clock; // @[m_x280_outbuf_0.scala 27:17:@33906.4]
  wire  x280_outbuf_0_reset; // @[m_x280_outbuf_0.scala 27:17:@33906.4]
  wire [20:0] x280_outbuf_0_io_rPort_0_ofs_0; // @[m_x280_outbuf_0.scala 27:17:@33906.4]
  wire  x280_outbuf_0_io_rPort_0_en_0; // @[m_x280_outbuf_0.scala 27:17:@33906.4]
  wire  x280_outbuf_0_io_rPort_0_backpressure; // @[m_x280_outbuf_0.scala 27:17:@33906.4]
  wire [7:0] x280_outbuf_0_io_rPort_0_output_0; // @[m_x280_outbuf_0.scala 27:17:@33906.4]
  wire  x556_sm_clock; // @[sm_x556.scala 37:18:@33964.4]
  wire  x556_sm_reset; // @[sm_x556.scala 37:18:@33964.4]
  wire  x556_sm_io_enable; // @[sm_x556.scala 37:18:@33964.4]
  wire  x556_sm_io_done; // @[sm_x556.scala 37:18:@33964.4]
  wire  x556_sm_io_ctrDone; // @[sm_x556.scala 37:18:@33964.4]
  wire  x556_sm_io_ctrInc; // @[sm_x556.scala 37:18:@33964.4]
  wire  x556_sm_io_parentAck; // @[sm_x556.scala 37:18:@33964.4]
  wire  x556_sm_io_doneIn_0; // @[sm_x556.scala 37:18:@33964.4]
  wire  x556_sm_io_doneIn_1; // @[sm_x556.scala 37:18:@33964.4]
  wire  x556_sm_io_enableOut_0; // @[sm_x556.scala 37:18:@33964.4]
  wire  x556_sm_io_enableOut_1; // @[sm_x556.scala 37:18:@33964.4]
  wire  x556_sm_io_childAck_0; // @[sm_x556.scala 37:18:@33964.4]
  wire  x556_sm_io_childAck_1; // @[sm_x556.scala 37:18:@33964.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@34031.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@34031.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@34031.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@34031.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@34031.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@34039.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@34039.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@34039.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@34039.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@34039.4]
  wire  x556_kernelx556_concrete1_clock; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_reset; // @[sm_x556.scala 102:24:@34068.4]
  wire [63:0] x556_kernelx556_concrete1_io_in_x276_outdram_number; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_in_x421_ready; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_in_x421_valid; // @[sm_x556.scala 102:24:@34068.4]
  wire [20:0] x556_kernelx556_concrete1_io_in_x280_outbuf_0_rPort_0_ofs_0; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_in_x280_outbuf_0_rPort_0_en_0; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_in_x280_outbuf_0_rPort_0_backpressure; // @[sm_x556.scala 102:24:@34068.4]
  wire [7:0] x556_kernelx556_concrete1_io_in_x280_outbuf_0_rPort_0_output_0; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_in_x420_ready; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_in_x420_valid; // @[sm_x556.scala 102:24:@34068.4]
  wire [7:0] x556_kernelx556_concrete1_io_in_x420_bits_wdata_0; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_in_x420_bits_wstrb; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_in_x279_TVALID; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_in_x279_TREADY; // @[sm_x556.scala 102:24:@34068.4]
  wire [255:0] x556_kernelx556_concrete1_io_in_x279_TDATA; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_in_x419_ready; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_in_x419_valid; // @[sm_x556.scala 102:24:@34068.4]
  wire [63:0] x556_kernelx556_concrete1_io_in_x419_bits_addr; // @[sm_x556.scala 102:24:@34068.4]
  wire [31:0] x556_kernelx556_concrete1_io_in_x419_bits_size; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_in_x278_TVALID; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_in_x278_TREADY; // @[sm_x556.scala 102:24:@34068.4]
  wire [255:0] x556_kernelx556_concrete1_io_in_x278_TDATA; // @[sm_x556.scala 102:24:@34068.4]
  wire [7:0] x556_kernelx556_concrete1_io_in_x278_TID; // @[sm_x556.scala 102:24:@34068.4]
  wire [7:0] x556_kernelx556_concrete1_io_in_x278_TDEST; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x556.scala 102:24:@34068.4]
  wire  x556_kernelx556_concrete1_io_rr; // @[sm_x556.scala 102:24:@34068.4]
  wire  _T_266; // @[package.scala 100:49:@33997.4]
  reg  _T_269; // @[package.scala 48:56:@33998.4]
  reg [31:0] _RAND_0;
  wire  _T_283; // @[package.scala 96:25:@34036.4 package.scala 96:25:@34037.4]
  wire  _T_289; // @[package.scala 96:25:@34044.4 package.scala 96:25:@34045.4]
  wire  _T_292; // @[SpatialBlocks.scala 138:93:@34047.4]
  x280_outbuf_0 x280_outbuf_0 ( // @[m_x280_outbuf_0.scala 27:17:@33906.4]
    .clock(x280_outbuf_0_clock),
    .reset(x280_outbuf_0_reset),
    .io_rPort_0_ofs_0(x280_outbuf_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x280_outbuf_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x280_outbuf_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x280_outbuf_0_io_rPort_0_output_0)
  );
  x556_sm x556_sm ( // @[sm_x556.scala 37:18:@33964.4]
    .clock(x556_sm_clock),
    .reset(x556_sm_reset),
    .io_enable(x556_sm_io_enable),
    .io_done(x556_sm_io_done),
    .io_ctrDone(x556_sm_io_ctrDone),
    .io_ctrInc(x556_sm_io_ctrInc),
    .io_parentAck(x556_sm_io_parentAck),
    .io_doneIn_0(x556_sm_io_doneIn_0),
    .io_doneIn_1(x556_sm_io_doneIn_1),
    .io_enableOut_0(x556_sm_io_enableOut_0),
    .io_enableOut_1(x556_sm_io_enableOut_1),
    .io_childAck_0(x556_sm_io_childAck_0),
    .io_childAck_1(x556_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@34031.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@34039.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x556_kernelx556_concrete1 x556_kernelx556_concrete1 ( // @[sm_x556.scala 102:24:@34068.4]
    .clock(x556_kernelx556_concrete1_clock),
    .reset(x556_kernelx556_concrete1_reset),
    .io_in_x276_outdram_number(x556_kernelx556_concrete1_io_in_x276_outdram_number),
    .io_in_x421_ready(x556_kernelx556_concrete1_io_in_x421_ready),
    .io_in_x421_valid(x556_kernelx556_concrete1_io_in_x421_valid),
    .io_in_x280_outbuf_0_rPort_0_ofs_0(x556_kernelx556_concrete1_io_in_x280_outbuf_0_rPort_0_ofs_0),
    .io_in_x280_outbuf_0_rPort_0_en_0(x556_kernelx556_concrete1_io_in_x280_outbuf_0_rPort_0_en_0),
    .io_in_x280_outbuf_0_rPort_0_backpressure(x556_kernelx556_concrete1_io_in_x280_outbuf_0_rPort_0_backpressure),
    .io_in_x280_outbuf_0_rPort_0_output_0(x556_kernelx556_concrete1_io_in_x280_outbuf_0_rPort_0_output_0),
    .io_in_x420_ready(x556_kernelx556_concrete1_io_in_x420_ready),
    .io_in_x420_valid(x556_kernelx556_concrete1_io_in_x420_valid),
    .io_in_x420_bits_wdata_0(x556_kernelx556_concrete1_io_in_x420_bits_wdata_0),
    .io_in_x420_bits_wstrb(x556_kernelx556_concrete1_io_in_x420_bits_wstrb),
    .io_in_x279_TVALID(x556_kernelx556_concrete1_io_in_x279_TVALID),
    .io_in_x279_TREADY(x556_kernelx556_concrete1_io_in_x279_TREADY),
    .io_in_x279_TDATA(x556_kernelx556_concrete1_io_in_x279_TDATA),
    .io_in_x419_ready(x556_kernelx556_concrete1_io_in_x419_ready),
    .io_in_x419_valid(x556_kernelx556_concrete1_io_in_x419_valid),
    .io_in_x419_bits_addr(x556_kernelx556_concrete1_io_in_x419_bits_addr),
    .io_in_x419_bits_size(x556_kernelx556_concrete1_io_in_x419_bits_size),
    .io_in_x278_TVALID(x556_kernelx556_concrete1_io_in_x278_TVALID),
    .io_in_x278_TREADY(x556_kernelx556_concrete1_io_in_x278_TREADY),
    .io_in_x278_TDATA(x556_kernelx556_concrete1_io_in_x278_TDATA),
    .io_in_x278_TID(x556_kernelx556_concrete1_io_in_x278_TID),
    .io_in_x278_TDEST(x556_kernelx556_concrete1_io_in_x278_TDEST),
    .io_sigsIn_smEnableOuts_0(x556_kernelx556_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x556_kernelx556_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x556_kernelx556_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x556_kernelx556_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x556_kernelx556_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x556_kernelx556_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(x556_kernelx556_concrete1_io_rr)
  );
  assign _T_266 = x556_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@33997.4]
  assign _T_283 = RetimeWrapper_io_out; // @[package.scala 96:25:@34036.4 package.scala 96:25:@34037.4]
  assign _T_289 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@34044.4 package.scala 96:25:@34045.4]
  assign _T_292 = ~ _T_289; // @[SpatialBlocks.scala 138:93:@34047.4]
  assign io_in_x421_ready = x556_kernelx556_concrete1_io_in_x421_ready; // @[sm_x556.scala 64:23:@34150.4]
  assign io_in_x420_valid = x556_kernelx556_concrete1_io_in_x420_valid; // @[sm_x556.scala 66:23:@34158.4]
  assign io_in_x420_bits_wdata_0 = x556_kernelx556_concrete1_io_in_x420_bits_wdata_0; // @[sm_x556.scala 66:23:@34157.4]
  assign io_in_x420_bits_wstrb = x556_kernelx556_concrete1_io_in_x420_bits_wstrb; // @[sm_x556.scala 66:23:@34156.4]
  assign io_in_x279_TVALID = x556_kernelx556_concrete1_io_in_x279_TVALID; // @[sm_x556.scala 67:23:@34168.4]
  assign io_in_x279_TDATA = x556_kernelx556_concrete1_io_in_x279_TDATA; // @[sm_x556.scala 67:23:@34166.4]
  assign io_in_x419_valid = x556_kernelx556_concrete1_io_in_x419_valid; // @[sm_x556.scala 68:23:@34171.4]
  assign io_in_x419_bits_addr = x556_kernelx556_concrete1_io_in_x419_bits_addr; // @[sm_x556.scala 68:23:@34170.4]
  assign io_in_x419_bits_size = x556_kernelx556_concrete1_io_in_x419_bits_size; // @[sm_x556.scala 68:23:@34169.4]
  assign io_in_x278_TREADY = x556_kernelx556_concrete1_io_in_x278_TREADY; // @[sm_x556.scala 69:23:@34180.4]
  assign io_sigsOut_smDoneIn_0 = x556_sm_io_done; // @[SpatialBlocks.scala 156:53:@34054.4]
  assign x280_outbuf_0_clock = clock; // @[:@33907.4]
  assign x280_outbuf_0_reset = reset; // @[:@33908.4]
  assign x280_outbuf_0_io_rPort_0_ofs_0 = x556_kernelx556_concrete1_io_in_x280_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@34154.4]
  assign x280_outbuf_0_io_rPort_0_en_0 = x556_kernelx556_concrete1_io_in_x280_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@34153.4]
  assign x280_outbuf_0_io_rPort_0_backpressure = x556_kernelx556_concrete1_io_in_x280_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@34152.4]
  assign x556_sm_clock = clock; // @[:@33965.4]
  assign x556_sm_reset = reset; // @[:@33966.4]
  assign x556_sm_io_enable = _T_283 & _T_292; // @[SpatialBlocks.scala 140:18:@34051.4]
  assign x556_sm_io_ctrDone = x556_sm_io_ctrInc & _T_269; // @[sm_RootController.scala 82:26:@34001.4]
  assign x556_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@34053.4]
  assign x556_sm_io_doneIn_0 = x556_kernelx556_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@34021.4]
  assign x556_sm_io_doneIn_1 = x556_kernelx556_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@34022.4]
  assign RetimeWrapper_clock = clock; // @[:@34032.4]
  assign RetimeWrapper_reset = reset; // @[:@34033.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@34035.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@34034.4]
  assign RetimeWrapper_1_clock = clock; // @[:@34040.4]
  assign RetimeWrapper_1_reset = reset; // @[:@34041.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@34043.4]
  assign RetimeWrapper_1_io_in = x556_sm_io_done; // @[package.scala 94:16:@34042.4]
  assign x556_kernelx556_concrete1_clock = clock; // @[:@34069.4]
  assign x556_kernelx556_concrete1_reset = reset; // @[:@34070.4]
  assign x556_kernelx556_concrete1_io_in_x276_outdram_number = io_in_x276_outdram_number; // @[sm_x556.scala 63:31:@34147.4]
  assign x556_kernelx556_concrete1_io_in_x421_valid = io_in_x421_valid; // @[sm_x556.scala 64:23:@34149.4]
  assign x556_kernelx556_concrete1_io_in_x280_outbuf_0_rPort_0_output_0 = x280_outbuf_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@34151.4]
  assign x556_kernelx556_concrete1_io_in_x420_ready = io_in_x420_ready; // @[sm_x556.scala 66:23:@34159.4]
  assign x556_kernelx556_concrete1_io_in_x279_TREADY = io_in_x279_TREADY; // @[sm_x556.scala 67:23:@34167.4]
  assign x556_kernelx556_concrete1_io_in_x419_ready = io_in_x419_ready; // @[sm_x556.scala 68:23:@34172.4]
  assign x556_kernelx556_concrete1_io_in_x278_TVALID = io_in_x278_TVALID; // @[sm_x556.scala 69:23:@34181.4]
  assign x556_kernelx556_concrete1_io_in_x278_TDATA = io_in_x278_TDATA; // @[sm_x556.scala 69:23:@34179.4]
  assign x556_kernelx556_concrete1_io_in_x278_TID = io_in_x278_TID; // @[sm_x556.scala 69:23:@34175.4]
  assign x556_kernelx556_concrete1_io_in_x278_TDEST = io_in_x278_TDEST; // @[sm_x556.scala 69:23:@34174.4]
  assign x556_kernelx556_concrete1_io_sigsIn_smEnableOuts_0 = x556_sm_io_enableOut_0; // @[sm_x556.scala 107:22:@34192.4]
  assign x556_kernelx556_concrete1_io_sigsIn_smEnableOuts_1 = x556_sm_io_enableOut_1; // @[sm_x556.scala 107:22:@34193.4]
  assign x556_kernelx556_concrete1_io_sigsIn_smChildAcks_0 = x556_sm_io_childAck_0; // @[sm_x556.scala 107:22:@34188.4]
  assign x556_kernelx556_concrete1_io_sigsIn_smChildAcks_1 = x556_sm_io_childAck_1; // @[sm_x556.scala 107:22:@34189.4]
  assign x556_kernelx556_concrete1_io_rr = io_rr; // @[sm_x556.scala 106:18:@34182.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_269 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_269 <= 1'h0;
    end else begin
      _T_269 <= _T_266;
    end
  end
endmodule
module AccelUnit( // @[:@34215.2]
  input          clock, // @[:@34216.4]
  input          reset, // @[:@34217.4]
  input          io_enable, // @[:@34218.4]
  output         io_done, // @[:@34218.4]
  input          io_reset, // @[:@34218.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@34218.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@34218.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@34218.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@34218.4]
  output         io_memStreams_loads_0_data_ready, // @[:@34218.4]
  input          io_memStreams_loads_0_data_valid, // @[:@34218.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@34218.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@34218.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@34218.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@34218.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@34218.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@34218.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@34218.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@34218.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@34218.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@34218.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@34218.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@34218.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@34218.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@34218.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@34218.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@34218.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@34218.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@34218.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@34218.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@34218.4]
  input          io_memStreams_stores_0_data_ready, // @[:@34218.4]
  output         io_memStreams_stores_0_data_valid, // @[:@34218.4]
  output [7:0]   io_memStreams_stores_0_data_bits_wdata_0, // @[:@34218.4]
  output         io_memStreams_stores_0_data_bits_wstrb, // @[:@34218.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@34218.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@34218.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@34218.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@34218.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@34218.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@34218.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@34218.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@34218.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@34218.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@34218.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@34218.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@34218.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@34218.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@34218.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@34218.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@34218.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@34218.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@34218.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@34218.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@34218.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@34218.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@34218.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@34218.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@34218.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@34218.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@34218.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@34218.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@34218.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@34218.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@34218.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@34218.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@34218.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@34218.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@34218.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@34218.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@34218.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@34218.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@34218.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@34218.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@34218.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@34218.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@34218.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@34218.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@34218.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@34218.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@34218.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@34218.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@34218.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@34218.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@34218.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@34218.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@34218.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@34218.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@34218.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@34218.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@34218.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@34218.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@34218.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@34218.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@34218.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@34218.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@34218.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@34218.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@34218.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@34218.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@34218.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@34218.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@34218.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@34218.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@34218.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@34218.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@34218.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@34218.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@34218.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@34218.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@34218.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@34218.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@34218.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@34218.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@34218.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@34218.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@34218.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@34218.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@34218.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@34218.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@34218.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@34218.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@34218.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@34218.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@34218.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@34218.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@34218.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@34218.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@34218.4]
  output         io_heap_0_req_valid, // @[:@34218.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@34218.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@34218.4]
  input          io_heap_0_resp_valid, // @[:@34218.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@34218.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@34218.4]
  input  [63:0]  io_argIns_0, // @[:@34218.4]
  input  [63:0]  io_argIns_1, // @[:@34218.4]
  input          io_argOuts_0_port_ready, // @[:@34218.4]
  output         io_argOuts_0_port_valid, // @[:@34218.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@34218.4]
  input  [63:0]  io_argOuts_0_echo // @[:@34218.4]
);
  wire  SingleCounter_clock; // @[Main.scala 40:32:@34366.4]
  wire  SingleCounter_reset; // @[Main.scala 40:32:@34366.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 40:32:@34366.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 40:32:@34366.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@34384.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@34384.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@34384.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@34384.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@34384.4]
  wire  SRFF_clock; // @[Main.scala 44:28:@34393.4]
  wire  SRFF_reset; // @[Main.scala 44:28:@34393.4]
  wire  SRFF_io_input_set; // @[Main.scala 44:28:@34393.4]
  wire  SRFF_io_input_reset; // @[Main.scala 44:28:@34393.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 44:28:@34393.4]
  wire  SRFF_io_output; // @[Main.scala 44:28:@34393.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 36:18:@34432.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 36:18:@34432.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 36:18:@34432.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 36:18:@34432.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 36:18:@34432.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 36:18:@34432.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 36:18:@34432.4]
  wire  RootController_sm_io_parentAck; // @[sm_RootController.scala 36:18:@34432.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 36:18:@34432.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 36:18:@34432.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 36:18:@34432.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@34464.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@34464.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@34464.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@34464.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@34464.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 91:24:@34526.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 91:24:@34526.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x276_outdram_number; // @[sm_RootController.scala 91:24:@34526.4]
  wire  RootController_kernelRootController_concrete1_io_in_x421_ready; // @[sm_RootController.scala 91:24:@34526.4]
  wire  RootController_kernelRootController_concrete1_io_in_x421_valid; // @[sm_RootController.scala 91:24:@34526.4]
  wire  RootController_kernelRootController_concrete1_io_in_x420_ready; // @[sm_RootController.scala 91:24:@34526.4]
  wire  RootController_kernelRootController_concrete1_io_in_x420_valid; // @[sm_RootController.scala 91:24:@34526.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x420_bits_wdata_0; // @[sm_RootController.scala 91:24:@34526.4]
  wire  RootController_kernelRootController_concrete1_io_in_x420_bits_wstrb; // @[sm_RootController.scala 91:24:@34526.4]
  wire  RootController_kernelRootController_concrete1_io_in_x279_TVALID; // @[sm_RootController.scala 91:24:@34526.4]
  wire  RootController_kernelRootController_concrete1_io_in_x279_TREADY; // @[sm_RootController.scala 91:24:@34526.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x279_TDATA; // @[sm_RootController.scala 91:24:@34526.4]
  wire  RootController_kernelRootController_concrete1_io_in_x419_ready; // @[sm_RootController.scala 91:24:@34526.4]
  wire  RootController_kernelRootController_concrete1_io_in_x419_valid; // @[sm_RootController.scala 91:24:@34526.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x419_bits_addr; // @[sm_RootController.scala 91:24:@34526.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x419_bits_size; // @[sm_RootController.scala 91:24:@34526.4]
  wire  RootController_kernelRootController_concrete1_io_in_x278_TVALID; // @[sm_RootController.scala 91:24:@34526.4]
  wire  RootController_kernelRootController_concrete1_io_in_x278_TREADY; // @[sm_RootController.scala 91:24:@34526.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x278_TDATA; // @[sm_RootController.scala 91:24:@34526.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x278_TID; // @[sm_RootController.scala 91:24:@34526.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x278_TDEST; // @[sm_RootController.scala 91:24:@34526.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 91:24:@34526.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 91:24:@34526.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 91:24:@34526.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 91:24:@34526.4]
  wire  _T_599; // @[package.scala 96:25:@34389.4 package.scala 96:25:@34390.4]
  wire  _T_664; // @[Main.scala 46:50:@34460.4]
  wire  _T_665; // @[Main.scala 46:59:@34461.4]
  wire  _T_677; // @[package.scala 100:49:@34481.4]
  reg  _T_680; // @[package.scala 48:56:@34482.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 40:32:@34366.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@34384.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 44:28:@34393.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 36:18:@34432.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_parentAck(RootController_sm_io_parentAck),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@34464.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 91:24:@34526.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x276_outdram_number(RootController_kernelRootController_concrete1_io_in_x276_outdram_number),
    .io_in_x421_ready(RootController_kernelRootController_concrete1_io_in_x421_ready),
    .io_in_x421_valid(RootController_kernelRootController_concrete1_io_in_x421_valid),
    .io_in_x420_ready(RootController_kernelRootController_concrete1_io_in_x420_ready),
    .io_in_x420_valid(RootController_kernelRootController_concrete1_io_in_x420_valid),
    .io_in_x420_bits_wdata_0(RootController_kernelRootController_concrete1_io_in_x420_bits_wdata_0),
    .io_in_x420_bits_wstrb(RootController_kernelRootController_concrete1_io_in_x420_bits_wstrb),
    .io_in_x279_TVALID(RootController_kernelRootController_concrete1_io_in_x279_TVALID),
    .io_in_x279_TREADY(RootController_kernelRootController_concrete1_io_in_x279_TREADY),
    .io_in_x279_TDATA(RootController_kernelRootController_concrete1_io_in_x279_TDATA),
    .io_in_x419_ready(RootController_kernelRootController_concrete1_io_in_x419_ready),
    .io_in_x419_valid(RootController_kernelRootController_concrete1_io_in_x419_valid),
    .io_in_x419_bits_addr(RootController_kernelRootController_concrete1_io_in_x419_bits_addr),
    .io_in_x419_bits_size(RootController_kernelRootController_concrete1_io_in_x419_bits_size),
    .io_in_x278_TVALID(RootController_kernelRootController_concrete1_io_in_x278_TVALID),
    .io_in_x278_TREADY(RootController_kernelRootController_concrete1_io_in_x278_TREADY),
    .io_in_x278_TDATA(RootController_kernelRootController_concrete1_io_in_x278_TDATA),
    .io_in_x278_TID(RootController_kernelRootController_concrete1_io_in_x278_TID),
    .io_in_x278_TDEST(RootController_kernelRootController_concrete1_io_in_x278_TDEST),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@34389.4 package.scala 96:25:@34390.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 46:50:@34460.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 46:59:@34461.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@34481.4]
  assign io_done = SRFF_io_output; // @[Main.scala 53:23:@34480.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x419_valid; // @[sm_RootController.scala 64:23:@34606.4]
  assign io_memStreams_stores_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x419_bits_addr; // @[sm_RootController.scala 64:23:@34605.4]
  assign io_memStreams_stores_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x419_bits_size; // @[sm_RootController.scala 64:23:@34604.4]
  assign io_memStreams_stores_0_data_valid = RootController_kernelRootController_concrete1_io_in_x420_valid; // @[sm_RootController.scala 62:23:@34593.4]
  assign io_memStreams_stores_0_data_bits_wdata_0 = RootController_kernelRootController_concrete1_io_in_x420_bits_wdata_0; // @[sm_RootController.scala 62:23:@34592.4]
  assign io_memStreams_stores_0_data_bits_wstrb = RootController_kernelRootController_concrete1_io_in_x420_bits_wstrb; // @[sm_RootController.scala 62:23:@34591.4]
  assign io_memStreams_stores_0_wresp_ready = RootController_kernelRootController_concrete1_io_in_x421_ready; // @[sm_RootController.scala 61:23:@34590.4]
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x278_TREADY; // @[sm_RootController.scala 65:23:@34615.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x279_TVALID; // @[sm_RootController.scala 63:23:@34603.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x279_TDATA; // @[sm_RootController.scala 63:23:@34601.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 63:23:@34600.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 63:23:@34599.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 63:23:@34598.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 63:23:@34597.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 63:23:@34596.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 63:23:@34595.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@34367.4]
  assign SingleCounter_reset = reset; // @[:@34368.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 41:79:@34382.4]
  assign RetimeWrapper_clock = clock; // @[:@34385.4]
  assign RetimeWrapper_reset = reset; // @[:@34386.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@34388.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@34387.4]
  assign SRFF_clock = clock; // @[:@34394.4]
  assign SRFF_reset = reset; // @[:@34395.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 62:29:@34644.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 51:31:@34478.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 52:36:@34479.4]
  assign RootController_sm_clock = clock; // @[:@34433.4]
  assign RootController_sm_reset = reset; // @[:@34434.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 50:33:@34477.4 SpatialBlocks.scala 140:18:@34511.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@34505.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 54:34:@34485.4]
  assign RootController_sm_io_parentAck = 1'h0; // @[Main.scala 49:36:@34473.4 SpatialBlocks.scala 142:21:@34513.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@34502.4]
  assign RetimeWrapper_1_clock = clock; // @[:@34465.4]
  assign RetimeWrapper_1_reset = reset; // @[:@34466.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@34468.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@34467.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@34527.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@34528.4]
  assign RootController_kernelRootController_concrete1_io_in_x276_outdram_number = io_argIns_1; // @[sm_RootController.scala 60:31:@34587.4]
  assign RootController_kernelRootController_concrete1_io_in_x421_valid = io_memStreams_stores_0_wresp_valid; // @[sm_RootController.scala 61:23:@34589.4]
  assign RootController_kernelRootController_concrete1_io_in_x420_ready = io_memStreams_stores_0_data_ready; // @[sm_RootController.scala 62:23:@34594.4]
  assign RootController_kernelRootController_concrete1_io_in_x279_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 63:23:@34602.4]
  assign RootController_kernelRootController_concrete1_io_in_x419_ready = io_memStreams_stores_0_cmd_ready; // @[sm_RootController.scala 64:23:@34607.4]
  assign RootController_kernelRootController_concrete1_io_in_x278_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 65:23:@34616.4]
  assign RootController_kernelRootController_concrete1_io_in_x278_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 65:23:@34614.4]
  assign RootController_kernelRootController_concrete1_io_in_x278_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 65:23:@34610.4]
  assign RootController_kernelRootController_concrete1_io_in_x278_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 65:23:@34609.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 96:22:@34625.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 96:22:@34623.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 95:18:@34617.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module SpatialIP( // @[:@34646.2]
  input         clock, // @[:@34647.4]
  input         reset, // @[:@34648.4]
  input  [31:0] io_raddr, // @[:@34649.4]
  input         io_wen, // @[:@34649.4]
  input  [31:0] io_waddr, // @[:@34649.4]
  input  [63:0] io_wdata, // @[:@34649.4]
  output [63:0] io_rdata // @[:@34649.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@34651.4]
  wire [7:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@34651.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@34651.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@34651.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@34651.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@34651.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@34651.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@34651.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@34651.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@34651.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@34651.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@34651.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  assign io_rdata = 64'h0;
  assign accel_clock = clock; // @[:@34652.4]
  assign accel_reset = reset; // @[:@34653.4]
  assign accel_io_enable = 1'h0;
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_loads_0_data_valid = 1'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0;
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0;
  assign accel_io_memStreams_stores_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_stores_0_data_ready = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_stores_0_wresp_bits = 1'h0;
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0;
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0;
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0;
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0;
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0;
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = 1'h0;
  assign accel_io_heap_0_resp_bits_allocDealloc = 1'h0;
  assign accel_io_heap_0_resp_bits_sizeAddr = 64'h0;
  assign accel_io_argIns_0 = 64'h0;
  assign accel_io_argIns_1 = 64'h0;
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0;
endmodule
