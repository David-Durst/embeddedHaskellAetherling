module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  output [31:0] O_0,
  output [31:0] O_1
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(clock), // @[:@1296.4]
    .reset(reset), // @[:@1297.4]
    .io_in_x250_TREADY(dontcare), // @[:@1298.4]
    .io_in_x250_TDATA({I_0,I_1}), // @[:@1298.4]
    .io_in_x250_TID(8'h0),
    .io_in_x250_TDEST(8'h0),
    .io_in_x251_TVALID(valid_down), // @[:@1298.4]
    .io_in_x251_TDATA({O_0,O_1}), // @[:@1298.4]
    .io_in_x251_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x258_ctrchain cchain ( // @[:@2879.2]
    .clock(clock), // @[:@2880.4]
    .reset(reset), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule


module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 321:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 325:12:@24.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : io_wPort_0_data_0; // @[MemPrimitives.scala 325:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        ff <= io_wPort_0_data_0;
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh30); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh30); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_parentAck, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  _T_81; // @[Controllers.scala 86:43:@328.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_93; // @[Controllers.scala 92:52:@342.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_134; // @[Controllers.scala 129:57:@382.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  wire  _T_167; // @[package.scala 100:41:@414.4]
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign _T_81 = io_rst | done_0_io_output; // @[Controllers.scala 86:43:@328.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_93 = synchronize | io_rst; // @[Controllers.scala 92:52:@342.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_134 = _T_133 | io_parentAck; // @[Controllers.scala 129:57:@382.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign _T_167 = done_0_io_output & _T_166; // @[package.scala 100:41:@414.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_134 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = _T_81 | io_parentAck; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = _T_93 | io_parentAck; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = _T_167 | io_parentAck; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module SRAM( // @[:@507.2]
  input         clock, // @[:@508.4]
  input  [20:0] io_raddr, // @[:@510.4]
  output [31:0] io_rdata, // @[:@510.4]
  input         io_backpressure // @[:@510.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@512.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@512.4]
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(2073600), .AWIDTH(21)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@512.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign io_rdata = SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@539.4]
  assign SRAMVerilogAWS_wdata = 32'h0; // @[SRAM.scala 175:20:@526.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@527.4]
  assign SRAMVerilogAWS_wen = 1'h0; // @[SRAM.scala 173:18:@524.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@529.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@528.4]
  assign SRAMVerilogAWS_waddr = 21'h0; // @[SRAM.scala 174:20:@525.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@523.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@522.4]
endmodule
module RetimeWrapper_5( // @[:@553.2]
  input         clock, // @[:@554.4]
  input         reset, // @[:@555.4]
  input         io_flow, // @[:@556.4]
  input  [20:0] io_in, // @[:@556.4]
  output [20:0] io_out // @[:@556.4]
);
  wire [20:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@558.4]
  RetimeShiftRegister #(.WIDTH(21), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@558.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@571.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@570.4]
  assign sr_init = 21'h0; // @[RetimeShiftRegister.scala 19:16:@569.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@568.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@567.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@565.4]
endmodule
module Mem1D( // @[:@573.2]
  input         clock, // @[:@574.4]
  input         reset, // @[:@575.4]
  input  [20:0] io_r_ofs_0, // @[:@576.4]
  input         io_r_backpressure, // @[:@576.4]
  output [31:0] io_output // @[:@576.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@580.4]
  wire [20:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@580.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@580.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@580.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_in; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_out; // @[package.scala 93:22:@583.4]
  SRAM SRAM ( // @[MemPrimitives.scala 715:21:@580.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@583.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@596.4]
  assign SRAM_clock = clock; // @[:@581.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@590.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@595.4]
  assign RetimeWrapper_clock = clock; // @[:@584.4]
  assign RetimeWrapper_reset = reset; // @[:@585.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@587.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@586.4]
endmodule
module StickySelects( // @[:@598.2]
  input   io_ins_0, // @[:@601.4]
  output  io_outs_0 // @[:@601.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 34:26:@603.4]
endmodule
module RetimeWrapper_6( // @[:@617.2]
  input   clock, // @[:@618.4]
  input   reset, // @[:@619.4]
  input   io_flow, // @[:@620.4]
  input   io_in, // @[:@620.4]
  output  io_out // @[:@620.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@622.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@622.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@635.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@634.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@633.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@632.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@631.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@629.4]
endmodule
module x252_outbuf_0( // @[:@637.2]
  input         clock, // @[:@638.4]
  input         reset, // @[:@639.4]
  input  [20:0] io_rPort_0_ofs_0, // @[:@640.4]
  input         io_rPort_0_en_0, // @[:@640.4]
  input         io_rPort_0_backpressure, // @[:@640.4]
  output [31:0] io_rPort_0_output_0 // @[:@640.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@655.4]
  wire [20:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@655.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@655.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@695.4]
  wire  _T_76; // @[MemPrimitives.scala 126:35:@685.4]
  wire [22:0] _T_78; // @[Cat.scala 30:58:@687.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@655.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@681.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@695.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@685.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@687.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@702.4]
  assign Mem1D_clock = clock; // @[:@656.4]
  assign Mem1D_reset = reset; // @[:@657.4]
  assign Mem1D_io_r_ofs_0 = _T_78[20:0]; // @[MemPrimitives.scala 131:28:@691.4]
  assign Mem1D_io_r_backpressure = _T_78[21]; // @[MemPrimitives.scala 132:32:@692.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@684.4]
  assign RetimeWrapper_clock = clock; // @[:@696.4]
  assign RetimeWrapper_reset = reset; // @[:@697.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@699.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@698.4]
endmodule
module x538_sm( // @[:@846.2]
  input   clock, // @[:@847.4]
  input   reset, // @[:@848.4]
  input   io_enable, // @[:@849.4]
  output  io_done, // @[:@849.4]
  input   io_ctrDone, // @[:@849.4]
  output  io_ctrInc, // @[:@849.4]
  input   io_parentAck, // @[:@849.4]
  input   io_doneIn_0, // @[:@849.4]
  input   io_doneIn_1, // @[:@849.4]
  output  io_enableOut_0, // @[:@849.4]
  output  io_enableOut_1, // @[:@849.4]
  output  io_childAck_0, // @[:@849.4]
  output  io_childAck_1 // @[:@849.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@852.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@855.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@858.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@861.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@893.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1011.4]
  wire  allDone; // @[Controllers.scala 80:47:@864.4]
  wire  synchronize; // @[Controllers.scala 146:56:@918.4]
  wire  _T_127; // @[Controllers.scala 150:35:@920.4]
  wire  _T_129; // @[Controllers.scala 150:60:@921.4]
  wire  _T_130; // @[Controllers.scala 150:58:@922.4]
  wire  _T_132; // @[Controllers.scala 150:76:@923.4]
  wire  _T_133; // @[Controllers.scala 150:74:@924.4]
  wire  _T_135; // @[Controllers.scala 150:97:@925.4]
  wire  _T_136; // @[Controllers.scala 150:95:@926.4]
  wire  _T_152; // @[Controllers.scala 150:35:@944.4]
  wire  _T_154; // @[Controllers.scala 150:60:@945.4]
  wire  _T_155; // @[Controllers.scala 150:58:@946.4]
  wire  _T_157; // @[Controllers.scala 150:76:@947.4]
  wire  _T_158; // @[Controllers.scala 150:74:@948.4]
  wire  _T_161; // @[Controllers.scala 150:95:@950.4]
  wire  _T_179; // @[Controllers.scala 213:68:@972.4]
  wire  _T_181; // @[Controllers.scala 213:90:@974.4]
  wire  _T_183; // @[Controllers.scala 213:132:@976.4]
  wire  _T_184; // @[Controllers.scala 213:130:@977.4]
  wire  _T_185; // @[Controllers.scala 213:156:@978.4]
  wire  _T_187; // @[Controllers.scala 213:68:@981.4]
  wire  _T_189; // @[Controllers.scala 213:90:@983.4]
  wire  _T_196; // @[package.scala 100:49:@989.4]
  reg  _T_199; // @[package.scala 48:56:@990.4]
  reg [31:0] _RAND_0;
  wire  _T_200; // @[package.scala 100:41:@992.4]
  reg  _T_213; // @[package.scala 48:56:@1008.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@852.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@855.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@858.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@861.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@890.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@893.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@994.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1011.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@864.4]
  assign synchronize = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 146:56:@918.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 150:35:@920.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 150:60:@921.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 150:58:@922.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 150:76:@923.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 150:74:@924.4]
  assign _T_135 = io_ctrDone == 1'h0; // @[Controllers.scala 150:97:@925.4]
  assign _T_136 = _T_133 & _T_135; // @[Controllers.scala 150:95:@926.4]
  assign _T_152 = ~ iterDone_1_io_output; // @[Controllers.scala 150:35:@944.4]
  assign _T_154 = io_doneIn_1 == 1'h0; // @[Controllers.scala 150:60:@945.4]
  assign _T_155 = _T_152 & _T_154; // @[Controllers.scala 150:58:@946.4]
  assign _T_157 = done_1_io_output == 1'h0; // @[Controllers.scala 150:76:@947.4]
  assign _T_158 = _T_155 & _T_157; // @[Controllers.scala 150:74:@948.4]
  assign _T_161 = _T_158 & _T_135; // @[Controllers.scala 150:95:@950.4]
  assign _T_179 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@972.4]
  assign _T_181 = _T_179 & _T_127; // @[Controllers.scala 213:90:@974.4]
  assign _T_183 = ~ allDone; // @[Controllers.scala 213:132:@976.4]
  assign _T_184 = _T_181 & _T_183; // @[Controllers.scala 213:130:@977.4]
  assign _T_185 = ~ io_ctrDone; // @[Controllers.scala 213:156:@978.4]
  assign _T_187 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@981.4]
  assign _T_189 = _T_187 & _T_152; // @[Controllers.scala 213:90:@983.4]
  assign _T_196 = allDone == 1'h0; // @[package.scala 100:49:@989.4]
  assign _T_200 = allDone & _T_199; // @[package.scala 100:41:@992.4]
  assign io_done = RetimeWrapper_1_io_out; // @[Controllers.scala 245:13:@1018.4]
  assign io_ctrInc = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 143:17:@917.4]
  assign io_enableOut_0 = _T_184 & _T_185; // @[Controllers.scala 213:55:@980.4]
  assign io_enableOut_1 = _T_189 & _T_183; // @[Controllers.scala 213:55:@988.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@969.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@971.4]
  assign active_0_clock = clock; // @[:@853.4]
  assign active_0_reset = reset; // @[:@854.4]
  assign active_0_io_input_set = _T_136 & io_enable; // @[Controllers.scala 150:32:@929.4]
  assign active_0_io_input_reset = io_doneIn_0 | io_parentAck; // @[Controllers.scala 151:34:@933.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@867.4]
  assign active_1_clock = clock; // @[:@856.4]
  assign active_1_reset = reset; // @[:@857.4]
  assign active_1_io_input_set = _T_161 & io_enable; // @[Controllers.scala 150:32:@953.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_parentAck; // @[Controllers.scala 151:34:@957.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@868.4]
  assign done_0_clock = clock; // @[:@859.4]
  assign done_0_reset = reset; // @[:@860.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@943.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@879.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@869.4]
  assign done_1_clock = clock; // @[:@862.4]
  assign done_1_reset = reset; // @[:@863.4]
  assign done_1_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@967.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@888.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@870.4]
  assign iterDone_0_clock = clock; // @[:@891.4]
  assign iterDone_0_reset = reset; // @[:@892.4]
  assign iterDone_0_io_input_set = io_doneIn_0; // @[Controllers.scala 152:34:@939.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@906.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@896.4]
  assign iterDone_1_clock = clock; // @[:@894.4]
  assign iterDone_1_reset = reset; // @[:@895.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 152:34:@963.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@915.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@897.4]
  assign RetimeWrapper_clock = clock; // @[:@995.4]
  assign RetimeWrapper_reset = reset; // @[:@996.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@998.4]
  assign RetimeWrapper_io_in = _T_200 | io_parentAck; // @[package.scala 94:16:@997.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1012.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1013.4]
  assign RetimeWrapper_1_io_flow = io_enable; // @[package.scala 95:18:@1015.4]
  assign RetimeWrapper_1_io_in = allDone & _T_213; // @[package.scala 94:16:@1014.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_199 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_213 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_199 <= 1'h0;
    end else begin
      _T_199 <= _T_196;
    end
    if (reset) begin
      _T_213 <= 1'h0;
    end else begin
      _T_213 <= _T_196;
    end
  end
endmodule
module x467_outr_UnitPipe_sm( // @[:@1435.2]
  input   clock, // @[:@1436.4]
  input   reset, // @[:@1437.4]
  input   io_enable, // @[:@1438.4]
  output  io_done, // @[:@1438.4]
  input   io_parentAck, // @[:@1438.4]
  input   io_doneIn_0, // @[:@1438.4]
  input   io_doneIn_1, // @[:@1438.4]
  output  io_enableOut_0, // @[:@1438.4]
  output  io_enableOut_1, // @[:@1438.4]
  output  io_childAck_0, // @[:@1438.4]
  output  io_childAck_1, // @[:@1438.4]
  input   io_ctrCopyDone_0, // @[:@1438.4]
  input   io_ctrCopyDone_1 // @[:@1438.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@1441.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@1444.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@1447.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1450.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1482.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1688.4]
  wire  allDone; // @[Controllers.scala 80:47:@1453.4]
  wire  _T_127; // @[Controllers.scala 165:35:@1507.4]
  wire  _T_129; // @[Controllers.scala 165:60:@1508.4]
  wire  _T_130; // @[Controllers.scala 165:58:@1509.4]
  wire  _T_132; // @[Controllers.scala 165:76:@1510.4]
  wire  _T_133; // @[Controllers.scala 165:74:@1511.4]
  wire  _T_137; // @[Controllers.scala 165:109:@1514.4]
  wire  _T_140; // @[Controllers.scala 165:141:@1516.4]
  wire  _T_148; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  wire  _T_152; // @[Controllers.scala 167:54:@1531.4]
  wire  _T_153; // @[Controllers.scala 167:52:@1532.4]
  wire  _T_160; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  wire  _T_178; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  wire  _T_182; // @[Controllers.scala 169:67:@1563.4]
  wire  _T_183; // @[Controllers.scala 169:86:@1564.4]
  wire  _T_195; // @[Controllers.scala 165:35:@1576.4]
  wire  _T_197; // @[Controllers.scala 165:60:@1577.4]
  wire  _T_198; // @[Controllers.scala 165:58:@1578.4]
  wire  _T_200; // @[Controllers.scala 165:76:@1579.4]
  wire  _T_201; // @[Controllers.scala 165:74:@1580.4]
  wire  _T_205; // @[Controllers.scala 165:109:@1583.4]
  wire  _T_208; // @[Controllers.scala 165:141:@1585.4]
  wire  _T_216; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  wire  _T_220; // @[Controllers.scala 167:54:@1600.4]
  wire  _T_221; // @[Controllers.scala 167:52:@1601.4]
  wire  _T_228; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  wire  _T_246; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  wire  _T_250; // @[Controllers.scala 169:67:@1632.4]
  wire  _T_251; // @[Controllers.scala 169:86:@1633.4]
  wire  _T_265; // @[Controllers.scala 213:68:@1649.4]
  wire  _T_267; // @[Controllers.scala 213:90:@1651.4]
  wire  _T_269; // @[Controllers.scala 213:132:@1653.4]
  wire  _T_273; // @[Controllers.scala 213:68:@1658.4]
  wire  _T_275; // @[Controllers.scala 213:90:@1660.4]
  wire  _T_282; // @[package.scala 100:49:@1666.4]
  reg  _T_285; // @[package.scala 48:56:@1667.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@1669.4]
  reg  _T_299; // @[package.scala 48:56:@1685.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@1441.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@1444.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@1447.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1450.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1479.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1482.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1523.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1537.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1555.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1592.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1606.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1624.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1671.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1688.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1453.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1507.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1508.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@1509.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1510.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@1511.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@1514.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1516.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@1531.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@1532.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@1563.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@1564.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1576.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1577.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@1578.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1579.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@1580.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@1583.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1585.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@1600.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@1601.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@1632.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@1633.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1649.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@1651.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@1653.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1658.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@1660.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@1666.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@1669.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@1695.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@1657.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@1665.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1646.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1648.4]
  assign active_0_clock = clock; // @[:@1442.4]
  assign active_0_reset = reset; // @[:@1443.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@1518.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1522.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1456.4]
  assign active_1_clock = clock; // @[:@1445.4]
  assign active_1_reset = reset; // @[:@1446.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@1587.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1591.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1457.4]
  assign done_0_clock = clock; // @[:@1448.4]
  assign done_0_reset = reset; // @[:@1449.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@1568.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1468.4 Controllers.scala 170:32:@1575.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1458.4]
  assign done_1_clock = clock; // @[:@1451.4]
  assign done_1_reset = reset; // @[:@1452.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@1637.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1477.4 Controllers.scala 170:32:@1644.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1459.4]
  assign iterDone_0_clock = clock; // @[:@1480.4]
  assign iterDone_0_reset = reset; // @[:@1481.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@1536.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@1495.4 Controllers.scala 168:36:@1552.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1485.4]
  assign iterDone_1_clock = clock; // @[:@1483.4]
  assign iterDone_1_reset = reset; // @[:@1484.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@1605.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@1504.4 Controllers.scala 168:36:@1621.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1486.4]
  assign RetimeWrapper_clock = clock; // @[:@1524.4]
  assign RetimeWrapper_reset = reset; // @[:@1525.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1527.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1526.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1538.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1539.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1541.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1540.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1556.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1557.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1559.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1558.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1593.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1594.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1596.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1595.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1607.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1608.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1610.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1609.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1625.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1626.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1628.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1627.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1672.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1673.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1675.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@1674.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1689.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1690.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@1692.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@1691.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module CompactingIncDincCtr( // @[:@1924.2]
  input   clock, // @[:@1925.4]
  input   reset, // @[:@1926.4]
  input   io_input_inc_en_0, // @[:@1927.4]
  input   io_input_dinc_en_0, // @[:@1927.4]
  output  io_output_full // @[:@1927.4]
);
  reg [31:0] cnt; // @[Counter.scala 170:20:@1929.4]
  reg [31:0] _RAND_0;
  wire [14:0] numPushed; // @[Counter.scala 172:47:@1930.4]
  wire [14:0] numPopped; // @[Counter.scala 173:48:@1931.4]
  wire [31:0] _GEN_0; // @[Counter.scala 174:14:@1932.4]
  wire [32:0] _T_37; // @[Counter.scala 174:14:@1932.4]
  wire [31:0] _T_38; // @[Counter.scala 174:14:@1933.4]
  wire [31:0] _T_39; // @[Counter.scala 174:14:@1934.4]
  wire [31:0] _GEN_1; // @[Counter.scala 174:26:@1935.4]
  wire [32:0] _T_40; // @[Counter.scala 174:26:@1935.4]
  wire [31:0] _T_41; // @[Counter.scala 174:26:@1936.4]
  wire [31:0] _T_42; // @[Counter.scala 174:26:@1937.4]
  assign numPushed = io_input_inc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 172:47:@1930.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 173:48:@1931.4]
  assign _GEN_0 = {{17{numPushed[14]}},numPushed}; // @[Counter.scala 174:14:@1932.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1932.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1933.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 174:14:@1934.4]
  assign _GEN_1 = {{17{numPopped[14]}},numPopped}; // @[Counter.scala 174:26:@1935.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1935.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1936.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 174:26:@1937.4]
  assign io_output_full = $signed(cnt) > $signed(32'sh1dff); // @[Counter.scala 180:18:@1951.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module x253_fifoinraw_0( // @[:@2074.2]
  input   clock, // @[:@2075.4]
  input   reset // @[:@2076.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2121.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2121.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign elements_clock = clock; // @[:@2122.4]
  assign elements_reset = reset; // @[:@2123.4]
  assign elements_io_input_inc_en_0 = 1'h0; // @[MemPrimitives.scala 394:79:@2133.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2134.4]
endmodule
module x254_fifoinpacked_0( // @[:@2497.2]
  input   clock, // @[:@2498.4]
  input   reset, // @[:@2499.4]
  input   io_wPort_0_en_0, // @[:@2500.4]
  output  io_full, // @[:@2500.4]
  input   io_active_0_in, // @[:@2500.4]
  output  io_active_0_out // @[:@2500.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2544.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2544.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 439:39:@2618.4]
  assign io_active_0_out = io_active_0_in; // @[MemPrimitives.scala 437:129:@2616.4]
  assign elements_clock = clock; // @[:@2545.4]
  assign elements_reset = reset; // @[:@2546.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 394:79:@2556.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2557.4]
endmodule
module FF_7( // @[:@3047.2]
  input         clock, // @[:@3048.4]
  input         reset, // @[:@3049.4]
  output [12:0] io_rPort_0_output_0, // @[:@3050.4]
  input  [12:0] io_wPort_0_data_0, // @[:@3050.4]
  input         io_wPort_0_reset, // @[:@3050.4]
  input         io_wPort_0_en_0 // @[:@3050.4]
);
  reg [12:0] ff; // @[MemPrimitives.scala 321:19:@3065.4]
  reg [31:0] _RAND_0;
  wire [12:0] _T_68; // @[MemPrimitives.scala 325:32:@3067.4]
  wire [12:0] _T_69; // @[MemPrimitives.scala 325:12:@3068.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@3067.4]
  assign _T_69 = io_wPort_0_reset ? 13'h0 : _T_68; // @[MemPrimitives.scala 325:12:@3068.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@3070.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 13'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 13'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_1( // @[:@3085.2]
  input         clock, // @[:@3086.4]
  input         reset, // @[:@3087.4]
  input         io_setup_saturate, // @[:@3088.4]
  input         io_input_reset, // @[:@3088.4]
  input         io_input_enable, // @[:@3088.4]
  output [12:0] io_output_count_0, // @[:@3088.4]
  output        io_output_oobs_0, // @[:@3088.4]
  output        io_output_done, // @[:@3088.4]
  output        io_output_saturated // @[:@3088.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3101.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3117.4]
  wire  _T_36; // @[Counter.scala 264:45:@3120.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3145.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3146.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3147.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3148.4]
  wire  _T_57; // @[Counter.scala 293:18:@3150.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3158.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3160.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3161.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3162.4]
  wire  _T_75; // @[Counter.scala 322:102:@3166.4]
  wire  _T_77; // @[Counter.scala 322:130:@3167.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3101.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3117.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3120.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3145.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3146.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3147.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3148.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh438); // @[Counter.scala 293:18:@3150.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3158.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3160.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3161.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3162.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3166.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh438); // @[Counter.scala 322:130:@3167.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3165.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3169.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3171.4]
  assign io_output_saturated = io_setup_saturate & _T_57; // @[Counter.scala 340:25:@3174.4]
  assign bases_0_clock = clock; // @[:@3102.4]
  assign bases_0_reset = reset; // @[:@3103.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3164.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3143.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3144.4]
  assign SRFF_clock = clock; // @[:@3118.4]
  assign SRFF_reset = reset; // @[:@3119.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3122.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3124.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3125.4]
endmodule
module SingleCounter_2( // @[:@3214.2]
  input         clock, // @[:@3215.4]
  input         reset, // @[:@3216.4]
  input         io_setup_saturate, // @[:@3217.4]
  input         io_input_reset, // @[:@3217.4]
  input         io_input_enable, // @[:@3217.4]
  output [12:0] io_output_count_0, // @[:@3217.4]
  output        io_output_oobs_0, // @[:@3217.4]
  output        io_output_done // @[:@3217.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3230.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3246.4]
  wire  _T_36; // @[Counter.scala 264:45:@3249.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3274.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3275.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3276.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3277.4]
  wire  _T_57; // @[Counter.scala 293:18:@3279.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3287.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3289.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3290.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3291.4]
  wire  _T_75; // @[Counter.scala 322:102:@3295.4]
  wire  _T_77; // @[Counter.scala 322:130:@3296.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3230.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3246.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3249.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3274.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh2); // @[Counter.scala 291:33:@3275.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh2); // @[Counter.scala 291:33:@3276.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3277.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh780); // @[Counter.scala 293:18:@3279.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3287.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3289.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3290.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3291.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3295.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh780); // @[Counter.scala 322:130:@3296.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3294.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3298.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3300.4]
  assign bases_0_clock = clock; // @[:@3231.4]
  assign bases_0_reset = reset; // @[:@3232.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3293.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3272.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3273.4]
  assign SRFF_clock = clock; // @[:@3247.4]
  assign SRFF_reset = reset; // @[:@3248.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3251.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3253.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3254.4]
endmodule
module x258_ctrchain( // @[:@3305.2]
  input         clock, // @[:@3306.4]
  input         reset, // @[:@3307.4]
  input         io_input_reset, // @[:@3308.4]
  input         io_input_enable, // @[:@3308.4]
  output [12:0] io_output_counts_1, // @[:@3308.4]
  output [12:0] io_output_counts_0, // @[:@3308.4]
  output        io_output_oobs_0, // @[:@3308.4]
  output        io_output_oobs_1, // @[:@3308.4]
  output        io_output_done // @[:@3308.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@3310.4]
  wire [12:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@3313.4]
  wire [12:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@3313.4]
  wire  isDone; // @[Counter.scala 541:51:@3330.4]
  reg  wasDone; // @[Counter.scala 542:24:@3331.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@3339.4]
  wire  _T_66; // @[Counter.scala 546:80:@3340.4]
  reg  doneLatch; // @[Counter.scala 550:26:@3345.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@3346.4]
  wire  _T_74; // @[Counter.scala 551:19:@3347.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@3310.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@3313.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@3330.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@3339.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@3340.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@3346.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@3347.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@3352.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@3349.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3351.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3354.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@3342.4]
  assign ctrs_0_clock = clock; // @[:@3311.4]
  assign ctrs_0_reset = reset; // @[:@3312.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 530:29:@3327.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3319.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@3326.4]
  assign ctrs_1_clock = clock; // @[:@3314.4]
  assign ctrs_1_reset = reset; // @[:@3315.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@3329.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3323.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@3324.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_21( // @[:@3394.2]
  input   clock, // @[:@3395.4]
  input   reset, // @[:@3396.4]
  input   io_flow, // @[:@3397.4]
  input   io_in, // @[:@3397.4]
  output  io_out // @[:@3397.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@3399.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3412.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3411.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3410.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3409.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3408.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3406.4]
endmodule
module RetimeWrapper_25( // @[:@3522.2]
  input   clock, // @[:@3523.4]
  input   reset, // @[:@3524.4]
  input   io_flow, // @[:@3525.4]
  input   io_in, // @[:@3525.4]
  output  io_out // @[:@3525.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@3527.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3540.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3539.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3538.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3537.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3536.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3534.4]
endmodule
module x274_inr_Foreach_sm( // @[:@3542.2]
  input   clock, // @[:@3543.4]
  input   reset, // @[:@3544.4]
  input   io_enable, // @[:@3545.4]
  output  io_done, // @[:@3545.4]
  output  io_doneLatch, // @[:@3545.4]
  input   io_ctrDone, // @[:@3545.4]
  output  io_datapathEn, // @[:@3545.4]
  output  io_ctrInc, // @[:@3545.4]
  output  io_ctrRst, // @[:@3545.4]
  input   io_parentAck, // @[:@3545.4]
  input   io_backpressure, // @[:@3545.4]
  input   io_break // @[:@3545.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3547.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3547.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3550.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3550.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3642.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3555.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3556.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3557.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3558.4]
  wire  _T_100; // @[package.scala 100:49:@3575.4]
  reg  _T_103; // @[package.scala 48:56:@3576.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  wire  _T_110; // @[package.scala 100:49:@3591.4]
  reg  _T_113; // @[package.scala 48:56:@3592.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3594.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3599.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3600.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3603.4]
  wire  _T_124; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  wire  _T_126; // @[package.scala 100:49:@3613.4]
  reg  _T_129; // @[package.scala 48:56:@3614.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3636.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3638.4]
  reg  _T_153; // @[package.scala 48:56:@3639.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3649.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3650.4]
  SRFF active ( // @[Controllers.scala 261:22:@3547.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3550.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@3584.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3606.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3618.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3626.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@3642.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3555.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3556.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3557.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3558.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3575.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3591.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3594.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3599.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3600.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3603.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3613.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3638.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3649.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3650.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3617.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3652.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3602.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3605.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3597.4]
  assign active_clock = clock; // @[:@3548.4]
  assign active_reset = reset; // @[:@3549.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3560.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3564.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3565.4]
  assign done_clock = clock; // @[:@3551.4]
  assign done_reset = reset; // @[:@3552.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3580.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3573.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3574.4]
  assign RetimeWrapper_clock = clock; // @[:@3585.4]
  assign RetimeWrapper_reset = reset; // @[:@3586.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3588.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3587.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3607.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3608.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3610.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3609.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3619.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3620.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3622.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3621.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3627.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3628.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3630.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3629.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3643.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3644.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3646.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3645.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module fix2fixBox( // @[:@3759.2]
  input  [31:0] io_a, // @[:@3762.4]
  output [31:0] io_b // @[:@3762.4]
);
  assign io_b = io_a; // @[Converter.scala 95:38:@3775.4]
endmodule
module _( // @[:@3777.2]
  input  [31:0] io_b, // @[:@3780.4]
  output [31:0] io_result // @[:@3780.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3785.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3785.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@3785.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3793.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3788.4]
endmodule
module fix2fixBox_2( // @[:@3831.2]
  input  [31:0] io_a, // @[:@3834.4]
  output [32:0] io_b // @[:@3834.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@3844.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@3844.4]
  assign io_b = {_T_20,io_a}; // @[Converter.scala 95:38:@3849.4]
endmodule
module __2( // @[:@3851.2]
  input  [31:0] io_b, // @[:@3854.4]
  output [32:0] io_result // @[:@3854.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3859.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3859.4]
  fix2fixBox_2 fix2fixBox ( // @[BigIPZynq.scala 219:30:@3859.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3867.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3862.4]
endmodule
module RetimeWrapper_29( // @[:@3919.2]
  input         clock, // @[:@3920.4]
  input         reset, // @[:@3921.4]
  input         io_flow, // @[:@3922.4]
  input  [31:0] io_in, // @[:@3922.4]
  output [31:0] io_out // @[:@3922.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3924.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3937.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3936.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3935.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3934.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3933.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3931.4]
endmodule
module fix2fixBox_4( // @[:@3939.2]
  input         clock, // @[:@3940.4]
  input         reset, // @[:@3941.4]
  input  [32:0] io_a, // @[:@3942.4]
  input         io_flow, // @[:@3942.4]
  output [31:0] io_b // @[:@3942.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3955.4]
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@3955.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@3962.4]
  assign RetimeWrapper_clock = clock; // @[:@3956.4]
  assign RetimeWrapper_reset = reset; // @[:@3957.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@3959.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@3958.4]
endmodule
module x516_sub( // @[:@3964.2]
  input         clock, // @[:@3965.4]
  input         reset, // @[:@3966.4]
  input  [31:0] io_a, // @[:@3967.4]
  input  [31:0] io_b, // @[:@3967.4]
  input         io_flow, // @[:@3967.4]
  output [31:0] io_result // @[:@3967.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@3975.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@3975.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@3982.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@3982.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@4001.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@4001.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@4001.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@3989.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@3990.4]
  __2 _ ( // @[Math.scala 720:24:@3975.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@3982.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 182:30:@4001.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@3989.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@3990.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@4009.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@3978.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@3985.4]
  assign fix2fixBox_clock = clock; // @[:@4002.4]
  assign fix2fixBox_reset = reset; // @[:@4003.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@4004.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@4007.4]
endmodule
module x264_sum( // @[:@4176.2]
  input         clock, // @[:@4177.4]
  input         reset, // @[:@4178.4]
  input  [31:0] io_a, // @[:@4179.4]
  input  [31:0] io_b, // @[:@4179.4]
  input         io_flow, // @[:@4179.4]
  output [31:0] io_result // @[:@4179.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4187.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@4187.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@4194.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@4194.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4212.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4212.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4212.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@4201.4]
  __2 _ ( // @[Math.scala 720:24:@4187.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@4194.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@4212.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4201.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4220.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@4190.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@4197.4]
  assign fix2fixBox_clock = clock; // @[:@4213.4]
  assign fix2fixBox_reset = reset; // @[:@4214.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4215.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4218.4]
endmodule
module x274_inr_Foreach_kernelx274_inr_Foreach_concrete1( // @[:@4748.2]
  input         clock, // @[:@4749.4]
  input         reset, // @[:@4750.4]
  output        io_in_x254_fifoinpacked_0_wPort_0_en_0, // @[:@4751.4]
  input         io_in_x254_fifoinpacked_0_full, // @[:@4751.4]
  output        io_in_x254_fifoinpacked_0_active_0_in, // @[:@4751.4]
  input         io_in_x254_fifoinpacked_0_active_0_out, // @[:@4751.4]
  input         io_sigsIn_backpressure, // @[:@4751.4]
  input         io_sigsIn_datapathEn, // @[:@4751.4]
  input         io_sigsIn_break, // @[:@4751.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_1, // @[:@4751.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@4751.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@4751.4]
  input         io_sigsIn_cchainOutputs_0_oobs_1, // @[:@4751.4]
  input         io_rr // @[:@4751.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4785.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@4785.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@4797.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@4797.4]
  wire  x516_sub_1_clock; // @[Math.scala 191:24:@4824.4]
  wire  x516_sub_1_reset; // @[Math.scala 191:24:@4824.4]
  wire [31:0] x516_sub_1_io_a; // @[Math.scala 191:24:@4824.4]
  wire [31:0] x516_sub_1_io_b; // @[Math.scala 191:24:@4824.4]
  wire  x516_sub_1_io_flow; // @[Math.scala 191:24:@4824.4]
  wire [31:0] x516_sub_1_io_result; // @[Math.scala 191:24:@4824.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@4834.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@4834.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@4834.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@4834.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@4834.4]
  wire  x264_sum_1_clock; // @[Math.scala 150:24:@4843.4]
  wire  x264_sum_1_reset; // @[Math.scala 150:24:@4843.4]
  wire [31:0] x264_sum_1_io_a; // @[Math.scala 150:24:@4843.4]
  wire [31:0] x264_sum_1_io_b; // @[Math.scala 150:24:@4843.4]
  wire  x264_sum_1_io_flow; // @[Math.scala 150:24:@4843.4]
  wire [31:0] x264_sum_1_io_result; // @[Math.scala 150:24:@4843.4]
  wire  x265_sum_1_clock; // @[Math.scala 150:24:@4855.4]
  wire  x265_sum_1_reset; // @[Math.scala 150:24:@4855.4]
  wire [31:0] x265_sum_1_io_a; // @[Math.scala 150:24:@4855.4]
  wire [31:0] x265_sum_1_io_b; // @[Math.scala 150:24:@4855.4]
  wire  x265_sum_1_io_flow; // @[Math.scala 150:24:@4855.4]
  wire [31:0] x265_sum_1_io_result; // @[Math.scala 150:24:@4855.4]
  wire [31:0] x267_1_io_b; // @[Math.scala 720:24:@4876.4]
  wire [31:0] x267_1_io_result; // @[Math.scala 720:24:@4876.4]
  wire  x268_sum_1_clock; // @[Math.scala 150:24:@4887.4]
  wire  x268_sum_1_reset; // @[Math.scala 150:24:@4887.4]
  wire [31:0] x268_sum_1_io_a; // @[Math.scala 150:24:@4887.4]
  wire [31:0] x268_sum_1_io_b; // @[Math.scala 150:24:@4887.4]
  wire  x268_sum_1_io_flow; // @[Math.scala 150:24:@4887.4]
  wire [31:0] x268_sum_1_io_result; // @[Math.scala 150:24:@4887.4]
  wire [31:0] x270_1_io_b; // @[Math.scala 720:24:@4908.4]
  wire [31:0] x270_1_io_result; // @[Math.scala 720:24:@4908.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@4923.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@4923.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@4923.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@4923.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@4923.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@4932.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@4932.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@4932.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@4932.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@4932.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@4943.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@4943.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@4943.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@4943.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@4943.4]
  wire  _T_327; // @[sm_x274_inr_Foreach.scala 62:18:@4810.4]
  wire  _T_328; // @[sm_x274_inr_Foreach.scala 62:55:@4811.4]
  wire [31:0] b259_number; // @[Math.scala 723:22:@4790.4 Math.scala 724:14:@4791.4]
  wire [42:0] _GEN_0; // @[Math.scala 461:32:@4815.4]
  wire [42:0] _T_331; // @[Math.scala 461:32:@4815.4]
  wire [38:0] _GEN_1; // @[Math.scala 461:32:@4820.4]
  wire [38:0] _T_334; // @[Math.scala 461:32:@4820.4]
  wire [31:0] x265_sum_number; // @[Math.scala 154:22:@4861.4 Math.scala 155:14:@4862.4]
  wire [31:0] _T_358; // @[Math.scala 406:49:@4868.4]
  wire [31:0] _T_360; // @[Math.scala 406:56:@4870.4]
  wire [31:0] _T_361; // @[Math.scala 406:56:@4871.4]
  wire [31:0] x268_sum_number; // @[Math.scala 154:22:@4893.4 Math.scala 155:14:@4894.4]
  wire [31:0] _T_380; // @[Math.scala 406:49:@4900.4]
  wire [31:0] _T_382; // @[Math.scala 406:56:@4902.4]
  wire [31:0] _T_383; // @[Math.scala 406:56:@4903.4]
  wire  _T_403; // @[sm_x274_inr_Foreach.scala 95:131:@4940.4]
  wire  _T_407; // @[package.scala 96:25:@4948.4 package.scala 96:25:@4949.4]
  wire  _T_409; // @[implicits.scala 55:10:@4950.4]
  wire  _T_410; // @[sm_x274_inr_Foreach.scala 95:148:@4951.4]
  wire  _T_412; // @[sm_x274_inr_Foreach.scala 95:236:@4953.4]
  wire  _T_413; // @[sm_x274_inr_Foreach.scala 95:255:@4954.4]
  wire  x542_b261_D3; // @[package.scala 96:25:@4937.4 package.scala 96:25:@4938.4]
  wire  _T_416; // @[sm_x274_inr_Foreach.scala 95:291:@4956.4]
  wire  x541_b262_D3; // @[package.scala 96:25:@4928.4 package.scala 96:25:@4929.4]
  _ _ ( // @[Math.scala 720:24:@4785.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@4797.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x516_sub x516_sub_1 ( // @[Math.scala 191:24:@4824.4]
    .clock(x516_sub_1_clock),
    .reset(x516_sub_1_reset),
    .io_a(x516_sub_1_io_a),
    .io_b(x516_sub_1_io_b),
    .io_flow(x516_sub_1_io_flow),
    .io_result(x516_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@4834.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x264_sum x264_sum_1 ( // @[Math.scala 150:24:@4843.4]
    .clock(x264_sum_1_clock),
    .reset(x264_sum_1_reset),
    .io_a(x264_sum_1_io_a),
    .io_b(x264_sum_1_io_b),
    .io_flow(x264_sum_1_io_flow),
    .io_result(x264_sum_1_io_result)
  );
  x264_sum x265_sum_1 ( // @[Math.scala 150:24:@4855.4]
    .clock(x265_sum_1_clock),
    .reset(x265_sum_1_reset),
    .io_a(x265_sum_1_io_a),
    .io_b(x265_sum_1_io_b),
    .io_flow(x265_sum_1_io_flow),
    .io_result(x265_sum_1_io_result)
  );
  _ x267_1 ( // @[Math.scala 720:24:@4876.4]
    .io_b(x267_1_io_b),
    .io_result(x267_1_io_result)
  );
  x264_sum x268_sum_1 ( // @[Math.scala 150:24:@4887.4]
    .clock(x268_sum_1_clock),
    .reset(x268_sum_1_reset),
    .io_a(x268_sum_1_io_a),
    .io_b(x268_sum_1_io_b),
    .io_flow(x268_sum_1_io_flow),
    .io_result(x268_sum_1_io_result)
  );
  _ x270_1 ( // @[Math.scala 720:24:@4908.4]
    .io_b(x270_1_io_b),
    .io_result(x270_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@4923.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_2 ( // @[package.scala 93:22:@4932.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_3 ( // @[package.scala 93:22:@4943.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_327 = ~ io_in_x254_fifoinpacked_0_full; // @[sm_x274_inr_Foreach.scala 62:18:@4810.4]
  assign _T_328 = ~ io_in_x254_fifoinpacked_0_active_0_out; // @[sm_x274_inr_Foreach.scala 62:55:@4811.4]
  assign b259_number = __io_result; // @[Math.scala 723:22:@4790.4 Math.scala 724:14:@4791.4]
  assign _GEN_0 = {{11'd0}, b259_number}; // @[Math.scala 461:32:@4815.4]
  assign _T_331 = _GEN_0 << 11; // @[Math.scala 461:32:@4815.4]
  assign _GEN_1 = {{7'd0}, b259_number}; // @[Math.scala 461:32:@4820.4]
  assign _T_334 = _GEN_1 << 7; // @[Math.scala 461:32:@4820.4]
  assign x265_sum_number = x265_sum_1_io_result; // @[Math.scala 154:22:@4861.4 Math.scala 155:14:@4862.4]
  assign _T_358 = $signed(x265_sum_number); // @[Math.scala 406:49:@4868.4]
  assign _T_360 = $signed(_T_358) & $signed(32'shff); // @[Math.scala 406:56:@4870.4]
  assign _T_361 = $signed(_T_360); // @[Math.scala 406:56:@4871.4]
  assign x268_sum_number = x268_sum_1_io_result; // @[Math.scala 154:22:@4893.4 Math.scala 155:14:@4894.4]
  assign _T_380 = $signed(x268_sum_number); // @[Math.scala 406:49:@4900.4]
  assign _T_382 = $signed(_T_380) & $signed(32'shff); // @[Math.scala 406:56:@4902.4]
  assign _T_383 = $signed(_T_382); // @[Math.scala 406:56:@4903.4]
  assign _T_403 = ~ io_sigsIn_break; // @[sm_x274_inr_Foreach.scala 95:131:@4940.4]
  assign _T_407 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@4948.4 package.scala 96:25:@4949.4]
  assign _T_409 = io_rr ? _T_407 : 1'h0; // @[implicits.scala 55:10:@4950.4]
  assign _T_410 = _T_403 & _T_409; // @[sm_x274_inr_Foreach.scala 95:148:@4951.4]
  assign _T_412 = _T_410 & _T_403; // @[sm_x274_inr_Foreach.scala 95:236:@4953.4]
  assign _T_413 = _T_412 & io_sigsIn_backpressure; // @[sm_x274_inr_Foreach.scala 95:255:@4954.4]
  assign x542_b261_D3 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@4937.4 package.scala 96:25:@4938.4]
  assign _T_416 = _T_413 & x542_b261_D3; // @[sm_x274_inr_Foreach.scala 95:291:@4956.4]
  assign x541_b262_D3 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@4928.4 package.scala 96:25:@4929.4]
  assign io_in_x254_fifoinpacked_0_wPort_0_en_0 = _T_416 & x541_b262_D3; // @[MemInterfaceType.scala 93:57:@4960.4]
  assign io_in_x254_fifoinpacked_0_active_0_in = x542_b261_D3 & x541_b262_D3; // @[MemInterfaceType.scala 147:18:@4963.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@4788.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@4800.4]
  assign x516_sub_1_clock = clock; // @[:@4825.4]
  assign x516_sub_1_reset = reset; // @[:@4826.4]
  assign x516_sub_1_io_a = _T_331[31:0]; // @[Math.scala 192:17:@4827.4]
  assign x516_sub_1_io_b = _T_334[31:0]; // @[Math.scala 193:17:@4828.4]
  assign x516_sub_1_io_flow = _T_327 | _T_328; // @[Math.scala 194:20:@4829.4]
  assign RetimeWrapper_clock = clock; // @[:@4835.4]
  assign RetimeWrapper_reset = reset; // @[:@4836.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4838.4]
  assign RetimeWrapper_io_in = __1_io_result; // @[package.scala 94:16:@4837.4]
  assign x264_sum_1_clock = clock; // @[:@4844.4]
  assign x264_sum_1_reset = reset; // @[:@4845.4]
  assign x264_sum_1_io_a = x516_sub_1_io_result; // @[Math.scala 151:17:@4846.4]
  assign x264_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@4847.4]
  assign x264_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4848.4]
  assign x265_sum_1_clock = clock; // @[:@4856.4]
  assign x265_sum_1_reset = reset; // @[:@4857.4]
  assign x265_sum_1_io_a = x264_sum_1_io_result; // @[Math.scala 151:17:@4858.4]
  assign x265_sum_1_io_b = 32'h1; // @[Math.scala 152:17:@4859.4]
  assign x265_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4860.4]
  assign x267_1_io_b = $unsigned(_T_361); // @[Math.scala 721:17:@4879.4]
  assign x268_sum_1_clock = clock; // @[:@4888.4]
  assign x268_sum_1_reset = reset; // @[:@4889.4]
  assign x268_sum_1_io_a = x264_sum_1_io_result; // @[Math.scala 151:17:@4890.4]
  assign x268_sum_1_io_b = 32'h2; // @[Math.scala 152:17:@4891.4]
  assign x268_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@4892.4]
  assign x270_1_io_b = $unsigned(_T_383); // @[Math.scala 721:17:@4911.4]
  assign RetimeWrapper_1_clock = clock; // @[:@4924.4]
  assign RetimeWrapper_1_reset = reset; // @[:@4925.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4927.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@4926.4]
  assign RetimeWrapper_2_clock = clock; // @[:@4933.4]
  assign RetimeWrapper_2_reset = reset; // @[:@4934.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4936.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@4935.4]
  assign RetimeWrapper_3_clock = clock; // @[:@4944.4]
  assign RetimeWrapper_3_reset = reset; // @[:@4945.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@4947.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@4946.4]
endmodule
module RetimeWrapper_42( // @[:@6081.2]
  input   clock, // @[:@6082.4]
  input   reset, // @[:@6083.4]
  input   io_flow, // @[:@6084.4]
  input   io_in, // @[:@6084.4]
  output  io_out // @[:@6084.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6086.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6086.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6086.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6086.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6086.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6086.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(97)) sr ( // @[RetimeShiftRegister.scala 15:20:@6086.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6099.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6098.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6097.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6096.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6095.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6093.4]
endmodule
module RetimeWrapper_46( // @[:@6209.2]
  input   clock, // @[:@6210.4]
  input   reset, // @[:@6211.4]
  input   io_flow, // @[:@6212.4]
  input   io_in, // @[:@6212.4]
  output  io_out // @[:@6212.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6214.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6214.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6214.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6214.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6214.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6214.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(96)) sr ( // @[RetimeShiftRegister.scala 15:20:@6214.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6227.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6226.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6225.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6224.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6223.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6221.4]
endmodule
module x465_inr_Foreach_SAMPLER_BOX_sm( // @[:@6229.2]
  input   clock, // @[:@6230.4]
  input   reset, // @[:@6231.4]
  input   io_enable, // @[:@6232.4]
  output  io_done, // @[:@6232.4]
  output  io_doneLatch, // @[:@6232.4]
  input   io_ctrDone, // @[:@6232.4]
  output  io_datapathEn, // @[:@6232.4]
  output  io_ctrInc, // @[:@6232.4]
  output  io_ctrRst, // @[:@6232.4]
  input   io_parentAck, // @[:@6232.4]
  input   io_backpressure, // @[:@6232.4]
  input   io_break // @[:@6232.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@6234.4]
  wire  active_reset; // @[Controllers.scala 261:22:@6234.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@6234.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@6234.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@6234.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@6234.4]
  wire  done_clock; // @[Controllers.scala 262:20:@6237.4]
  wire  done_reset; // @[Controllers.scala 262:20:@6237.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@6237.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@6237.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@6237.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@6237.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6271.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6271.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6271.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@6271.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@6271.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6293.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6293.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6293.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6293.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6293.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6305.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6305.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6305.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6305.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6305.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6313.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6313.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6313.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6313.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6313.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@6329.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@6329.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@6329.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@6329.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@6329.4]
  wire  _T_80; // @[Controllers.scala 264:48:@6242.4]
  wire  _T_81; // @[Controllers.scala 264:46:@6243.4]
  wire  _T_82; // @[Controllers.scala 264:62:@6244.4]
  wire  _T_83; // @[Controllers.scala 264:60:@6245.4]
  wire  _T_100; // @[package.scala 100:49:@6262.4]
  reg  _T_103; // @[package.scala 48:56:@6263.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@6276.4 package.scala 96:25:@6277.4]
  wire  _T_110; // @[package.scala 100:49:@6278.4]
  reg  _T_113; // @[package.scala 48:56:@6279.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@6281.4]
  wire  _T_118; // @[Controllers.scala 283:41:@6286.4]
  wire  _T_119; // @[Controllers.scala 283:59:@6287.4]
  wire  _T_121; // @[Controllers.scala 284:37:@6290.4]
  wire  _T_124; // @[package.scala 96:25:@6298.4 package.scala 96:25:@6299.4]
  wire  _T_126; // @[package.scala 100:49:@6300.4]
  reg  _T_129; // @[package.scala 48:56:@6301.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@6323.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@6325.4]
  reg  _T_153; // @[package.scala 48:56:@6326.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@6334.4 package.scala 96:25:@6335.4]
  wire  _T_158; // @[Controllers.scala 292:61:@6336.4]
  wire  _T_159; // @[Controllers.scala 292:24:@6337.4]
  SRFF active ( // @[Controllers.scala 261:22:@6234.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@6237.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_42 RetimeWrapper ( // @[package.scala 93:22:@6271.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_42 RetimeWrapper_1 ( // @[package.scala 93:22:@6293.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@6305.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@6313.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_46 RetimeWrapper_4 ( // @[package.scala 93:22:@6329.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@6242.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@6243.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@6244.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@6245.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@6262.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@6276.4 package.scala 96:25:@6277.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@6278.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@6281.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@6286.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@6287.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@6290.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6298.4 package.scala 96:25:@6299.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@6300.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@6325.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@6334.4 package.scala 96:25:@6335.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@6336.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@6337.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@6304.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@6339.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@6289.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@6292.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@6284.4]
  assign active_clock = clock; // @[:@6235.4]
  assign active_reset = reset; // @[:@6236.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@6247.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@6251.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@6252.4]
  assign done_clock = clock; // @[:@6238.4]
  assign done_reset = reset; // @[:@6239.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@6267.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@6260.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@6261.4]
  assign RetimeWrapper_clock = clock; // @[:@6272.4]
  assign RetimeWrapper_reset = reset; // @[:@6273.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@6275.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@6274.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6294.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6295.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@6297.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@6296.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6306.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6307.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@6309.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@6308.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6314.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6315.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@6317.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@6316.4]
  assign RetimeWrapper_4_clock = clock; // @[:@6330.4]
  assign RetimeWrapper_4_reset = reset; // @[:@6331.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@6333.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@6332.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module RetimeWrapper_50( // @[:@6530.2]
  input         clock, // @[:@6531.4]
  input         reset, // @[:@6532.4]
  input         io_flow, // @[:@6533.4]
  input  [63:0] io_in, // @[:@6533.4]
  output [63:0] io_out // @[:@6533.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@6535.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@6535.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@6535.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6535.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6535.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6535.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@6535.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6548.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6547.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@6546.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6545.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6544.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6542.4]
endmodule
module SRAM_1( // @[:@6566.2]
  input         clock, // @[:@6567.4]
  input         reset, // @[:@6568.4]
  input  [8:0]  io_raddr, // @[:@6569.4]
  input         io_wen, // @[:@6569.4]
  input  [8:0]  io_waddr, // @[:@6569.4]
  input  [31:0] io_wdata, // @[:@6569.4]
  output [31:0] io_rdata, // @[:@6569.4]
  input         io_backpressure // @[:@6569.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@6571.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@6571.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@6571.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@6571.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@6571.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@6571.4]
  wire [8:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@6571.4]
  wire [8:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@6571.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@6571.4]
  wire  _T_19; // @[SRAM.scala 182:49:@6589.4]
  wire  _T_20; // @[SRAM.scala 182:37:@6590.4]
  reg  _T_23; // @[SRAM.scala 182:29:@6591.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@6593.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(480), .AWIDTH(9)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@6571.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@6589.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@6590.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@6598.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@6585.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@6586.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@6583.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@6588.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@6587.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@6584.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@6582.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@6581.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module RetimeWrapper_51( // @[:@6612.2]
  input        clock, // @[:@6613.4]
  input        reset, // @[:@6614.4]
  input        io_flow, // @[:@6615.4]
  input  [8:0] io_in, // @[:@6615.4]
  output [8:0] io_out // @[:@6615.4]
);
  wire [8:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@6617.4]
  wire [8:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@6617.4]
  wire [8:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@6617.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6617.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6617.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6617.4]
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@6617.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6630.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6629.4]
  assign sr_init = 9'h0; // @[RetimeShiftRegister.scala 19:16:@6628.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6627.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6626.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6624.4]
endmodule
module Mem1D_5( // @[:@6632.2]
  input         clock, // @[:@6633.4]
  input         reset, // @[:@6634.4]
  input  [8:0]  io_r_ofs_0, // @[:@6635.4]
  input         io_r_backpressure, // @[:@6635.4]
  input  [8:0]  io_w_ofs_0, // @[:@6635.4]
  input  [31:0] io_w_data_0, // @[:@6635.4]
  input         io_w_en_0, // @[:@6635.4]
  output [31:0] io_output // @[:@6635.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@6639.4]
  wire  SRAM_reset; // @[MemPrimitives.scala 715:21:@6639.4]
  wire [8:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@6639.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 715:21:@6639.4]
  wire [8:0] SRAM_io_waddr; // @[MemPrimitives.scala 715:21:@6639.4]
  wire [31:0] SRAM_io_wdata; // @[MemPrimitives.scala 715:21:@6639.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@6639.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@6639.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6642.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6642.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6642.4]
  wire [8:0] RetimeWrapper_io_in; // @[package.scala 93:22:@6642.4]
  wire [8:0] RetimeWrapper_io_out; // @[package.scala 93:22:@6642.4]
  wire  wInBound; // @[MemPrimitives.scala 702:32:@6637.4]
  SRAM_1 SRAM ( // @[MemPrimitives.scala 715:21:@6639.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_51 RetimeWrapper ( // @[package.scala 93:22:@6642.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 9'h1e0; // @[MemPrimitives.scala 702:32:@6637.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@6655.4]
  assign SRAM_clock = clock; // @[:@6640.4]
  assign SRAM_reset = reset; // @[:@6641.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@6649.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 719:22:@6652.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 718:22:@6650.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 720:22:@6653.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@6654.4]
  assign RetimeWrapper_clock = clock; // @[:@6643.4]
  assign RetimeWrapper_reset = reset; // @[:@6644.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@6646.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@6645.4]
endmodule
module StickySelects_1( // @[:@8262.2]
  input   clock, // @[:@8263.4]
  input   reset, // @[:@8264.4]
  input   io_ins_0, // @[:@8265.4]
  input   io_ins_1, // @[:@8265.4]
  input   io_ins_2, // @[:@8265.4]
  input   io_ins_3, // @[:@8265.4]
  input   io_ins_4, // @[:@8265.4]
  input   io_ins_5, // @[:@8265.4]
  output  io_outs_0, // @[:@8265.4]
  output  io_outs_1, // @[:@8265.4]
  output  io_outs_2, // @[:@8265.4]
  output  io_outs_3, // @[:@8265.4]
  output  io_outs_4, // @[:@8265.4]
  output  io_outs_5 // @[:@8265.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@8267.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@8268.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@8269.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@8270.4]
  reg [31:0] _RAND_3;
  reg  _T_31; // @[StickySelects.scala 37:46:@8271.4]
  reg [31:0] _RAND_4;
  reg  _T_34; // @[StickySelects.scala 37:46:@8272.4]
  reg [31:0] _RAND_5;
  wire  _T_35; // @[StickySelects.scala 47:46:@8273.4]
  wire  _T_36; // @[StickySelects.scala 47:46:@8274.4]
  wire  _T_37; // @[StickySelects.scala 47:46:@8275.4]
  wire  _T_38; // @[StickySelects.scala 47:46:@8276.4]
  wire  _T_39; // @[StickySelects.scala 49:53:@8277.4]
  wire  _T_40; // @[StickySelects.scala 49:21:@8278.4]
  wire  _T_41; // @[StickySelects.scala 47:46:@8280.4]
  wire  _T_42; // @[StickySelects.scala 47:46:@8281.4]
  wire  _T_43; // @[StickySelects.scala 47:46:@8282.4]
  wire  _T_44; // @[StickySelects.scala 47:46:@8283.4]
  wire  _T_45; // @[StickySelects.scala 49:53:@8284.4]
  wire  _T_46; // @[StickySelects.scala 49:21:@8285.4]
  wire  _T_47; // @[StickySelects.scala 47:46:@8287.4]
  wire  _T_48; // @[StickySelects.scala 47:46:@8288.4]
  wire  _T_49; // @[StickySelects.scala 47:46:@8289.4]
  wire  _T_50; // @[StickySelects.scala 47:46:@8290.4]
  wire  _T_51; // @[StickySelects.scala 49:53:@8291.4]
  wire  _T_52; // @[StickySelects.scala 49:21:@8292.4]
  wire  _T_54; // @[StickySelects.scala 47:46:@8295.4]
  wire  _T_55; // @[StickySelects.scala 47:46:@8296.4]
  wire  _T_56; // @[StickySelects.scala 47:46:@8297.4]
  wire  _T_57; // @[StickySelects.scala 49:53:@8298.4]
  wire  _T_58; // @[StickySelects.scala 49:21:@8299.4]
  wire  _T_61; // @[StickySelects.scala 47:46:@8303.4]
  wire  _T_62; // @[StickySelects.scala 47:46:@8304.4]
  wire  _T_63; // @[StickySelects.scala 49:53:@8305.4]
  wire  _T_64; // @[StickySelects.scala 49:21:@8306.4]
  wire  _T_68; // @[StickySelects.scala 47:46:@8311.4]
  wire  _T_69; // @[StickySelects.scala 49:53:@8312.4]
  wire  _T_70; // @[StickySelects.scala 49:21:@8313.4]
  assign _T_35 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@8273.4]
  assign _T_36 = _T_35 | io_ins_3; // @[StickySelects.scala 47:46:@8274.4]
  assign _T_37 = _T_36 | io_ins_4; // @[StickySelects.scala 47:46:@8275.4]
  assign _T_38 = _T_37 | io_ins_5; // @[StickySelects.scala 47:46:@8276.4]
  assign _T_39 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@8277.4]
  assign _T_40 = _T_38 ? io_ins_0 : _T_39; // @[StickySelects.scala 49:21:@8278.4]
  assign _T_41 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@8280.4]
  assign _T_42 = _T_41 | io_ins_3; // @[StickySelects.scala 47:46:@8281.4]
  assign _T_43 = _T_42 | io_ins_4; // @[StickySelects.scala 47:46:@8282.4]
  assign _T_44 = _T_43 | io_ins_5; // @[StickySelects.scala 47:46:@8283.4]
  assign _T_45 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@8284.4]
  assign _T_46 = _T_44 ? io_ins_1 : _T_45; // @[StickySelects.scala 49:21:@8285.4]
  assign _T_47 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@8287.4]
  assign _T_48 = _T_47 | io_ins_3; // @[StickySelects.scala 47:46:@8288.4]
  assign _T_49 = _T_48 | io_ins_4; // @[StickySelects.scala 47:46:@8289.4]
  assign _T_50 = _T_49 | io_ins_5; // @[StickySelects.scala 47:46:@8290.4]
  assign _T_51 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@8291.4]
  assign _T_52 = _T_50 ? io_ins_2 : _T_51; // @[StickySelects.scala 49:21:@8292.4]
  assign _T_54 = _T_47 | io_ins_2; // @[StickySelects.scala 47:46:@8295.4]
  assign _T_55 = _T_54 | io_ins_4; // @[StickySelects.scala 47:46:@8296.4]
  assign _T_56 = _T_55 | io_ins_5; // @[StickySelects.scala 47:46:@8297.4]
  assign _T_57 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@8298.4]
  assign _T_58 = _T_56 ? io_ins_3 : _T_57; // @[StickySelects.scala 49:21:@8299.4]
  assign _T_61 = _T_54 | io_ins_3; // @[StickySelects.scala 47:46:@8303.4]
  assign _T_62 = _T_61 | io_ins_5; // @[StickySelects.scala 47:46:@8304.4]
  assign _T_63 = io_ins_4 | _T_31; // @[StickySelects.scala 49:53:@8305.4]
  assign _T_64 = _T_62 ? io_ins_4 : _T_63; // @[StickySelects.scala 49:21:@8306.4]
  assign _T_68 = _T_61 | io_ins_4; // @[StickySelects.scala 47:46:@8311.4]
  assign _T_69 = io_ins_5 | _T_34; // @[StickySelects.scala 49:53:@8312.4]
  assign _T_70 = _T_68 ? io_ins_5 : _T_69; // @[StickySelects.scala 49:21:@8313.4]
  assign io_outs_0 = _T_38 ? io_ins_0 : _T_39; // @[StickySelects.scala 53:57:@8315.4]
  assign io_outs_1 = _T_44 ? io_ins_1 : _T_45; // @[StickySelects.scala 53:57:@8316.4]
  assign io_outs_2 = _T_50 ? io_ins_2 : _T_51; // @[StickySelects.scala 53:57:@8317.4]
  assign io_outs_3 = _T_56 ? io_ins_3 : _T_57; // @[StickySelects.scala 53:57:@8318.4]
  assign io_outs_4 = _T_62 ? io_ins_4 : _T_63; // @[StickySelects.scala 53:57:@8319.4]
  assign io_outs_5 = _T_68 ? io_ins_5 : _T_69; // @[StickySelects.scala 53:57:@8320.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_31 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_38) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_39;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_44) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_45;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_50) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_51;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_56) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_57;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_62) begin
        _T_31 <= io_ins_4;
      end else begin
        _T_31 <= _T_63;
      end
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (_T_68) begin
        _T_34 <= io_ins_5;
      end else begin
        _T_34 <= _T_69;
      end
    end
  end
endmodule
module x285_lb_0( // @[:@12294.2]
  input         clock, // @[:@12295.4]
  input         reset, // @[:@12296.4]
  input  [2:0]  io_rPort_11_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_11_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_11_ofs_0, // @[:@12297.4]
  input         io_rPort_11_en_0, // @[:@12297.4]
  input         io_rPort_11_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_11_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_10_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_10_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_10_ofs_0, // @[:@12297.4]
  input         io_rPort_10_en_0, // @[:@12297.4]
  input         io_rPort_10_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_10_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_9_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_9_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_9_ofs_0, // @[:@12297.4]
  input         io_rPort_9_en_0, // @[:@12297.4]
  input         io_rPort_9_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_9_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_8_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_8_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_8_ofs_0, // @[:@12297.4]
  input         io_rPort_8_en_0, // @[:@12297.4]
  input         io_rPort_8_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_8_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_7_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_7_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_7_ofs_0, // @[:@12297.4]
  input         io_rPort_7_en_0, // @[:@12297.4]
  input         io_rPort_7_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_7_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_6_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_6_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_6_ofs_0, // @[:@12297.4]
  input         io_rPort_6_en_0, // @[:@12297.4]
  input         io_rPort_6_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_6_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_5_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_5_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_5_ofs_0, // @[:@12297.4]
  input         io_rPort_5_en_0, // @[:@12297.4]
  input         io_rPort_5_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_5_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_4_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_4_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_4_ofs_0, // @[:@12297.4]
  input         io_rPort_4_en_0, // @[:@12297.4]
  input         io_rPort_4_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_4_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_3_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_3_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_3_ofs_0, // @[:@12297.4]
  input         io_rPort_3_en_0, // @[:@12297.4]
  input         io_rPort_3_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_3_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_2_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_2_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_2_ofs_0, // @[:@12297.4]
  input         io_rPort_2_en_0, // @[:@12297.4]
  input         io_rPort_2_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_2_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_1_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_1_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_1_ofs_0, // @[:@12297.4]
  input         io_rPort_1_en_0, // @[:@12297.4]
  input         io_rPort_1_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_1_output_0, // @[:@12297.4]
  input  [2:0]  io_rPort_0_banks_1, // @[:@12297.4]
  input  [2:0]  io_rPort_0_banks_0, // @[:@12297.4]
  input  [8:0]  io_rPort_0_ofs_0, // @[:@12297.4]
  input         io_rPort_0_en_0, // @[:@12297.4]
  input         io_rPort_0_backpressure, // @[:@12297.4]
  output [31:0] io_rPort_0_output_0, // @[:@12297.4]
  input  [2:0]  io_wPort_1_banks_1, // @[:@12297.4]
  input  [2:0]  io_wPort_1_banks_0, // @[:@12297.4]
  input  [8:0]  io_wPort_1_ofs_0, // @[:@12297.4]
  input  [31:0] io_wPort_1_data_0, // @[:@12297.4]
  input         io_wPort_1_en_0, // @[:@12297.4]
  input  [2:0]  io_wPort_0_banks_1, // @[:@12297.4]
  input  [2:0]  io_wPort_0_banks_0, // @[:@12297.4]
  input  [8:0]  io_wPort_0_ofs_0, // @[:@12297.4]
  input  [31:0] io_wPort_0_data_0, // @[:@12297.4]
  input         io_wPort_0_en_0 // @[:@12297.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@12388.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@12388.4]
  wire [8:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12388.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12388.4]
  wire [8:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12388.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@12388.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@12388.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@12388.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@12404.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@12404.4]
  wire [8:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12404.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12404.4]
  wire [8:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12404.4]
  wire [31:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@12404.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@12404.4]
  wire [31:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@12404.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@12420.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@12420.4]
  wire [8:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12420.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12420.4]
  wire [8:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12420.4]
  wire [31:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@12420.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@12420.4]
  wire [31:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@12420.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@12436.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@12436.4]
  wire [8:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12436.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12436.4]
  wire [8:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12436.4]
  wire [31:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@12436.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@12436.4]
  wire [31:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@12436.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@12452.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@12452.4]
  wire [8:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12452.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12452.4]
  wire [8:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12452.4]
  wire [31:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@12452.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@12452.4]
  wire [31:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@12452.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@12468.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@12468.4]
  wire [8:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12468.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12468.4]
  wire [8:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12468.4]
  wire [31:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@12468.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@12468.4]
  wire [31:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@12468.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@12484.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@12484.4]
  wire [8:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12484.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12484.4]
  wire [8:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12484.4]
  wire [31:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@12484.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@12484.4]
  wire [31:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@12484.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@12500.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@12500.4]
  wire [8:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12500.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12500.4]
  wire [8:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12500.4]
  wire [31:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@12500.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@12500.4]
  wire [31:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@12500.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@12516.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@12516.4]
  wire [8:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12516.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12516.4]
  wire [8:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12516.4]
  wire [31:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@12516.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@12516.4]
  wire [31:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@12516.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@12532.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@12532.4]
  wire [8:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12532.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12532.4]
  wire [8:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12532.4]
  wire [31:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@12532.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@12532.4]
  wire [31:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@12532.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@12548.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@12548.4]
  wire [8:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12548.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12548.4]
  wire [8:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12548.4]
  wire [31:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@12548.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@12548.4]
  wire [31:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@12548.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@12564.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@12564.4]
  wire [8:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12564.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12564.4]
  wire [8:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12564.4]
  wire [31:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@12564.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@12564.4]
  wire [31:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@12564.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@12580.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@12580.4]
  wire [8:0] Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12580.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12580.4]
  wire [8:0] Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12580.4]
  wire [31:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@12580.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@12580.4]
  wire [31:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@12580.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@12596.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@12596.4]
  wire [8:0] Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12596.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12596.4]
  wire [8:0] Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12596.4]
  wire [31:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@12596.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@12596.4]
  wire [31:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@12596.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@12612.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@12612.4]
  wire [8:0] Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12612.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12612.4]
  wire [8:0] Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12612.4]
  wire [31:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@12612.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@12612.4]
  wire [31:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@12612.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@12628.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@12628.4]
  wire [8:0] Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12628.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12628.4]
  wire [8:0] Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12628.4]
  wire [31:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@12628.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@12628.4]
  wire [31:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@12628.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 124:33:@12860.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 124:33:@12922.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 124:33:@12984.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 124:33:@13046.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 124:33:@13108.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 124:33:@13170.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 124:33:@13232.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 124:33:@13294.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 124:33:@13356.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 124:33:@13418.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 124:33:@13480.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 124:33:@13542.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_ins_4; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_ins_5; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_outs_4; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_12_io_outs_5; // @[MemPrimitives.scala 124:33:@13604.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_ins_4; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_ins_5; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_outs_4; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_13_io_outs_5; // @[MemPrimitives.scala 124:33:@13666.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 124:33:@13728.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 124:33:@13790.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@13853.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@13853.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@13853.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@13853.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@13853.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@13861.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@13861.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@13861.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@13861.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@13861.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@13869.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@13869.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@13869.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@13869.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@13869.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@13877.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@13877.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@13877.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@13877.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@13877.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@13885.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@13885.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@13885.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@13885.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@13885.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@13893.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@13893.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@13893.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@13893.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@13893.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@13901.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@13901.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@13901.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@13901.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@13901.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@13909.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@13909.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@13909.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@13909.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@13909.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@13949.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@13949.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@13949.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@13949.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@13949.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@13957.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@13957.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@13957.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@13957.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@13957.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@13965.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@13965.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@13965.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@13965.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@13965.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@13973.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@13973.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@13973.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@13973.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@13973.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@13981.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@13981.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@13981.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@13981.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@13981.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@13989.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@13989.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@13989.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@13989.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@13989.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@13997.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@13997.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@13997.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@13997.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@13997.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@14005.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@14005.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@14005.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@14005.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@14005.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@14045.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@14045.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@14045.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@14045.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@14045.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@14053.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@14053.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@14053.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@14053.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@14053.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@14061.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@14061.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@14061.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@14061.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@14061.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@14069.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@14069.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@14069.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@14069.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@14069.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@14077.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@14077.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@14077.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@14077.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@14077.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@14085.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@14085.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@14085.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@14085.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@14085.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@14093.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@14093.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@14093.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@14093.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@14093.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@14101.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@14101.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@14101.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@14101.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@14101.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@14141.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@14141.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@14141.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@14141.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@14141.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@14149.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@14149.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@14149.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@14149.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@14149.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@14157.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@14157.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@14157.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@14157.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@14157.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@14165.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@14165.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@14165.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@14165.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@14165.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@14173.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@14173.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@14173.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@14173.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@14173.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@14181.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@14181.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@14181.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@14181.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@14181.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@14189.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@14189.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@14189.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@14189.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@14189.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@14197.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@14197.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@14197.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@14197.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@14197.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@14237.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@14237.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@14237.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@14237.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@14237.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@14245.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@14245.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@14245.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@14245.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@14245.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@14253.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@14253.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@14253.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@14253.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@14253.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@14261.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@14261.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@14261.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@14261.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@14261.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@14269.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@14269.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@14269.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@14269.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@14269.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@14277.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@14277.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@14277.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@14277.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@14277.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@14285.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@14285.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@14285.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@14285.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@14285.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@14293.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@14293.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@14293.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@14293.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@14293.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@14333.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@14333.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@14333.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@14333.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@14333.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@14341.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@14341.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@14341.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@14341.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@14341.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@14349.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@14349.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@14349.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@14349.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@14349.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@14357.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@14357.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@14357.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@14357.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@14357.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@14365.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@14365.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@14365.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@14365.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@14365.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@14373.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@14373.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@14373.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@14373.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@14373.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@14381.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@14381.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@14381.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@14381.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@14381.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@14389.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@14389.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@14389.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@14389.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@14389.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@14429.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@14429.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@14429.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@14429.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@14429.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@14437.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@14437.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@14437.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@14437.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@14437.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@14445.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@14445.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@14445.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@14445.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@14445.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@14453.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@14453.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@14453.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@14453.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@14453.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@14461.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@14461.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@14461.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@14461.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@14461.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@14469.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@14469.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@14469.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@14469.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@14469.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@14477.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@14477.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@14477.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@14477.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@14477.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@14485.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@14485.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@14485.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@14485.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@14485.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@14525.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@14525.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@14525.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@14525.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@14525.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@14533.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@14533.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@14533.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@14533.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@14533.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@14541.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@14541.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@14541.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@14541.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@14541.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@14549.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@14549.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@14549.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@14549.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@14549.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@14557.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@14557.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@14557.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@14557.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@14557.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@14565.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@14565.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@14565.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@14565.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@14565.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@14573.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@14573.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@14573.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@14573.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@14573.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@14581.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@14581.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@14581.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@14581.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@14581.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@14621.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@14621.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@14621.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@14621.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@14621.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@14629.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@14629.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@14629.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@14629.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@14629.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@14637.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@14637.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@14637.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@14637.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@14637.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@14645.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@14645.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@14645.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@14645.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@14645.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@14653.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@14653.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@14653.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@14653.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@14653.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@14661.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@14661.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@14661.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@14661.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@14661.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@14669.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@14669.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@14669.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@14669.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@14669.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@14677.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@14677.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@14677.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@14677.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@14677.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@14717.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@14717.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@14717.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@14717.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@14717.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@14725.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@14725.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@14725.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@14725.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@14725.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@14733.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@14741.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@14741.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@14741.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@14741.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@14741.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@14749.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@14749.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@14749.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@14749.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@14749.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@14757.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@14757.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@14757.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@14757.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@14757.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@14765.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@14765.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@14765.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@14765.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@14765.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@14773.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@14773.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@14773.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@14773.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@14773.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@14813.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@14813.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@14813.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@14813.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@14813.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@14821.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@14821.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@14821.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@14821.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@14821.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@14829.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@14829.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@14829.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@14829.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@14829.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@14837.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@14837.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@14837.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@14837.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@14837.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@14845.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@14845.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@14845.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@14845.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@14845.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@14853.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@14853.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@14853.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@14853.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@14853.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@14861.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@14861.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@14861.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@14861.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@14861.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@14869.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@14869.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@14869.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@14869.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@14869.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@14909.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@14909.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@14909.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@14909.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@14909.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@14917.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@14917.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@14917.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@14917.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@14917.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@14925.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@14925.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@14925.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@14925.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@14925.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@14933.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@14933.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@14933.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@14933.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@14933.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@14941.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@14941.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@14941.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@14941.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@14941.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@14949.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@14949.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@14949.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@14949.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@14949.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@14957.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@14957.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@14957.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@14957.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@14957.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@14965.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@14965.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@14965.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@14965.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@14965.4]
  wire  _T_444; // @[MemPrimitives.scala 82:210:@12644.4]
  wire  _T_446; // @[MemPrimitives.scala 82:210:@12645.4]
  wire  _T_447; // @[MemPrimitives.scala 82:228:@12646.4]
  wire  _T_448; // @[MemPrimitives.scala 83:102:@12647.4]
  wire [41:0] _T_450; // @[Cat.scala 30:58:@12649.4]
  wire  _T_455; // @[MemPrimitives.scala 82:210:@12656.4]
  wire  _T_457; // @[MemPrimitives.scala 82:210:@12657.4]
  wire  _T_458; // @[MemPrimitives.scala 82:228:@12658.4]
  wire  _T_459; // @[MemPrimitives.scala 83:102:@12659.4]
  wire [41:0] _T_461; // @[Cat.scala 30:58:@12661.4]
  wire  _T_468; // @[MemPrimitives.scala 82:210:@12669.4]
  wire  _T_469; // @[MemPrimitives.scala 82:228:@12670.4]
  wire  _T_470; // @[MemPrimitives.scala 83:102:@12671.4]
  wire [41:0] _T_472; // @[Cat.scala 30:58:@12673.4]
  wire  _T_479; // @[MemPrimitives.scala 82:210:@12681.4]
  wire  _T_480; // @[MemPrimitives.scala 82:228:@12682.4]
  wire  _T_481; // @[MemPrimitives.scala 83:102:@12683.4]
  wire [41:0] _T_483; // @[Cat.scala 30:58:@12685.4]
  wire  _T_488; // @[MemPrimitives.scala 82:210:@12692.4]
  wire  _T_491; // @[MemPrimitives.scala 82:228:@12694.4]
  wire  _T_492; // @[MemPrimitives.scala 83:102:@12695.4]
  wire [41:0] _T_494; // @[Cat.scala 30:58:@12697.4]
  wire  _T_499; // @[MemPrimitives.scala 82:210:@12704.4]
  wire  _T_502; // @[MemPrimitives.scala 82:228:@12706.4]
  wire  _T_503; // @[MemPrimitives.scala 83:102:@12707.4]
  wire [41:0] _T_505; // @[Cat.scala 30:58:@12709.4]
  wire  _T_513; // @[MemPrimitives.scala 82:228:@12718.4]
  wire  _T_514; // @[MemPrimitives.scala 83:102:@12719.4]
  wire [41:0] _T_516; // @[Cat.scala 30:58:@12721.4]
  wire  _T_524; // @[MemPrimitives.scala 82:228:@12730.4]
  wire  _T_525; // @[MemPrimitives.scala 83:102:@12731.4]
  wire [41:0] _T_527; // @[Cat.scala 30:58:@12733.4]
  wire  _T_532; // @[MemPrimitives.scala 82:210:@12740.4]
  wire  _T_535; // @[MemPrimitives.scala 82:228:@12742.4]
  wire  _T_536; // @[MemPrimitives.scala 83:102:@12743.4]
  wire [41:0] _T_538; // @[Cat.scala 30:58:@12745.4]
  wire  _T_543; // @[MemPrimitives.scala 82:210:@12752.4]
  wire  _T_546; // @[MemPrimitives.scala 82:228:@12754.4]
  wire  _T_547; // @[MemPrimitives.scala 83:102:@12755.4]
  wire [41:0] _T_549; // @[Cat.scala 30:58:@12757.4]
  wire  _T_557; // @[MemPrimitives.scala 82:228:@12766.4]
  wire  _T_558; // @[MemPrimitives.scala 83:102:@12767.4]
  wire [41:0] _T_560; // @[Cat.scala 30:58:@12769.4]
  wire  _T_568; // @[MemPrimitives.scala 82:228:@12778.4]
  wire  _T_569; // @[MemPrimitives.scala 83:102:@12779.4]
  wire [41:0] _T_571; // @[Cat.scala 30:58:@12781.4]
  wire  _T_576; // @[MemPrimitives.scala 82:210:@12788.4]
  wire  _T_579; // @[MemPrimitives.scala 82:228:@12790.4]
  wire  _T_580; // @[MemPrimitives.scala 83:102:@12791.4]
  wire [41:0] _T_582; // @[Cat.scala 30:58:@12793.4]
  wire  _T_587; // @[MemPrimitives.scala 82:210:@12800.4]
  wire  _T_590; // @[MemPrimitives.scala 82:228:@12802.4]
  wire  _T_591; // @[MemPrimitives.scala 83:102:@12803.4]
  wire [41:0] _T_593; // @[Cat.scala 30:58:@12805.4]
  wire  _T_601; // @[MemPrimitives.scala 82:228:@12814.4]
  wire  _T_602; // @[MemPrimitives.scala 83:102:@12815.4]
  wire [41:0] _T_604; // @[Cat.scala 30:58:@12817.4]
  wire  _T_612; // @[MemPrimitives.scala 82:228:@12826.4]
  wire  _T_613; // @[MemPrimitives.scala 83:102:@12827.4]
  wire [41:0] _T_615; // @[Cat.scala 30:58:@12829.4]
  wire  _T_620; // @[MemPrimitives.scala 110:210:@12836.4]
  wire  _T_622; // @[MemPrimitives.scala 110:210:@12837.4]
  wire  _T_623; // @[MemPrimitives.scala 110:228:@12838.4]
  wire  _T_626; // @[MemPrimitives.scala 110:210:@12840.4]
  wire  _T_628; // @[MemPrimitives.scala 110:210:@12841.4]
  wire  _T_629; // @[MemPrimitives.scala 110:228:@12842.4]
  wire  _T_632; // @[MemPrimitives.scala 110:210:@12844.4]
  wire  _T_634; // @[MemPrimitives.scala 110:210:@12845.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@12846.4]
  wire  _T_638; // @[MemPrimitives.scala 110:210:@12848.4]
  wire  _T_640; // @[MemPrimitives.scala 110:210:@12849.4]
  wire  _T_641; // @[MemPrimitives.scala 110:228:@12850.4]
  wire  _T_644; // @[MemPrimitives.scala 110:210:@12852.4]
  wire  _T_646; // @[MemPrimitives.scala 110:210:@12853.4]
  wire  _T_647; // @[MemPrimitives.scala 110:228:@12854.4]
  wire  _T_650; // @[MemPrimitives.scala 110:210:@12856.4]
  wire  _T_652; // @[MemPrimitives.scala 110:210:@12857.4]
  wire  _T_653; // @[MemPrimitives.scala 110:228:@12858.4]
  wire  _T_655; // @[MemPrimitives.scala 126:35:@12869.4]
  wire  _T_656; // @[MemPrimitives.scala 126:35:@12870.4]
  wire  _T_657; // @[MemPrimitives.scala 126:35:@12871.4]
  wire  _T_658; // @[MemPrimitives.scala 126:35:@12872.4]
  wire  _T_659; // @[MemPrimitives.scala 126:35:@12873.4]
  wire  _T_660; // @[MemPrimitives.scala 126:35:@12874.4]
  wire [10:0] _T_662; // @[Cat.scala 30:58:@12876.4]
  wire [10:0] _T_664; // @[Cat.scala 30:58:@12878.4]
  wire [10:0] _T_666; // @[Cat.scala 30:58:@12880.4]
  wire [10:0] _T_668; // @[Cat.scala 30:58:@12882.4]
  wire [10:0] _T_670; // @[Cat.scala 30:58:@12884.4]
  wire [10:0] _T_672; // @[Cat.scala 30:58:@12886.4]
  wire [10:0] _T_673; // @[Mux.scala 31:69:@12887.4]
  wire [10:0] _T_674; // @[Mux.scala 31:69:@12888.4]
  wire [10:0] _T_675; // @[Mux.scala 31:69:@12889.4]
  wire [10:0] _T_676; // @[Mux.scala 31:69:@12890.4]
  wire [10:0] _T_677; // @[Mux.scala 31:69:@12891.4]
  wire  _T_682; // @[MemPrimitives.scala 110:210:@12898.4]
  wire  _T_684; // @[MemPrimitives.scala 110:210:@12899.4]
  wire  _T_685; // @[MemPrimitives.scala 110:228:@12900.4]
  wire  _T_688; // @[MemPrimitives.scala 110:210:@12902.4]
  wire  _T_690; // @[MemPrimitives.scala 110:210:@12903.4]
  wire  _T_691; // @[MemPrimitives.scala 110:228:@12904.4]
  wire  _T_694; // @[MemPrimitives.scala 110:210:@12906.4]
  wire  _T_696; // @[MemPrimitives.scala 110:210:@12907.4]
  wire  _T_697; // @[MemPrimitives.scala 110:228:@12908.4]
  wire  _T_700; // @[MemPrimitives.scala 110:210:@12910.4]
  wire  _T_702; // @[MemPrimitives.scala 110:210:@12911.4]
  wire  _T_703; // @[MemPrimitives.scala 110:228:@12912.4]
  wire  _T_706; // @[MemPrimitives.scala 110:210:@12914.4]
  wire  _T_708; // @[MemPrimitives.scala 110:210:@12915.4]
  wire  _T_709; // @[MemPrimitives.scala 110:228:@12916.4]
  wire  _T_712; // @[MemPrimitives.scala 110:210:@12918.4]
  wire  _T_714; // @[MemPrimitives.scala 110:210:@12919.4]
  wire  _T_715; // @[MemPrimitives.scala 110:228:@12920.4]
  wire  _T_717; // @[MemPrimitives.scala 126:35:@12931.4]
  wire  _T_718; // @[MemPrimitives.scala 126:35:@12932.4]
  wire  _T_719; // @[MemPrimitives.scala 126:35:@12933.4]
  wire  _T_720; // @[MemPrimitives.scala 126:35:@12934.4]
  wire  _T_721; // @[MemPrimitives.scala 126:35:@12935.4]
  wire  _T_722; // @[MemPrimitives.scala 126:35:@12936.4]
  wire [10:0] _T_724; // @[Cat.scala 30:58:@12938.4]
  wire [10:0] _T_726; // @[Cat.scala 30:58:@12940.4]
  wire [10:0] _T_728; // @[Cat.scala 30:58:@12942.4]
  wire [10:0] _T_730; // @[Cat.scala 30:58:@12944.4]
  wire [10:0] _T_732; // @[Cat.scala 30:58:@12946.4]
  wire [10:0] _T_734; // @[Cat.scala 30:58:@12948.4]
  wire [10:0] _T_735; // @[Mux.scala 31:69:@12949.4]
  wire [10:0] _T_736; // @[Mux.scala 31:69:@12950.4]
  wire [10:0] _T_737; // @[Mux.scala 31:69:@12951.4]
  wire [10:0] _T_738; // @[Mux.scala 31:69:@12952.4]
  wire [10:0] _T_739; // @[Mux.scala 31:69:@12953.4]
  wire  _T_746; // @[MemPrimitives.scala 110:210:@12961.4]
  wire  _T_747; // @[MemPrimitives.scala 110:228:@12962.4]
  wire  _T_752; // @[MemPrimitives.scala 110:210:@12965.4]
  wire  _T_753; // @[MemPrimitives.scala 110:228:@12966.4]
  wire  _T_758; // @[MemPrimitives.scala 110:210:@12969.4]
  wire  _T_759; // @[MemPrimitives.scala 110:228:@12970.4]
  wire  _T_764; // @[MemPrimitives.scala 110:210:@12973.4]
  wire  _T_765; // @[MemPrimitives.scala 110:228:@12974.4]
  wire  _T_770; // @[MemPrimitives.scala 110:210:@12977.4]
  wire  _T_771; // @[MemPrimitives.scala 110:228:@12978.4]
  wire  _T_776; // @[MemPrimitives.scala 110:210:@12981.4]
  wire  _T_777; // @[MemPrimitives.scala 110:228:@12982.4]
  wire  _T_779; // @[MemPrimitives.scala 126:35:@12993.4]
  wire  _T_780; // @[MemPrimitives.scala 126:35:@12994.4]
  wire  _T_781; // @[MemPrimitives.scala 126:35:@12995.4]
  wire  _T_782; // @[MemPrimitives.scala 126:35:@12996.4]
  wire  _T_783; // @[MemPrimitives.scala 126:35:@12997.4]
  wire  _T_784; // @[MemPrimitives.scala 126:35:@12998.4]
  wire [10:0] _T_786; // @[Cat.scala 30:58:@13000.4]
  wire [10:0] _T_788; // @[Cat.scala 30:58:@13002.4]
  wire [10:0] _T_790; // @[Cat.scala 30:58:@13004.4]
  wire [10:0] _T_792; // @[Cat.scala 30:58:@13006.4]
  wire [10:0] _T_794; // @[Cat.scala 30:58:@13008.4]
  wire [10:0] _T_796; // @[Cat.scala 30:58:@13010.4]
  wire [10:0] _T_797; // @[Mux.scala 31:69:@13011.4]
  wire [10:0] _T_798; // @[Mux.scala 31:69:@13012.4]
  wire [10:0] _T_799; // @[Mux.scala 31:69:@13013.4]
  wire [10:0] _T_800; // @[Mux.scala 31:69:@13014.4]
  wire [10:0] _T_801; // @[Mux.scala 31:69:@13015.4]
  wire  _T_808; // @[MemPrimitives.scala 110:210:@13023.4]
  wire  _T_809; // @[MemPrimitives.scala 110:228:@13024.4]
  wire  _T_814; // @[MemPrimitives.scala 110:210:@13027.4]
  wire  _T_815; // @[MemPrimitives.scala 110:228:@13028.4]
  wire  _T_820; // @[MemPrimitives.scala 110:210:@13031.4]
  wire  _T_821; // @[MemPrimitives.scala 110:228:@13032.4]
  wire  _T_826; // @[MemPrimitives.scala 110:210:@13035.4]
  wire  _T_827; // @[MemPrimitives.scala 110:228:@13036.4]
  wire  _T_832; // @[MemPrimitives.scala 110:210:@13039.4]
  wire  _T_833; // @[MemPrimitives.scala 110:228:@13040.4]
  wire  _T_838; // @[MemPrimitives.scala 110:210:@13043.4]
  wire  _T_839; // @[MemPrimitives.scala 110:228:@13044.4]
  wire  _T_841; // @[MemPrimitives.scala 126:35:@13055.4]
  wire  _T_842; // @[MemPrimitives.scala 126:35:@13056.4]
  wire  _T_843; // @[MemPrimitives.scala 126:35:@13057.4]
  wire  _T_844; // @[MemPrimitives.scala 126:35:@13058.4]
  wire  _T_845; // @[MemPrimitives.scala 126:35:@13059.4]
  wire  _T_846; // @[MemPrimitives.scala 126:35:@13060.4]
  wire [10:0] _T_848; // @[Cat.scala 30:58:@13062.4]
  wire [10:0] _T_850; // @[Cat.scala 30:58:@13064.4]
  wire [10:0] _T_852; // @[Cat.scala 30:58:@13066.4]
  wire [10:0] _T_854; // @[Cat.scala 30:58:@13068.4]
  wire [10:0] _T_856; // @[Cat.scala 30:58:@13070.4]
  wire [10:0] _T_858; // @[Cat.scala 30:58:@13072.4]
  wire [10:0] _T_859; // @[Mux.scala 31:69:@13073.4]
  wire [10:0] _T_860; // @[Mux.scala 31:69:@13074.4]
  wire [10:0] _T_861; // @[Mux.scala 31:69:@13075.4]
  wire [10:0] _T_862; // @[Mux.scala 31:69:@13076.4]
  wire [10:0] _T_863; // @[Mux.scala 31:69:@13077.4]
  wire  _T_868; // @[MemPrimitives.scala 110:210:@13084.4]
  wire  _T_871; // @[MemPrimitives.scala 110:228:@13086.4]
  wire  _T_874; // @[MemPrimitives.scala 110:210:@13088.4]
  wire  _T_877; // @[MemPrimitives.scala 110:228:@13090.4]
  wire  _T_880; // @[MemPrimitives.scala 110:210:@13092.4]
  wire  _T_883; // @[MemPrimitives.scala 110:228:@13094.4]
  wire  _T_886; // @[MemPrimitives.scala 110:210:@13096.4]
  wire  _T_889; // @[MemPrimitives.scala 110:228:@13098.4]
  wire  _T_892; // @[MemPrimitives.scala 110:210:@13100.4]
  wire  _T_895; // @[MemPrimitives.scala 110:228:@13102.4]
  wire  _T_898; // @[MemPrimitives.scala 110:210:@13104.4]
  wire  _T_901; // @[MemPrimitives.scala 110:228:@13106.4]
  wire  _T_903; // @[MemPrimitives.scala 126:35:@13117.4]
  wire  _T_904; // @[MemPrimitives.scala 126:35:@13118.4]
  wire  _T_905; // @[MemPrimitives.scala 126:35:@13119.4]
  wire  _T_906; // @[MemPrimitives.scala 126:35:@13120.4]
  wire  _T_907; // @[MemPrimitives.scala 126:35:@13121.4]
  wire  _T_908; // @[MemPrimitives.scala 126:35:@13122.4]
  wire [10:0] _T_910; // @[Cat.scala 30:58:@13124.4]
  wire [10:0] _T_912; // @[Cat.scala 30:58:@13126.4]
  wire [10:0] _T_914; // @[Cat.scala 30:58:@13128.4]
  wire [10:0] _T_916; // @[Cat.scala 30:58:@13130.4]
  wire [10:0] _T_918; // @[Cat.scala 30:58:@13132.4]
  wire [10:0] _T_920; // @[Cat.scala 30:58:@13134.4]
  wire [10:0] _T_921; // @[Mux.scala 31:69:@13135.4]
  wire [10:0] _T_922; // @[Mux.scala 31:69:@13136.4]
  wire [10:0] _T_923; // @[Mux.scala 31:69:@13137.4]
  wire [10:0] _T_924; // @[Mux.scala 31:69:@13138.4]
  wire [10:0] _T_925; // @[Mux.scala 31:69:@13139.4]
  wire  _T_930; // @[MemPrimitives.scala 110:210:@13146.4]
  wire  _T_933; // @[MemPrimitives.scala 110:228:@13148.4]
  wire  _T_936; // @[MemPrimitives.scala 110:210:@13150.4]
  wire  _T_939; // @[MemPrimitives.scala 110:228:@13152.4]
  wire  _T_942; // @[MemPrimitives.scala 110:210:@13154.4]
  wire  _T_945; // @[MemPrimitives.scala 110:228:@13156.4]
  wire  _T_948; // @[MemPrimitives.scala 110:210:@13158.4]
  wire  _T_951; // @[MemPrimitives.scala 110:228:@13160.4]
  wire  _T_954; // @[MemPrimitives.scala 110:210:@13162.4]
  wire  _T_957; // @[MemPrimitives.scala 110:228:@13164.4]
  wire  _T_960; // @[MemPrimitives.scala 110:210:@13166.4]
  wire  _T_963; // @[MemPrimitives.scala 110:228:@13168.4]
  wire  _T_965; // @[MemPrimitives.scala 126:35:@13179.4]
  wire  _T_966; // @[MemPrimitives.scala 126:35:@13180.4]
  wire  _T_967; // @[MemPrimitives.scala 126:35:@13181.4]
  wire  _T_968; // @[MemPrimitives.scala 126:35:@13182.4]
  wire  _T_969; // @[MemPrimitives.scala 126:35:@13183.4]
  wire  _T_970; // @[MemPrimitives.scala 126:35:@13184.4]
  wire [10:0] _T_972; // @[Cat.scala 30:58:@13186.4]
  wire [10:0] _T_974; // @[Cat.scala 30:58:@13188.4]
  wire [10:0] _T_976; // @[Cat.scala 30:58:@13190.4]
  wire [10:0] _T_978; // @[Cat.scala 30:58:@13192.4]
  wire [10:0] _T_980; // @[Cat.scala 30:58:@13194.4]
  wire [10:0] _T_982; // @[Cat.scala 30:58:@13196.4]
  wire [10:0] _T_983; // @[Mux.scala 31:69:@13197.4]
  wire [10:0] _T_984; // @[Mux.scala 31:69:@13198.4]
  wire [10:0] _T_985; // @[Mux.scala 31:69:@13199.4]
  wire [10:0] _T_986; // @[Mux.scala 31:69:@13200.4]
  wire [10:0] _T_987; // @[Mux.scala 31:69:@13201.4]
  wire  _T_995; // @[MemPrimitives.scala 110:228:@13210.4]
  wire  _T_1001; // @[MemPrimitives.scala 110:228:@13214.4]
  wire  _T_1007; // @[MemPrimitives.scala 110:228:@13218.4]
  wire  _T_1013; // @[MemPrimitives.scala 110:228:@13222.4]
  wire  _T_1019; // @[MemPrimitives.scala 110:228:@13226.4]
  wire  _T_1025; // @[MemPrimitives.scala 110:228:@13230.4]
  wire  _T_1027; // @[MemPrimitives.scala 126:35:@13241.4]
  wire  _T_1028; // @[MemPrimitives.scala 126:35:@13242.4]
  wire  _T_1029; // @[MemPrimitives.scala 126:35:@13243.4]
  wire  _T_1030; // @[MemPrimitives.scala 126:35:@13244.4]
  wire  _T_1031; // @[MemPrimitives.scala 126:35:@13245.4]
  wire  _T_1032; // @[MemPrimitives.scala 126:35:@13246.4]
  wire [10:0] _T_1034; // @[Cat.scala 30:58:@13248.4]
  wire [10:0] _T_1036; // @[Cat.scala 30:58:@13250.4]
  wire [10:0] _T_1038; // @[Cat.scala 30:58:@13252.4]
  wire [10:0] _T_1040; // @[Cat.scala 30:58:@13254.4]
  wire [10:0] _T_1042; // @[Cat.scala 30:58:@13256.4]
  wire [10:0] _T_1044; // @[Cat.scala 30:58:@13258.4]
  wire [10:0] _T_1045; // @[Mux.scala 31:69:@13259.4]
  wire [10:0] _T_1046; // @[Mux.scala 31:69:@13260.4]
  wire [10:0] _T_1047; // @[Mux.scala 31:69:@13261.4]
  wire [10:0] _T_1048; // @[Mux.scala 31:69:@13262.4]
  wire [10:0] _T_1049; // @[Mux.scala 31:69:@13263.4]
  wire  _T_1057; // @[MemPrimitives.scala 110:228:@13272.4]
  wire  _T_1063; // @[MemPrimitives.scala 110:228:@13276.4]
  wire  _T_1069; // @[MemPrimitives.scala 110:228:@13280.4]
  wire  _T_1075; // @[MemPrimitives.scala 110:228:@13284.4]
  wire  _T_1081; // @[MemPrimitives.scala 110:228:@13288.4]
  wire  _T_1087; // @[MemPrimitives.scala 110:228:@13292.4]
  wire  _T_1089; // @[MemPrimitives.scala 126:35:@13303.4]
  wire  _T_1090; // @[MemPrimitives.scala 126:35:@13304.4]
  wire  _T_1091; // @[MemPrimitives.scala 126:35:@13305.4]
  wire  _T_1092; // @[MemPrimitives.scala 126:35:@13306.4]
  wire  _T_1093; // @[MemPrimitives.scala 126:35:@13307.4]
  wire  _T_1094; // @[MemPrimitives.scala 126:35:@13308.4]
  wire [10:0] _T_1096; // @[Cat.scala 30:58:@13310.4]
  wire [10:0] _T_1098; // @[Cat.scala 30:58:@13312.4]
  wire [10:0] _T_1100; // @[Cat.scala 30:58:@13314.4]
  wire [10:0] _T_1102; // @[Cat.scala 30:58:@13316.4]
  wire [10:0] _T_1104; // @[Cat.scala 30:58:@13318.4]
  wire [10:0] _T_1106; // @[Cat.scala 30:58:@13320.4]
  wire [10:0] _T_1107; // @[Mux.scala 31:69:@13321.4]
  wire [10:0] _T_1108; // @[Mux.scala 31:69:@13322.4]
  wire [10:0] _T_1109; // @[Mux.scala 31:69:@13323.4]
  wire [10:0] _T_1110; // @[Mux.scala 31:69:@13324.4]
  wire [10:0] _T_1111; // @[Mux.scala 31:69:@13325.4]
  wire  _T_1116; // @[MemPrimitives.scala 110:210:@13332.4]
  wire  _T_1119; // @[MemPrimitives.scala 110:228:@13334.4]
  wire  _T_1122; // @[MemPrimitives.scala 110:210:@13336.4]
  wire  _T_1125; // @[MemPrimitives.scala 110:228:@13338.4]
  wire  _T_1128; // @[MemPrimitives.scala 110:210:@13340.4]
  wire  _T_1131; // @[MemPrimitives.scala 110:228:@13342.4]
  wire  _T_1134; // @[MemPrimitives.scala 110:210:@13344.4]
  wire  _T_1137; // @[MemPrimitives.scala 110:228:@13346.4]
  wire  _T_1140; // @[MemPrimitives.scala 110:210:@13348.4]
  wire  _T_1143; // @[MemPrimitives.scala 110:228:@13350.4]
  wire  _T_1146; // @[MemPrimitives.scala 110:210:@13352.4]
  wire  _T_1149; // @[MemPrimitives.scala 110:228:@13354.4]
  wire  _T_1151; // @[MemPrimitives.scala 126:35:@13365.4]
  wire  _T_1152; // @[MemPrimitives.scala 126:35:@13366.4]
  wire  _T_1153; // @[MemPrimitives.scala 126:35:@13367.4]
  wire  _T_1154; // @[MemPrimitives.scala 126:35:@13368.4]
  wire  _T_1155; // @[MemPrimitives.scala 126:35:@13369.4]
  wire  _T_1156; // @[MemPrimitives.scala 126:35:@13370.4]
  wire [10:0] _T_1158; // @[Cat.scala 30:58:@13372.4]
  wire [10:0] _T_1160; // @[Cat.scala 30:58:@13374.4]
  wire [10:0] _T_1162; // @[Cat.scala 30:58:@13376.4]
  wire [10:0] _T_1164; // @[Cat.scala 30:58:@13378.4]
  wire [10:0] _T_1166; // @[Cat.scala 30:58:@13380.4]
  wire [10:0] _T_1168; // @[Cat.scala 30:58:@13382.4]
  wire [10:0] _T_1169; // @[Mux.scala 31:69:@13383.4]
  wire [10:0] _T_1170; // @[Mux.scala 31:69:@13384.4]
  wire [10:0] _T_1171; // @[Mux.scala 31:69:@13385.4]
  wire [10:0] _T_1172; // @[Mux.scala 31:69:@13386.4]
  wire [10:0] _T_1173; // @[Mux.scala 31:69:@13387.4]
  wire  _T_1178; // @[MemPrimitives.scala 110:210:@13394.4]
  wire  _T_1181; // @[MemPrimitives.scala 110:228:@13396.4]
  wire  _T_1184; // @[MemPrimitives.scala 110:210:@13398.4]
  wire  _T_1187; // @[MemPrimitives.scala 110:228:@13400.4]
  wire  _T_1190; // @[MemPrimitives.scala 110:210:@13402.4]
  wire  _T_1193; // @[MemPrimitives.scala 110:228:@13404.4]
  wire  _T_1196; // @[MemPrimitives.scala 110:210:@13406.4]
  wire  _T_1199; // @[MemPrimitives.scala 110:228:@13408.4]
  wire  _T_1202; // @[MemPrimitives.scala 110:210:@13410.4]
  wire  _T_1205; // @[MemPrimitives.scala 110:228:@13412.4]
  wire  _T_1208; // @[MemPrimitives.scala 110:210:@13414.4]
  wire  _T_1211; // @[MemPrimitives.scala 110:228:@13416.4]
  wire  _T_1213; // @[MemPrimitives.scala 126:35:@13427.4]
  wire  _T_1214; // @[MemPrimitives.scala 126:35:@13428.4]
  wire  _T_1215; // @[MemPrimitives.scala 126:35:@13429.4]
  wire  _T_1216; // @[MemPrimitives.scala 126:35:@13430.4]
  wire  _T_1217; // @[MemPrimitives.scala 126:35:@13431.4]
  wire  _T_1218; // @[MemPrimitives.scala 126:35:@13432.4]
  wire [10:0] _T_1220; // @[Cat.scala 30:58:@13434.4]
  wire [10:0] _T_1222; // @[Cat.scala 30:58:@13436.4]
  wire [10:0] _T_1224; // @[Cat.scala 30:58:@13438.4]
  wire [10:0] _T_1226; // @[Cat.scala 30:58:@13440.4]
  wire [10:0] _T_1228; // @[Cat.scala 30:58:@13442.4]
  wire [10:0] _T_1230; // @[Cat.scala 30:58:@13444.4]
  wire [10:0] _T_1231; // @[Mux.scala 31:69:@13445.4]
  wire [10:0] _T_1232; // @[Mux.scala 31:69:@13446.4]
  wire [10:0] _T_1233; // @[Mux.scala 31:69:@13447.4]
  wire [10:0] _T_1234; // @[Mux.scala 31:69:@13448.4]
  wire [10:0] _T_1235; // @[Mux.scala 31:69:@13449.4]
  wire  _T_1243; // @[MemPrimitives.scala 110:228:@13458.4]
  wire  _T_1249; // @[MemPrimitives.scala 110:228:@13462.4]
  wire  _T_1255; // @[MemPrimitives.scala 110:228:@13466.4]
  wire  _T_1261; // @[MemPrimitives.scala 110:228:@13470.4]
  wire  _T_1267; // @[MemPrimitives.scala 110:228:@13474.4]
  wire  _T_1273; // @[MemPrimitives.scala 110:228:@13478.4]
  wire  _T_1275; // @[MemPrimitives.scala 126:35:@13489.4]
  wire  _T_1276; // @[MemPrimitives.scala 126:35:@13490.4]
  wire  _T_1277; // @[MemPrimitives.scala 126:35:@13491.4]
  wire  _T_1278; // @[MemPrimitives.scala 126:35:@13492.4]
  wire  _T_1279; // @[MemPrimitives.scala 126:35:@13493.4]
  wire  _T_1280; // @[MemPrimitives.scala 126:35:@13494.4]
  wire [10:0] _T_1282; // @[Cat.scala 30:58:@13496.4]
  wire [10:0] _T_1284; // @[Cat.scala 30:58:@13498.4]
  wire [10:0] _T_1286; // @[Cat.scala 30:58:@13500.4]
  wire [10:0] _T_1288; // @[Cat.scala 30:58:@13502.4]
  wire [10:0] _T_1290; // @[Cat.scala 30:58:@13504.4]
  wire [10:0] _T_1292; // @[Cat.scala 30:58:@13506.4]
  wire [10:0] _T_1293; // @[Mux.scala 31:69:@13507.4]
  wire [10:0] _T_1294; // @[Mux.scala 31:69:@13508.4]
  wire [10:0] _T_1295; // @[Mux.scala 31:69:@13509.4]
  wire [10:0] _T_1296; // @[Mux.scala 31:69:@13510.4]
  wire [10:0] _T_1297; // @[Mux.scala 31:69:@13511.4]
  wire  _T_1305; // @[MemPrimitives.scala 110:228:@13520.4]
  wire  _T_1311; // @[MemPrimitives.scala 110:228:@13524.4]
  wire  _T_1317; // @[MemPrimitives.scala 110:228:@13528.4]
  wire  _T_1323; // @[MemPrimitives.scala 110:228:@13532.4]
  wire  _T_1329; // @[MemPrimitives.scala 110:228:@13536.4]
  wire  _T_1335; // @[MemPrimitives.scala 110:228:@13540.4]
  wire  _T_1337; // @[MemPrimitives.scala 126:35:@13551.4]
  wire  _T_1338; // @[MemPrimitives.scala 126:35:@13552.4]
  wire  _T_1339; // @[MemPrimitives.scala 126:35:@13553.4]
  wire  _T_1340; // @[MemPrimitives.scala 126:35:@13554.4]
  wire  _T_1341; // @[MemPrimitives.scala 126:35:@13555.4]
  wire  _T_1342; // @[MemPrimitives.scala 126:35:@13556.4]
  wire [10:0] _T_1344; // @[Cat.scala 30:58:@13558.4]
  wire [10:0] _T_1346; // @[Cat.scala 30:58:@13560.4]
  wire [10:0] _T_1348; // @[Cat.scala 30:58:@13562.4]
  wire [10:0] _T_1350; // @[Cat.scala 30:58:@13564.4]
  wire [10:0] _T_1352; // @[Cat.scala 30:58:@13566.4]
  wire [10:0] _T_1354; // @[Cat.scala 30:58:@13568.4]
  wire [10:0] _T_1355; // @[Mux.scala 31:69:@13569.4]
  wire [10:0] _T_1356; // @[Mux.scala 31:69:@13570.4]
  wire [10:0] _T_1357; // @[Mux.scala 31:69:@13571.4]
  wire [10:0] _T_1358; // @[Mux.scala 31:69:@13572.4]
  wire [10:0] _T_1359; // @[Mux.scala 31:69:@13573.4]
  wire  _T_1364; // @[MemPrimitives.scala 110:210:@13580.4]
  wire  _T_1367; // @[MemPrimitives.scala 110:228:@13582.4]
  wire  _T_1370; // @[MemPrimitives.scala 110:210:@13584.4]
  wire  _T_1373; // @[MemPrimitives.scala 110:228:@13586.4]
  wire  _T_1376; // @[MemPrimitives.scala 110:210:@13588.4]
  wire  _T_1379; // @[MemPrimitives.scala 110:228:@13590.4]
  wire  _T_1382; // @[MemPrimitives.scala 110:210:@13592.4]
  wire  _T_1385; // @[MemPrimitives.scala 110:228:@13594.4]
  wire  _T_1388; // @[MemPrimitives.scala 110:210:@13596.4]
  wire  _T_1391; // @[MemPrimitives.scala 110:228:@13598.4]
  wire  _T_1394; // @[MemPrimitives.scala 110:210:@13600.4]
  wire  _T_1397; // @[MemPrimitives.scala 110:228:@13602.4]
  wire  _T_1399; // @[MemPrimitives.scala 126:35:@13613.4]
  wire  _T_1400; // @[MemPrimitives.scala 126:35:@13614.4]
  wire  _T_1401; // @[MemPrimitives.scala 126:35:@13615.4]
  wire  _T_1402; // @[MemPrimitives.scala 126:35:@13616.4]
  wire  _T_1403; // @[MemPrimitives.scala 126:35:@13617.4]
  wire  _T_1404; // @[MemPrimitives.scala 126:35:@13618.4]
  wire [10:0] _T_1406; // @[Cat.scala 30:58:@13620.4]
  wire [10:0] _T_1408; // @[Cat.scala 30:58:@13622.4]
  wire [10:0] _T_1410; // @[Cat.scala 30:58:@13624.4]
  wire [10:0] _T_1412; // @[Cat.scala 30:58:@13626.4]
  wire [10:0] _T_1414; // @[Cat.scala 30:58:@13628.4]
  wire [10:0] _T_1416; // @[Cat.scala 30:58:@13630.4]
  wire [10:0] _T_1417; // @[Mux.scala 31:69:@13631.4]
  wire [10:0] _T_1418; // @[Mux.scala 31:69:@13632.4]
  wire [10:0] _T_1419; // @[Mux.scala 31:69:@13633.4]
  wire [10:0] _T_1420; // @[Mux.scala 31:69:@13634.4]
  wire [10:0] _T_1421; // @[Mux.scala 31:69:@13635.4]
  wire  _T_1426; // @[MemPrimitives.scala 110:210:@13642.4]
  wire  _T_1429; // @[MemPrimitives.scala 110:228:@13644.4]
  wire  _T_1432; // @[MemPrimitives.scala 110:210:@13646.4]
  wire  _T_1435; // @[MemPrimitives.scala 110:228:@13648.4]
  wire  _T_1438; // @[MemPrimitives.scala 110:210:@13650.4]
  wire  _T_1441; // @[MemPrimitives.scala 110:228:@13652.4]
  wire  _T_1444; // @[MemPrimitives.scala 110:210:@13654.4]
  wire  _T_1447; // @[MemPrimitives.scala 110:228:@13656.4]
  wire  _T_1450; // @[MemPrimitives.scala 110:210:@13658.4]
  wire  _T_1453; // @[MemPrimitives.scala 110:228:@13660.4]
  wire  _T_1456; // @[MemPrimitives.scala 110:210:@13662.4]
  wire  _T_1459; // @[MemPrimitives.scala 110:228:@13664.4]
  wire  _T_1461; // @[MemPrimitives.scala 126:35:@13675.4]
  wire  _T_1462; // @[MemPrimitives.scala 126:35:@13676.4]
  wire  _T_1463; // @[MemPrimitives.scala 126:35:@13677.4]
  wire  _T_1464; // @[MemPrimitives.scala 126:35:@13678.4]
  wire  _T_1465; // @[MemPrimitives.scala 126:35:@13679.4]
  wire  _T_1466; // @[MemPrimitives.scala 126:35:@13680.4]
  wire [10:0] _T_1468; // @[Cat.scala 30:58:@13682.4]
  wire [10:0] _T_1470; // @[Cat.scala 30:58:@13684.4]
  wire [10:0] _T_1472; // @[Cat.scala 30:58:@13686.4]
  wire [10:0] _T_1474; // @[Cat.scala 30:58:@13688.4]
  wire [10:0] _T_1476; // @[Cat.scala 30:58:@13690.4]
  wire [10:0] _T_1478; // @[Cat.scala 30:58:@13692.4]
  wire [10:0] _T_1479; // @[Mux.scala 31:69:@13693.4]
  wire [10:0] _T_1480; // @[Mux.scala 31:69:@13694.4]
  wire [10:0] _T_1481; // @[Mux.scala 31:69:@13695.4]
  wire [10:0] _T_1482; // @[Mux.scala 31:69:@13696.4]
  wire [10:0] _T_1483; // @[Mux.scala 31:69:@13697.4]
  wire  _T_1491; // @[MemPrimitives.scala 110:228:@13706.4]
  wire  _T_1497; // @[MemPrimitives.scala 110:228:@13710.4]
  wire  _T_1503; // @[MemPrimitives.scala 110:228:@13714.4]
  wire  _T_1509; // @[MemPrimitives.scala 110:228:@13718.4]
  wire  _T_1515; // @[MemPrimitives.scala 110:228:@13722.4]
  wire  _T_1521; // @[MemPrimitives.scala 110:228:@13726.4]
  wire  _T_1523; // @[MemPrimitives.scala 126:35:@13737.4]
  wire  _T_1524; // @[MemPrimitives.scala 126:35:@13738.4]
  wire  _T_1525; // @[MemPrimitives.scala 126:35:@13739.4]
  wire  _T_1526; // @[MemPrimitives.scala 126:35:@13740.4]
  wire  _T_1527; // @[MemPrimitives.scala 126:35:@13741.4]
  wire  _T_1528; // @[MemPrimitives.scala 126:35:@13742.4]
  wire [10:0] _T_1530; // @[Cat.scala 30:58:@13744.4]
  wire [10:0] _T_1532; // @[Cat.scala 30:58:@13746.4]
  wire [10:0] _T_1534; // @[Cat.scala 30:58:@13748.4]
  wire [10:0] _T_1536; // @[Cat.scala 30:58:@13750.4]
  wire [10:0] _T_1538; // @[Cat.scala 30:58:@13752.4]
  wire [10:0] _T_1540; // @[Cat.scala 30:58:@13754.4]
  wire [10:0] _T_1541; // @[Mux.scala 31:69:@13755.4]
  wire [10:0] _T_1542; // @[Mux.scala 31:69:@13756.4]
  wire [10:0] _T_1543; // @[Mux.scala 31:69:@13757.4]
  wire [10:0] _T_1544; // @[Mux.scala 31:69:@13758.4]
  wire [10:0] _T_1545; // @[Mux.scala 31:69:@13759.4]
  wire  _T_1553; // @[MemPrimitives.scala 110:228:@13768.4]
  wire  _T_1559; // @[MemPrimitives.scala 110:228:@13772.4]
  wire  _T_1565; // @[MemPrimitives.scala 110:228:@13776.4]
  wire  _T_1571; // @[MemPrimitives.scala 110:228:@13780.4]
  wire  _T_1577; // @[MemPrimitives.scala 110:228:@13784.4]
  wire  _T_1583; // @[MemPrimitives.scala 110:228:@13788.4]
  wire  _T_1585; // @[MemPrimitives.scala 126:35:@13799.4]
  wire  _T_1586; // @[MemPrimitives.scala 126:35:@13800.4]
  wire  _T_1587; // @[MemPrimitives.scala 126:35:@13801.4]
  wire  _T_1588; // @[MemPrimitives.scala 126:35:@13802.4]
  wire  _T_1589; // @[MemPrimitives.scala 126:35:@13803.4]
  wire  _T_1590; // @[MemPrimitives.scala 126:35:@13804.4]
  wire [10:0] _T_1592; // @[Cat.scala 30:58:@13806.4]
  wire [10:0] _T_1594; // @[Cat.scala 30:58:@13808.4]
  wire [10:0] _T_1596; // @[Cat.scala 30:58:@13810.4]
  wire [10:0] _T_1598; // @[Cat.scala 30:58:@13812.4]
  wire [10:0] _T_1600; // @[Cat.scala 30:58:@13814.4]
  wire [10:0] _T_1602; // @[Cat.scala 30:58:@13816.4]
  wire [10:0] _T_1603; // @[Mux.scala 31:69:@13817.4]
  wire [10:0] _T_1604; // @[Mux.scala 31:69:@13818.4]
  wire [10:0] _T_1605; // @[Mux.scala 31:69:@13819.4]
  wire [10:0] _T_1606; // @[Mux.scala 31:69:@13820.4]
  wire [10:0] _T_1607; // @[Mux.scala 31:69:@13821.4]
  wire  _T_1671; // @[package.scala 96:25:@13906.4 package.scala 96:25:@13907.4]
  wire [31:0] _T_1675; // @[Mux.scala 31:69:@13916.4]
  wire  _T_1668; // @[package.scala 96:25:@13898.4 package.scala 96:25:@13899.4]
  wire [31:0] _T_1676; // @[Mux.scala 31:69:@13917.4]
  wire  _T_1665; // @[package.scala 96:25:@13890.4 package.scala 96:25:@13891.4]
  wire [31:0] _T_1677; // @[Mux.scala 31:69:@13918.4]
  wire  _T_1662; // @[package.scala 96:25:@13882.4 package.scala 96:25:@13883.4]
  wire [31:0] _T_1678; // @[Mux.scala 31:69:@13919.4]
  wire  _T_1659; // @[package.scala 96:25:@13874.4 package.scala 96:25:@13875.4]
  wire [31:0] _T_1679; // @[Mux.scala 31:69:@13920.4]
  wire  _T_1656; // @[package.scala 96:25:@13866.4 package.scala 96:25:@13867.4]
  wire [31:0] _T_1680; // @[Mux.scala 31:69:@13921.4]
  wire  _T_1653; // @[package.scala 96:25:@13858.4 package.scala 96:25:@13859.4]
  wire  _T_1742; // @[package.scala 96:25:@14002.4 package.scala 96:25:@14003.4]
  wire [31:0] _T_1746; // @[Mux.scala 31:69:@14012.4]
  wire  _T_1739; // @[package.scala 96:25:@13994.4 package.scala 96:25:@13995.4]
  wire [31:0] _T_1747; // @[Mux.scala 31:69:@14013.4]
  wire  _T_1736; // @[package.scala 96:25:@13986.4 package.scala 96:25:@13987.4]
  wire [31:0] _T_1748; // @[Mux.scala 31:69:@14014.4]
  wire  _T_1733; // @[package.scala 96:25:@13978.4 package.scala 96:25:@13979.4]
  wire [31:0] _T_1749; // @[Mux.scala 31:69:@14015.4]
  wire  _T_1730; // @[package.scala 96:25:@13970.4 package.scala 96:25:@13971.4]
  wire [31:0] _T_1750; // @[Mux.scala 31:69:@14016.4]
  wire  _T_1727; // @[package.scala 96:25:@13962.4 package.scala 96:25:@13963.4]
  wire [31:0] _T_1751; // @[Mux.scala 31:69:@14017.4]
  wire  _T_1724; // @[package.scala 96:25:@13954.4 package.scala 96:25:@13955.4]
  wire  _T_1813; // @[package.scala 96:25:@14098.4 package.scala 96:25:@14099.4]
  wire [31:0] _T_1817; // @[Mux.scala 31:69:@14108.4]
  wire  _T_1810; // @[package.scala 96:25:@14090.4 package.scala 96:25:@14091.4]
  wire [31:0] _T_1818; // @[Mux.scala 31:69:@14109.4]
  wire  _T_1807; // @[package.scala 96:25:@14082.4 package.scala 96:25:@14083.4]
  wire [31:0] _T_1819; // @[Mux.scala 31:69:@14110.4]
  wire  _T_1804; // @[package.scala 96:25:@14074.4 package.scala 96:25:@14075.4]
  wire [31:0] _T_1820; // @[Mux.scala 31:69:@14111.4]
  wire  _T_1801; // @[package.scala 96:25:@14066.4 package.scala 96:25:@14067.4]
  wire [31:0] _T_1821; // @[Mux.scala 31:69:@14112.4]
  wire  _T_1798; // @[package.scala 96:25:@14058.4 package.scala 96:25:@14059.4]
  wire [31:0] _T_1822; // @[Mux.scala 31:69:@14113.4]
  wire  _T_1795; // @[package.scala 96:25:@14050.4 package.scala 96:25:@14051.4]
  wire  _T_1884; // @[package.scala 96:25:@14194.4 package.scala 96:25:@14195.4]
  wire [31:0] _T_1888; // @[Mux.scala 31:69:@14204.4]
  wire  _T_1881; // @[package.scala 96:25:@14186.4 package.scala 96:25:@14187.4]
  wire [31:0] _T_1889; // @[Mux.scala 31:69:@14205.4]
  wire  _T_1878; // @[package.scala 96:25:@14178.4 package.scala 96:25:@14179.4]
  wire [31:0] _T_1890; // @[Mux.scala 31:69:@14206.4]
  wire  _T_1875; // @[package.scala 96:25:@14170.4 package.scala 96:25:@14171.4]
  wire [31:0] _T_1891; // @[Mux.scala 31:69:@14207.4]
  wire  _T_1872; // @[package.scala 96:25:@14162.4 package.scala 96:25:@14163.4]
  wire [31:0] _T_1892; // @[Mux.scala 31:69:@14208.4]
  wire  _T_1869; // @[package.scala 96:25:@14154.4 package.scala 96:25:@14155.4]
  wire [31:0] _T_1893; // @[Mux.scala 31:69:@14209.4]
  wire  _T_1866; // @[package.scala 96:25:@14146.4 package.scala 96:25:@14147.4]
  wire  _T_1955; // @[package.scala 96:25:@14290.4 package.scala 96:25:@14291.4]
  wire [31:0] _T_1959; // @[Mux.scala 31:69:@14300.4]
  wire  _T_1952; // @[package.scala 96:25:@14282.4 package.scala 96:25:@14283.4]
  wire [31:0] _T_1960; // @[Mux.scala 31:69:@14301.4]
  wire  _T_1949; // @[package.scala 96:25:@14274.4 package.scala 96:25:@14275.4]
  wire [31:0] _T_1961; // @[Mux.scala 31:69:@14302.4]
  wire  _T_1946; // @[package.scala 96:25:@14266.4 package.scala 96:25:@14267.4]
  wire [31:0] _T_1962; // @[Mux.scala 31:69:@14303.4]
  wire  _T_1943; // @[package.scala 96:25:@14258.4 package.scala 96:25:@14259.4]
  wire [31:0] _T_1963; // @[Mux.scala 31:69:@14304.4]
  wire  _T_1940; // @[package.scala 96:25:@14250.4 package.scala 96:25:@14251.4]
  wire [31:0] _T_1964; // @[Mux.scala 31:69:@14305.4]
  wire  _T_1937; // @[package.scala 96:25:@14242.4 package.scala 96:25:@14243.4]
  wire  _T_2026; // @[package.scala 96:25:@14386.4 package.scala 96:25:@14387.4]
  wire [31:0] _T_2030; // @[Mux.scala 31:69:@14396.4]
  wire  _T_2023; // @[package.scala 96:25:@14378.4 package.scala 96:25:@14379.4]
  wire [31:0] _T_2031; // @[Mux.scala 31:69:@14397.4]
  wire  _T_2020; // @[package.scala 96:25:@14370.4 package.scala 96:25:@14371.4]
  wire [31:0] _T_2032; // @[Mux.scala 31:69:@14398.4]
  wire  _T_2017; // @[package.scala 96:25:@14362.4 package.scala 96:25:@14363.4]
  wire [31:0] _T_2033; // @[Mux.scala 31:69:@14399.4]
  wire  _T_2014; // @[package.scala 96:25:@14354.4 package.scala 96:25:@14355.4]
  wire [31:0] _T_2034; // @[Mux.scala 31:69:@14400.4]
  wire  _T_2011; // @[package.scala 96:25:@14346.4 package.scala 96:25:@14347.4]
  wire [31:0] _T_2035; // @[Mux.scala 31:69:@14401.4]
  wire  _T_2008; // @[package.scala 96:25:@14338.4 package.scala 96:25:@14339.4]
  wire  _T_2097; // @[package.scala 96:25:@14482.4 package.scala 96:25:@14483.4]
  wire [31:0] _T_2101; // @[Mux.scala 31:69:@14492.4]
  wire  _T_2094; // @[package.scala 96:25:@14474.4 package.scala 96:25:@14475.4]
  wire [31:0] _T_2102; // @[Mux.scala 31:69:@14493.4]
  wire  _T_2091; // @[package.scala 96:25:@14466.4 package.scala 96:25:@14467.4]
  wire [31:0] _T_2103; // @[Mux.scala 31:69:@14494.4]
  wire  _T_2088; // @[package.scala 96:25:@14458.4 package.scala 96:25:@14459.4]
  wire [31:0] _T_2104; // @[Mux.scala 31:69:@14495.4]
  wire  _T_2085; // @[package.scala 96:25:@14450.4 package.scala 96:25:@14451.4]
  wire [31:0] _T_2105; // @[Mux.scala 31:69:@14496.4]
  wire  _T_2082; // @[package.scala 96:25:@14442.4 package.scala 96:25:@14443.4]
  wire [31:0] _T_2106; // @[Mux.scala 31:69:@14497.4]
  wire  _T_2079; // @[package.scala 96:25:@14434.4 package.scala 96:25:@14435.4]
  wire  _T_2168; // @[package.scala 96:25:@14578.4 package.scala 96:25:@14579.4]
  wire [31:0] _T_2172; // @[Mux.scala 31:69:@14588.4]
  wire  _T_2165; // @[package.scala 96:25:@14570.4 package.scala 96:25:@14571.4]
  wire [31:0] _T_2173; // @[Mux.scala 31:69:@14589.4]
  wire  _T_2162; // @[package.scala 96:25:@14562.4 package.scala 96:25:@14563.4]
  wire [31:0] _T_2174; // @[Mux.scala 31:69:@14590.4]
  wire  _T_2159; // @[package.scala 96:25:@14554.4 package.scala 96:25:@14555.4]
  wire [31:0] _T_2175; // @[Mux.scala 31:69:@14591.4]
  wire  _T_2156; // @[package.scala 96:25:@14546.4 package.scala 96:25:@14547.4]
  wire [31:0] _T_2176; // @[Mux.scala 31:69:@14592.4]
  wire  _T_2153; // @[package.scala 96:25:@14538.4 package.scala 96:25:@14539.4]
  wire [31:0] _T_2177; // @[Mux.scala 31:69:@14593.4]
  wire  _T_2150; // @[package.scala 96:25:@14530.4 package.scala 96:25:@14531.4]
  wire  _T_2239; // @[package.scala 96:25:@14674.4 package.scala 96:25:@14675.4]
  wire [31:0] _T_2243; // @[Mux.scala 31:69:@14684.4]
  wire  _T_2236; // @[package.scala 96:25:@14666.4 package.scala 96:25:@14667.4]
  wire [31:0] _T_2244; // @[Mux.scala 31:69:@14685.4]
  wire  _T_2233; // @[package.scala 96:25:@14658.4 package.scala 96:25:@14659.4]
  wire [31:0] _T_2245; // @[Mux.scala 31:69:@14686.4]
  wire  _T_2230; // @[package.scala 96:25:@14650.4 package.scala 96:25:@14651.4]
  wire [31:0] _T_2246; // @[Mux.scala 31:69:@14687.4]
  wire  _T_2227; // @[package.scala 96:25:@14642.4 package.scala 96:25:@14643.4]
  wire [31:0] _T_2247; // @[Mux.scala 31:69:@14688.4]
  wire  _T_2224; // @[package.scala 96:25:@14634.4 package.scala 96:25:@14635.4]
  wire [31:0] _T_2248; // @[Mux.scala 31:69:@14689.4]
  wire  _T_2221; // @[package.scala 96:25:@14626.4 package.scala 96:25:@14627.4]
  wire  _T_2310; // @[package.scala 96:25:@14770.4 package.scala 96:25:@14771.4]
  wire [31:0] _T_2314; // @[Mux.scala 31:69:@14780.4]
  wire  _T_2307; // @[package.scala 96:25:@14762.4 package.scala 96:25:@14763.4]
  wire [31:0] _T_2315; // @[Mux.scala 31:69:@14781.4]
  wire  _T_2304; // @[package.scala 96:25:@14754.4 package.scala 96:25:@14755.4]
  wire [31:0] _T_2316; // @[Mux.scala 31:69:@14782.4]
  wire  _T_2301; // @[package.scala 96:25:@14746.4 package.scala 96:25:@14747.4]
  wire [31:0] _T_2317; // @[Mux.scala 31:69:@14783.4]
  wire  _T_2298; // @[package.scala 96:25:@14738.4 package.scala 96:25:@14739.4]
  wire [31:0] _T_2318; // @[Mux.scala 31:69:@14784.4]
  wire  _T_2295; // @[package.scala 96:25:@14730.4 package.scala 96:25:@14731.4]
  wire [31:0] _T_2319; // @[Mux.scala 31:69:@14785.4]
  wire  _T_2292; // @[package.scala 96:25:@14722.4 package.scala 96:25:@14723.4]
  wire  _T_2381; // @[package.scala 96:25:@14866.4 package.scala 96:25:@14867.4]
  wire [31:0] _T_2385; // @[Mux.scala 31:69:@14876.4]
  wire  _T_2378; // @[package.scala 96:25:@14858.4 package.scala 96:25:@14859.4]
  wire [31:0] _T_2386; // @[Mux.scala 31:69:@14877.4]
  wire  _T_2375; // @[package.scala 96:25:@14850.4 package.scala 96:25:@14851.4]
  wire [31:0] _T_2387; // @[Mux.scala 31:69:@14878.4]
  wire  _T_2372; // @[package.scala 96:25:@14842.4 package.scala 96:25:@14843.4]
  wire [31:0] _T_2388; // @[Mux.scala 31:69:@14879.4]
  wire  _T_2369; // @[package.scala 96:25:@14834.4 package.scala 96:25:@14835.4]
  wire [31:0] _T_2389; // @[Mux.scala 31:69:@14880.4]
  wire  _T_2366; // @[package.scala 96:25:@14826.4 package.scala 96:25:@14827.4]
  wire [31:0] _T_2390; // @[Mux.scala 31:69:@14881.4]
  wire  _T_2363; // @[package.scala 96:25:@14818.4 package.scala 96:25:@14819.4]
  wire  _T_2452; // @[package.scala 96:25:@14962.4 package.scala 96:25:@14963.4]
  wire [31:0] _T_2456; // @[Mux.scala 31:69:@14972.4]
  wire  _T_2449; // @[package.scala 96:25:@14954.4 package.scala 96:25:@14955.4]
  wire [31:0] _T_2457; // @[Mux.scala 31:69:@14973.4]
  wire  _T_2446; // @[package.scala 96:25:@14946.4 package.scala 96:25:@14947.4]
  wire [31:0] _T_2458; // @[Mux.scala 31:69:@14974.4]
  wire  _T_2443; // @[package.scala 96:25:@14938.4 package.scala 96:25:@14939.4]
  wire [31:0] _T_2459; // @[Mux.scala 31:69:@14975.4]
  wire  _T_2440; // @[package.scala 96:25:@14930.4 package.scala 96:25:@14931.4]
  wire [31:0] _T_2460; // @[Mux.scala 31:69:@14976.4]
  wire  _T_2437; // @[package.scala 96:25:@14922.4 package.scala 96:25:@14923.4]
  wire [31:0] _T_2461; // @[Mux.scala 31:69:@14977.4]
  wire  _T_2434; // @[package.scala 96:25:@14914.4 package.scala 96:25:@14915.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@12388.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@12404.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@12420.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@12436.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@12452.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@12468.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@12484.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@12500.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@12516.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@12532.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@12548.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@12564.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_5 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@12580.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_5 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@12596.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_5 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@12612.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_5 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@12628.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects_1 StickySelects ( // @[MemPrimitives.scala 124:33:@12860.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5)
  );
  StickySelects_1 StickySelects_1 ( // @[MemPrimitives.scala 124:33:@12922.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5)
  );
  StickySelects_1 StickySelects_2 ( // @[MemPrimitives.scala 124:33:@12984.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5)
  );
  StickySelects_1 StickySelects_3 ( // @[MemPrimitives.scala 124:33:@13046.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5)
  );
  StickySelects_1 StickySelects_4 ( // @[MemPrimitives.scala 124:33:@13108.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5)
  );
  StickySelects_1 StickySelects_5 ( // @[MemPrimitives.scala 124:33:@13170.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5)
  );
  StickySelects_1 StickySelects_6 ( // @[MemPrimitives.scala 124:33:@13232.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5)
  );
  StickySelects_1 StickySelects_7 ( // @[MemPrimitives.scala 124:33:@13294.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5)
  );
  StickySelects_1 StickySelects_8 ( // @[MemPrimitives.scala 124:33:@13356.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5)
  );
  StickySelects_1 StickySelects_9 ( // @[MemPrimitives.scala 124:33:@13418.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5)
  );
  StickySelects_1 StickySelects_10 ( // @[MemPrimitives.scala 124:33:@13480.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5)
  );
  StickySelects_1 StickySelects_11 ( // @[MemPrimitives.scala 124:33:@13542.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5)
  );
  StickySelects_1 StickySelects_12 ( // @[MemPrimitives.scala 124:33:@13604.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_ins_4(StickySelects_12_io_ins_4),
    .io_ins_5(StickySelects_12_io_ins_5),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3),
    .io_outs_4(StickySelects_12_io_outs_4),
    .io_outs_5(StickySelects_12_io_outs_5)
  );
  StickySelects_1 StickySelects_13 ( // @[MemPrimitives.scala 124:33:@13666.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_ins_4(StickySelects_13_io_ins_4),
    .io_ins_5(StickySelects_13_io_ins_5),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3),
    .io_outs_4(StickySelects_13_io_outs_4),
    .io_outs_5(StickySelects_13_io_outs_5)
  );
  StickySelects_1 StickySelects_14 ( // @[MemPrimitives.scala 124:33:@13728.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5)
  );
  StickySelects_1 StickySelects_15 ( // @[MemPrimitives.scala 124:33:@13790.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@13853.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@13861.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@13869.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@13877.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@13885.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@13893.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@13901.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@13909.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@13949.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@13957.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@13965.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@13973.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@13981.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@13989.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@13997.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@14005.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@14045.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@14053.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@14061.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@14069.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@14077.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@14085.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@14093.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@14101.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@14141.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@14149.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@14157.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@14165.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@14173.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@14181.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@14189.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@14197.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@14237.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@14245.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@14253.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@14261.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@14269.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@14277.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@14285.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@14293.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@14333.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@14341.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@14349.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@14357.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@14365.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@14373.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@14381.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@14389.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_48 ( // @[package.scala 93:22:@14429.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@14437.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_50 ( // @[package.scala 93:22:@14445.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@14453.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@14461.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_53 ( // @[package.scala 93:22:@14469.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@14477.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_55 ( // @[package.scala 93:22:@14485.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@14525.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_57 ( // @[package.scala 93:22:@14533.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@14541.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_59 ( // @[package.scala 93:22:@14549.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_60 ( // @[package.scala 93:22:@14557.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_61 ( // @[package.scala 93:22:@14565.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_62 ( // @[package.scala 93:22:@14573.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_63 ( // @[package.scala 93:22:@14581.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_64 ( // @[package.scala 93:22:@14621.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_65 ( // @[package.scala 93:22:@14629.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_66 ( // @[package.scala 93:22:@14637.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_67 ( // @[package.scala 93:22:@14645.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_68 ( // @[package.scala 93:22:@14653.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_69 ( // @[package.scala 93:22:@14661.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_70 ( // @[package.scala 93:22:@14669.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_71 ( // @[package.scala 93:22:@14677.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_72 ( // @[package.scala 93:22:@14717.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_73 ( // @[package.scala 93:22:@14725.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_74 ( // @[package.scala 93:22:@14733.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_75 ( // @[package.scala 93:22:@14741.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_76 ( // @[package.scala 93:22:@14749.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_77 ( // @[package.scala 93:22:@14757.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_78 ( // @[package.scala 93:22:@14765.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_79 ( // @[package.scala 93:22:@14773.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_80 ( // @[package.scala 93:22:@14813.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_81 ( // @[package.scala 93:22:@14821.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_82 ( // @[package.scala 93:22:@14829.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_83 ( // @[package.scala 93:22:@14837.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_84 ( // @[package.scala 93:22:@14845.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_85 ( // @[package.scala 93:22:@14853.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_86 ( // @[package.scala 93:22:@14861.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_87 ( // @[package.scala 93:22:@14869.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_88 ( // @[package.scala 93:22:@14909.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_89 ( // @[package.scala 93:22:@14917.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_90 ( // @[package.scala 93:22:@14925.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_91 ( // @[package.scala 93:22:@14933.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_92 ( // @[package.scala 93:22:@14941.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_93 ( // @[package.scala 93:22:@14949.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_94 ( // @[package.scala 93:22:@14957.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_95 ( // @[package.scala 93:22:@14965.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  assign _T_444 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@12644.4]
  assign _T_446 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@12645.4]
  assign _T_447 = _T_444 & _T_446; // @[MemPrimitives.scala 82:228:@12646.4]
  assign _T_448 = io_wPort_0_en_0 & _T_447; // @[MemPrimitives.scala 83:102:@12647.4]
  assign _T_450 = {_T_448,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12649.4]
  assign _T_455 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@12656.4]
  assign _T_457 = io_wPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@12657.4]
  assign _T_458 = _T_455 & _T_457; // @[MemPrimitives.scala 82:228:@12658.4]
  assign _T_459 = io_wPort_1_en_0 & _T_458; // @[MemPrimitives.scala 83:102:@12659.4]
  assign _T_461 = {_T_459,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@12661.4]
  assign _T_468 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@12669.4]
  assign _T_469 = _T_444 & _T_468; // @[MemPrimitives.scala 82:228:@12670.4]
  assign _T_470 = io_wPort_0_en_0 & _T_469; // @[MemPrimitives.scala 83:102:@12671.4]
  assign _T_472 = {_T_470,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12673.4]
  assign _T_479 = io_wPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@12681.4]
  assign _T_480 = _T_455 & _T_479; // @[MemPrimitives.scala 82:228:@12682.4]
  assign _T_481 = io_wPort_1_en_0 & _T_480; // @[MemPrimitives.scala 83:102:@12683.4]
  assign _T_483 = {_T_481,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@12685.4]
  assign _T_488 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@12692.4]
  assign _T_491 = _T_488 & _T_446; // @[MemPrimitives.scala 82:228:@12694.4]
  assign _T_492 = io_wPort_0_en_0 & _T_491; // @[MemPrimitives.scala 83:102:@12695.4]
  assign _T_494 = {_T_492,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12697.4]
  assign _T_499 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@12704.4]
  assign _T_502 = _T_499 & _T_457; // @[MemPrimitives.scala 82:228:@12706.4]
  assign _T_503 = io_wPort_1_en_0 & _T_502; // @[MemPrimitives.scala 83:102:@12707.4]
  assign _T_505 = {_T_503,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@12709.4]
  assign _T_513 = _T_488 & _T_468; // @[MemPrimitives.scala 82:228:@12718.4]
  assign _T_514 = io_wPort_0_en_0 & _T_513; // @[MemPrimitives.scala 83:102:@12719.4]
  assign _T_516 = {_T_514,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12721.4]
  assign _T_524 = _T_499 & _T_479; // @[MemPrimitives.scala 82:228:@12730.4]
  assign _T_525 = io_wPort_1_en_0 & _T_524; // @[MemPrimitives.scala 83:102:@12731.4]
  assign _T_527 = {_T_525,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@12733.4]
  assign _T_532 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@12740.4]
  assign _T_535 = _T_532 & _T_446; // @[MemPrimitives.scala 82:228:@12742.4]
  assign _T_536 = io_wPort_0_en_0 & _T_535; // @[MemPrimitives.scala 83:102:@12743.4]
  assign _T_538 = {_T_536,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12745.4]
  assign _T_543 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@12752.4]
  assign _T_546 = _T_543 & _T_457; // @[MemPrimitives.scala 82:228:@12754.4]
  assign _T_547 = io_wPort_1_en_0 & _T_546; // @[MemPrimitives.scala 83:102:@12755.4]
  assign _T_549 = {_T_547,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@12757.4]
  assign _T_557 = _T_532 & _T_468; // @[MemPrimitives.scala 82:228:@12766.4]
  assign _T_558 = io_wPort_0_en_0 & _T_557; // @[MemPrimitives.scala 83:102:@12767.4]
  assign _T_560 = {_T_558,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12769.4]
  assign _T_568 = _T_543 & _T_479; // @[MemPrimitives.scala 82:228:@12778.4]
  assign _T_569 = io_wPort_1_en_0 & _T_568; // @[MemPrimitives.scala 83:102:@12779.4]
  assign _T_571 = {_T_569,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@12781.4]
  assign _T_576 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@12788.4]
  assign _T_579 = _T_576 & _T_446; // @[MemPrimitives.scala 82:228:@12790.4]
  assign _T_580 = io_wPort_0_en_0 & _T_579; // @[MemPrimitives.scala 83:102:@12791.4]
  assign _T_582 = {_T_580,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12793.4]
  assign _T_587 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@12800.4]
  assign _T_590 = _T_587 & _T_457; // @[MemPrimitives.scala 82:228:@12802.4]
  assign _T_591 = io_wPort_1_en_0 & _T_590; // @[MemPrimitives.scala 83:102:@12803.4]
  assign _T_593 = {_T_591,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@12805.4]
  assign _T_601 = _T_576 & _T_468; // @[MemPrimitives.scala 82:228:@12814.4]
  assign _T_602 = io_wPort_0_en_0 & _T_601; // @[MemPrimitives.scala 83:102:@12815.4]
  assign _T_604 = {_T_602,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@12817.4]
  assign _T_612 = _T_587 & _T_479; // @[MemPrimitives.scala 82:228:@12826.4]
  assign _T_613 = io_wPort_1_en_0 & _T_612; // @[MemPrimitives.scala 83:102:@12827.4]
  assign _T_615 = {_T_613,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@12829.4]
  assign _T_620 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12836.4]
  assign _T_622 = io_rPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@12837.4]
  assign _T_623 = _T_620 & _T_622; // @[MemPrimitives.scala 110:228:@12838.4]
  assign _T_626 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12840.4]
  assign _T_628 = io_rPort_3_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@12841.4]
  assign _T_629 = _T_626 & _T_628; // @[MemPrimitives.scala 110:228:@12842.4]
  assign _T_632 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12844.4]
  assign _T_634 = io_rPort_4_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@12845.4]
  assign _T_635 = _T_632 & _T_634; // @[MemPrimitives.scala 110:228:@12846.4]
  assign _T_638 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12848.4]
  assign _T_640 = io_rPort_6_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@12849.4]
  assign _T_641 = _T_638 & _T_640; // @[MemPrimitives.scala 110:228:@12850.4]
  assign _T_644 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12852.4]
  assign _T_646 = io_rPort_9_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@12853.4]
  assign _T_647 = _T_644 & _T_646; // @[MemPrimitives.scala 110:228:@12854.4]
  assign _T_650 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12856.4]
  assign _T_652 = io_rPort_10_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@12857.4]
  assign _T_653 = _T_650 & _T_652; // @[MemPrimitives.scala 110:228:@12858.4]
  assign _T_655 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@12869.4]
  assign _T_656 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@12870.4]
  assign _T_657 = StickySelects_io_outs_2; // @[MemPrimitives.scala 126:35:@12871.4]
  assign _T_658 = StickySelects_io_outs_3; // @[MemPrimitives.scala 126:35:@12872.4]
  assign _T_659 = StickySelects_io_outs_4; // @[MemPrimitives.scala 126:35:@12873.4]
  assign _T_660 = StickySelects_io_outs_5; // @[MemPrimitives.scala 126:35:@12874.4]
  assign _T_662 = {_T_655,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@12876.4]
  assign _T_664 = {_T_656,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@12878.4]
  assign _T_666 = {_T_657,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@12880.4]
  assign _T_668 = {_T_658,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@12882.4]
  assign _T_670 = {_T_659,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@12884.4]
  assign _T_672 = {_T_660,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@12886.4]
  assign _T_673 = _T_659 ? _T_670 : _T_672; // @[Mux.scala 31:69:@12887.4]
  assign _T_674 = _T_658 ? _T_668 : _T_673; // @[Mux.scala 31:69:@12888.4]
  assign _T_675 = _T_657 ? _T_666 : _T_674; // @[Mux.scala 31:69:@12889.4]
  assign _T_676 = _T_656 ? _T_664 : _T_675; // @[Mux.scala 31:69:@12890.4]
  assign _T_677 = _T_655 ? _T_662 : _T_676; // @[Mux.scala 31:69:@12891.4]
  assign _T_682 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12898.4]
  assign _T_684 = io_rPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@12899.4]
  assign _T_685 = _T_682 & _T_684; // @[MemPrimitives.scala 110:228:@12900.4]
  assign _T_688 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12902.4]
  assign _T_690 = io_rPort_2_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@12903.4]
  assign _T_691 = _T_688 & _T_690; // @[MemPrimitives.scala 110:228:@12904.4]
  assign _T_694 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12906.4]
  assign _T_696 = io_rPort_5_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@12907.4]
  assign _T_697 = _T_694 & _T_696; // @[MemPrimitives.scala 110:228:@12908.4]
  assign _T_700 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12910.4]
  assign _T_702 = io_rPort_7_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@12911.4]
  assign _T_703 = _T_700 & _T_702; // @[MemPrimitives.scala 110:228:@12912.4]
  assign _T_706 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12914.4]
  assign _T_708 = io_rPort_8_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@12915.4]
  assign _T_709 = _T_706 & _T_708; // @[MemPrimitives.scala 110:228:@12916.4]
  assign _T_712 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@12918.4]
  assign _T_714 = io_rPort_11_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@12919.4]
  assign _T_715 = _T_712 & _T_714; // @[MemPrimitives.scala 110:228:@12920.4]
  assign _T_717 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 126:35:@12931.4]
  assign _T_718 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 126:35:@12932.4]
  assign _T_719 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 126:35:@12933.4]
  assign _T_720 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 126:35:@12934.4]
  assign _T_721 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 126:35:@12935.4]
  assign _T_722 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 126:35:@12936.4]
  assign _T_724 = {_T_717,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@12938.4]
  assign _T_726 = {_T_718,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@12940.4]
  assign _T_728 = {_T_719,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@12942.4]
  assign _T_730 = {_T_720,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@12944.4]
  assign _T_732 = {_T_721,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@12946.4]
  assign _T_734 = {_T_722,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@12948.4]
  assign _T_735 = _T_721 ? _T_732 : _T_734; // @[Mux.scala 31:69:@12949.4]
  assign _T_736 = _T_720 ? _T_730 : _T_735; // @[Mux.scala 31:69:@12950.4]
  assign _T_737 = _T_719 ? _T_728 : _T_736; // @[Mux.scala 31:69:@12951.4]
  assign _T_738 = _T_718 ? _T_726 : _T_737; // @[Mux.scala 31:69:@12952.4]
  assign _T_739 = _T_717 ? _T_724 : _T_738; // @[Mux.scala 31:69:@12953.4]
  assign _T_746 = io_rPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12961.4]
  assign _T_747 = _T_620 & _T_746; // @[MemPrimitives.scala 110:228:@12962.4]
  assign _T_752 = io_rPort_3_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12965.4]
  assign _T_753 = _T_626 & _T_752; // @[MemPrimitives.scala 110:228:@12966.4]
  assign _T_758 = io_rPort_4_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12969.4]
  assign _T_759 = _T_632 & _T_758; // @[MemPrimitives.scala 110:228:@12970.4]
  assign _T_764 = io_rPort_6_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12973.4]
  assign _T_765 = _T_638 & _T_764; // @[MemPrimitives.scala 110:228:@12974.4]
  assign _T_770 = io_rPort_9_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12977.4]
  assign _T_771 = _T_644 & _T_770; // @[MemPrimitives.scala 110:228:@12978.4]
  assign _T_776 = io_rPort_10_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@12981.4]
  assign _T_777 = _T_650 & _T_776; // @[MemPrimitives.scala 110:228:@12982.4]
  assign _T_779 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 126:35:@12993.4]
  assign _T_780 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 126:35:@12994.4]
  assign _T_781 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 126:35:@12995.4]
  assign _T_782 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 126:35:@12996.4]
  assign _T_783 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 126:35:@12997.4]
  assign _T_784 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 126:35:@12998.4]
  assign _T_786 = {_T_779,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13000.4]
  assign _T_788 = {_T_780,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13002.4]
  assign _T_790 = {_T_781,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13004.4]
  assign _T_792 = {_T_782,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13006.4]
  assign _T_794 = {_T_783,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13008.4]
  assign _T_796 = {_T_784,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13010.4]
  assign _T_797 = _T_783 ? _T_794 : _T_796; // @[Mux.scala 31:69:@13011.4]
  assign _T_798 = _T_782 ? _T_792 : _T_797; // @[Mux.scala 31:69:@13012.4]
  assign _T_799 = _T_781 ? _T_790 : _T_798; // @[Mux.scala 31:69:@13013.4]
  assign _T_800 = _T_780 ? _T_788 : _T_799; // @[Mux.scala 31:69:@13014.4]
  assign _T_801 = _T_779 ? _T_786 : _T_800; // @[Mux.scala 31:69:@13015.4]
  assign _T_808 = io_rPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13023.4]
  assign _T_809 = _T_682 & _T_808; // @[MemPrimitives.scala 110:228:@13024.4]
  assign _T_814 = io_rPort_2_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13027.4]
  assign _T_815 = _T_688 & _T_814; // @[MemPrimitives.scala 110:228:@13028.4]
  assign _T_820 = io_rPort_5_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13031.4]
  assign _T_821 = _T_694 & _T_820; // @[MemPrimitives.scala 110:228:@13032.4]
  assign _T_826 = io_rPort_7_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13035.4]
  assign _T_827 = _T_700 & _T_826; // @[MemPrimitives.scala 110:228:@13036.4]
  assign _T_832 = io_rPort_8_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13039.4]
  assign _T_833 = _T_706 & _T_832; // @[MemPrimitives.scala 110:228:@13040.4]
  assign _T_838 = io_rPort_11_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13043.4]
  assign _T_839 = _T_712 & _T_838; // @[MemPrimitives.scala 110:228:@13044.4]
  assign _T_841 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 126:35:@13055.4]
  assign _T_842 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 126:35:@13056.4]
  assign _T_843 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 126:35:@13057.4]
  assign _T_844 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 126:35:@13058.4]
  assign _T_845 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 126:35:@13059.4]
  assign _T_846 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 126:35:@13060.4]
  assign _T_848 = {_T_841,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13062.4]
  assign _T_850 = {_T_842,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13064.4]
  assign _T_852 = {_T_843,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13066.4]
  assign _T_854 = {_T_844,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13068.4]
  assign _T_856 = {_T_845,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13070.4]
  assign _T_858 = {_T_846,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13072.4]
  assign _T_859 = _T_845 ? _T_856 : _T_858; // @[Mux.scala 31:69:@13073.4]
  assign _T_860 = _T_844 ? _T_854 : _T_859; // @[Mux.scala 31:69:@13074.4]
  assign _T_861 = _T_843 ? _T_852 : _T_860; // @[Mux.scala 31:69:@13075.4]
  assign _T_862 = _T_842 ? _T_850 : _T_861; // @[Mux.scala 31:69:@13076.4]
  assign _T_863 = _T_841 ? _T_848 : _T_862; // @[Mux.scala 31:69:@13077.4]
  assign _T_868 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13084.4]
  assign _T_871 = _T_868 & _T_622; // @[MemPrimitives.scala 110:228:@13086.4]
  assign _T_874 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13088.4]
  assign _T_877 = _T_874 & _T_628; // @[MemPrimitives.scala 110:228:@13090.4]
  assign _T_880 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13092.4]
  assign _T_883 = _T_880 & _T_634; // @[MemPrimitives.scala 110:228:@13094.4]
  assign _T_886 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13096.4]
  assign _T_889 = _T_886 & _T_640; // @[MemPrimitives.scala 110:228:@13098.4]
  assign _T_892 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13100.4]
  assign _T_895 = _T_892 & _T_646; // @[MemPrimitives.scala 110:228:@13102.4]
  assign _T_898 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13104.4]
  assign _T_901 = _T_898 & _T_652; // @[MemPrimitives.scala 110:228:@13106.4]
  assign _T_903 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 126:35:@13117.4]
  assign _T_904 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 126:35:@13118.4]
  assign _T_905 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 126:35:@13119.4]
  assign _T_906 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 126:35:@13120.4]
  assign _T_907 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 126:35:@13121.4]
  assign _T_908 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 126:35:@13122.4]
  assign _T_910 = {_T_903,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13124.4]
  assign _T_912 = {_T_904,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13126.4]
  assign _T_914 = {_T_905,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13128.4]
  assign _T_916 = {_T_906,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13130.4]
  assign _T_918 = {_T_907,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13132.4]
  assign _T_920 = {_T_908,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13134.4]
  assign _T_921 = _T_907 ? _T_918 : _T_920; // @[Mux.scala 31:69:@13135.4]
  assign _T_922 = _T_906 ? _T_916 : _T_921; // @[Mux.scala 31:69:@13136.4]
  assign _T_923 = _T_905 ? _T_914 : _T_922; // @[Mux.scala 31:69:@13137.4]
  assign _T_924 = _T_904 ? _T_912 : _T_923; // @[Mux.scala 31:69:@13138.4]
  assign _T_925 = _T_903 ? _T_910 : _T_924; // @[Mux.scala 31:69:@13139.4]
  assign _T_930 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13146.4]
  assign _T_933 = _T_930 & _T_684; // @[MemPrimitives.scala 110:228:@13148.4]
  assign _T_936 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13150.4]
  assign _T_939 = _T_936 & _T_690; // @[MemPrimitives.scala 110:228:@13152.4]
  assign _T_942 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13154.4]
  assign _T_945 = _T_942 & _T_696; // @[MemPrimitives.scala 110:228:@13156.4]
  assign _T_948 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13158.4]
  assign _T_951 = _T_948 & _T_702; // @[MemPrimitives.scala 110:228:@13160.4]
  assign _T_954 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13162.4]
  assign _T_957 = _T_954 & _T_708; // @[MemPrimitives.scala 110:228:@13164.4]
  assign _T_960 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13166.4]
  assign _T_963 = _T_960 & _T_714; // @[MemPrimitives.scala 110:228:@13168.4]
  assign _T_965 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 126:35:@13179.4]
  assign _T_966 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 126:35:@13180.4]
  assign _T_967 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 126:35:@13181.4]
  assign _T_968 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 126:35:@13182.4]
  assign _T_969 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 126:35:@13183.4]
  assign _T_970 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 126:35:@13184.4]
  assign _T_972 = {_T_965,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13186.4]
  assign _T_974 = {_T_966,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13188.4]
  assign _T_976 = {_T_967,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13190.4]
  assign _T_978 = {_T_968,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13192.4]
  assign _T_980 = {_T_969,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13194.4]
  assign _T_982 = {_T_970,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13196.4]
  assign _T_983 = _T_969 ? _T_980 : _T_982; // @[Mux.scala 31:69:@13197.4]
  assign _T_984 = _T_968 ? _T_978 : _T_983; // @[Mux.scala 31:69:@13198.4]
  assign _T_985 = _T_967 ? _T_976 : _T_984; // @[Mux.scala 31:69:@13199.4]
  assign _T_986 = _T_966 ? _T_974 : _T_985; // @[Mux.scala 31:69:@13200.4]
  assign _T_987 = _T_965 ? _T_972 : _T_986; // @[Mux.scala 31:69:@13201.4]
  assign _T_995 = _T_868 & _T_746; // @[MemPrimitives.scala 110:228:@13210.4]
  assign _T_1001 = _T_874 & _T_752; // @[MemPrimitives.scala 110:228:@13214.4]
  assign _T_1007 = _T_880 & _T_758; // @[MemPrimitives.scala 110:228:@13218.4]
  assign _T_1013 = _T_886 & _T_764; // @[MemPrimitives.scala 110:228:@13222.4]
  assign _T_1019 = _T_892 & _T_770; // @[MemPrimitives.scala 110:228:@13226.4]
  assign _T_1025 = _T_898 & _T_776; // @[MemPrimitives.scala 110:228:@13230.4]
  assign _T_1027 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 126:35:@13241.4]
  assign _T_1028 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 126:35:@13242.4]
  assign _T_1029 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 126:35:@13243.4]
  assign _T_1030 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 126:35:@13244.4]
  assign _T_1031 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 126:35:@13245.4]
  assign _T_1032 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 126:35:@13246.4]
  assign _T_1034 = {_T_1027,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13248.4]
  assign _T_1036 = {_T_1028,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13250.4]
  assign _T_1038 = {_T_1029,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13252.4]
  assign _T_1040 = {_T_1030,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13254.4]
  assign _T_1042 = {_T_1031,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13256.4]
  assign _T_1044 = {_T_1032,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13258.4]
  assign _T_1045 = _T_1031 ? _T_1042 : _T_1044; // @[Mux.scala 31:69:@13259.4]
  assign _T_1046 = _T_1030 ? _T_1040 : _T_1045; // @[Mux.scala 31:69:@13260.4]
  assign _T_1047 = _T_1029 ? _T_1038 : _T_1046; // @[Mux.scala 31:69:@13261.4]
  assign _T_1048 = _T_1028 ? _T_1036 : _T_1047; // @[Mux.scala 31:69:@13262.4]
  assign _T_1049 = _T_1027 ? _T_1034 : _T_1048; // @[Mux.scala 31:69:@13263.4]
  assign _T_1057 = _T_930 & _T_808; // @[MemPrimitives.scala 110:228:@13272.4]
  assign _T_1063 = _T_936 & _T_814; // @[MemPrimitives.scala 110:228:@13276.4]
  assign _T_1069 = _T_942 & _T_820; // @[MemPrimitives.scala 110:228:@13280.4]
  assign _T_1075 = _T_948 & _T_826; // @[MemPrimitives.scala 110:228:@13284.4]
  assign _T_1081 = _T_954 & _T_832; // @[MemPrimitives.scala 110:228:@13288.4]
  assign _T_1087 = _T_960 & _T_838; // @[MemPrimitives.scala 110:228:@13292.4]
  assign _T_1089 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 126:35:@13303.4]
  assign _T_1090 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 126:35:@13304.4]
  assign _T_1091 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 126:35:@13305.4]
  assign _T_1092 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 126:35:@13306.4]
  assign _T_1093 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 126:35:@13307.4]
  assign _T_1094 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 126:35:@13308.4]
  assign _T_1096 = {_T_1089,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13310.4]
  assign _T_1098 = {_T_1090,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13312.4]
  assign _T_1100 = {_T_1091,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13314.4]
  assign _T_1102 = {_T_1092,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13316.4]
  assign _T_1104 = {_T_1093,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13318.4]
  assign _T_1106 = {_T_1094,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13320.4]
  assign _T_1107 = _T_1093 ? _T_1104 : _T_1106; // @[Mux.scala 31:69:@13321.4]
  assign _T_1108 = _T_1092 ? _T_1102 : _T_1107; // @[Mux.scala 31:69:@13322.4]
  assign _T_1109 = _T_1091 ? _T_1100 : _T_1108; // @[Mux.scala 31:69:@13323.4]
  assign _T_1110 = _T_1090 ? _T_1098 : _T_1109; // @[Mux.scala 31:69:@13324.4]
  assign _T_1111 = _T_1089 ? _T_1096 : _T_1110; // @[Mux.scala 31:69:@13325.4]
  assign _T_1116 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13332.4]
  assign _T_1119 = _T_1116 & _T_622; // @[MemPrimitives.scala 110:228:@13334.4]
  assign _T_1122 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13336.4]
  assign _T_1125 = _T_1122 & _T_628; // @[MemPrimitives.scala 110:228:@13338.4]
  assign _T_1128 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13340.4]
  assign _T_1131 = _T_1128 & _T_634; // @[MemPrimitives.scala 110:228:@13342.4]
  assign _T_1134 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13344.4]
  assign _T_1137 = _T_1134 & _T_640; // @[MemPrimitives.scala 110:228:@13346.4]
  assign _T_1140 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13348.4]
  assign _T_1143 = _T_1140 & _T_646; // @[MemPrimitives.scala 110:228:@13350.4]
  assign _T_1146 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13352.4]
  assign _T_1149 = _T_1146 & _T_652; // @[MemPrimitives.scala 110:228:@13354.4]
  assign _T_1151 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 126:35:@13365.4]
  assign _T_1152 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 126:35:@13366.4]
  assign _T_1153 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 126:35:@13367.4]
  assign _T_1154 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 126:35:@13368.4]
  assign _T_1155 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 126:35:@13369.4]
  assign _T_1156 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 126:35:@13370.4]
  assign _T_1158 = {_T_1151,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13372.4]
  assign _T_1160 = {_T_1152,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13374.4]
  assign _T_1162 = {_T_1153,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13376.4]
  assign _T_1164 = {_T_1154,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13378.4]
  assign _T_1166 = {_T_1155,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13380.4]
  assign _T_1168 = {_T_1156,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13382.4]
  assign _T_1169 = _T_1155 ? _T_1166 : _T_1168; // @[Mux.scala 31:69:@13383.4]
  assign _T_1170 = _T_1154 ? _T_1164 : _T_1169; // @[Mux.scala 31:69:@13384.4]
  assign _T_1171 = _T_1153 ? _T_1162 : _T_1170; // @[Mux.scala 31:69:@13385.4]
  assign _T_1172 = _T_1152 ? _T_1160 : _T_1171; // @[Mux.scala 31:69:@13386.4]
  assign _T_1173 = _T_1151 ? _T_1158 : _T_1172; // @[Mux.scala 31:69:@13387.4]
  assign _T_1178 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13394.4]
  assign _T_1181 = _T_1178 & _T_684; // @[MemPrimitives.scala 110:228:@13396.4]
  assign _T_1184 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13398.4]
  assign _T_1187 = _T_1184 & _T_690; // @[MemPrimitives.scala 110:228:@13400.4]
  assign _T_1190 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13402.4]
  assign _T_1193 = _T_1190 & _T_696; // @[MemPrimitives.scala 110:228:@13404.4]
  assign _T_1196 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13406.4]
  assign _T_1199 = _T_1196 & _T_702; // @[MemPrimitives.scala 110:228:@13408.4]
  assign _T_1202 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13410.4]
  assign _T_1205 = _T_1202 & _T_708; // @[MemPrimitives.scala 110:228:@13412.4]
  assign _T_1208 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13414.4]
  assign _T_1211 = _T_1208 & _T_714; // @[MemPrimitives.scala 110:228:@13416.4]
  assign _T_1213 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 126:35:@13427.4]
  assign _T_1214 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 126:35:@13428.4]
  assign _T_1215 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 126:35:@13429.4]
  assign _T_1216 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 126:35:@13430.4]
  assign _T_1217 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 126:35:@13431.4]
  assign _T_1218 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 126:35:@13432.4]
  assign _T_1220 = {_T_1213,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13434.4]
  assign _T_1222 = {_T_1214,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13436.4]
  assign _T_1224 = {_T_1215,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13438.4]
  assign _T_1226 = {_T_1216,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13440.4]
  assign _T_1228 = {_T_1217,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13442.4]
  assign _T_1230 = {_T_1218,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13444.4]
  assign _T_1231 = _T_1217 ? _T_1228 : _T_1230; // @[Mux.scala 31:69:@13445.4]
  assign _T_1232 = _T_1216 ? _T_1226 : _T_1231; // @[Mux.scala 31:69:@13446.4]
  assign _T_1233 = _T_1215 ? _T_1224 : _T_1232; // @[Mux.scala 31:69:@13447.4]
  assign _T_1234 = _T_1214 ? _T_1222 : _T_1233; // @[Mux.scala 31:69:@13448.4]
  assign _T_1235 = _T_1213 ? _T_1220 : _T_1234; // @[Mux.scala 31:69:@13449.4]
  assign _T_1243 = _T_1116 & _T_746; // @[MemPrimitives.scala 110:228:@13458.4]
  assign _T_1249 = _T_1122 & _T_752; // @[MemPrimitives.scala 110:228:@13462.4]
  assign _T_1255 = _T_1128 & _T_758; // @[MemPrimitives.scala 110:228:@13466.4]
  assign _T_1261 = _T_1134 & _T_764; // @[MemPrimitives.scala 110:228:@13470.4]
  assign _T_1267 = _T_1140 & _T_770; // @[MemPrimitives.scala 110:228:@13474.4]
  assign _T_1273 = _T_1146 & _T_776; // @[MemPrimitives.scala 110:228:@13478.4]
  assign _T_1275 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 126:35:@13489.4]
  assign _T_1276 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 126:35:@13490.4]
  assign _T_1277 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 126:35:@13491.4]
  assign _T_1278 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 126:35:@13492.4]
  assign _T_1279 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 126:35:@13493.4]
  assign _T_1280 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 126:35:@13494.4]
  assign _T_1282 = {_T_1275,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13496.4]
  assign _T_1284 = {_T_1276,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13498.4]
  assign _T_1286 = {_T_1277,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13500.4]
  assign _T_1288 = {_T_1278,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13502.4]
  assign _T_1290 = {_T_1279,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13504.4]
  assign _T_1292 = {_T_1280,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13506.4]
  assign _T_1293 = _T_1279 ? _T_1290 : _T_1292; // @[Mux.scala 31:69:@13507.4]
  assign _T_1294 = _T_1278 ? _T_1288 : _T_1293; // @[Mux.scala 31:69:@13508.4]
  assign _T_1295 = _T_1277 ? _T_1286 : _T_1294; // @[Mux.scala 31:69:@13509.4]
  assign _T_1296 = _T_1276 ? _T_1284 : _T_1295; // @[Mux.scala 31:69:@13510.4]
  assign _T_1297 = _T_1275 ? _T_1282 : _T_1296; // @[Mux.scala 31:69:@13511.4]
  assign _T_1305 = _T_1178 & _T_808; // @[MemPrimitives.scala 110:228:@13520.4]
  assign _T_1311 = _T_1184 & _T_814; // @[MemPrimitives.scala 110:228:@13524.4]
  assign _T_1317 = _T_1190 & _T_820; // @[MemPrimitives.scala 110:228:@13528.4]
  assign _T_1323 = _T_1196 & _T_826; // @[MemPrimitives.scala 110:228:@13532.4]
  assign _T_1329 = _T_1202 & _T_832; // @[MemPrimitives.scala 110:228:@13536.4]
  assign _T_1335 = _T_1208 & _T_838; // @[MemPrimitives.scala 110:228:@13540.4]
  assign _T_1337 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 126:35:@13551.4]
  assign _T_1338 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 126:35:@13552.4]
  assign _T_1339 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 126:35:@13553.4]
  assign _T_1340 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 126:35:@13554.4]
  assign _T_1341 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 126:35:@13555.4]
  assign _T_1342 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 126:35:@13556.4]
  assign _T_1344 = {_T_1337,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13558.4]
  assign _T_1346 = {_T_1338,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13560.4]
  assign _T_1348 = {_T_1339,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13562.4]
  assign _T_1350 = {_T_1340,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13564.4]
  assign _T_1352 = {_T_1341,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13566.4]
  assign _T_1354 = {_T_1342,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13568.4]
  assign _T_1355 = _T_1341 ? _T_1352 : _T_1354; // @[Mux.scala 31:69:@13569.4]
  assign _T_1356 = _T_1340 ? _T_1350 : _T_1355; // @[Mux.scala 31:69:@13570.4]
  assign _T_1357 = _T_1339 ? _T_1348 : _T_1356; // @[Mux.scala 31:69:@13571.4]
  assign _T_1358 = _T_1338 ? _T_1346 : _T_1357; // @[Mux.scala 31:69:@13572.4]
  assign _T_1359 = _T_1337 ? _T_1344 : _T_1358; // @[Mux.scala 31:69:@13573.4]
  assign _T_1364 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13580.4]
  assign _T_1367 = _T_1364 & _T_622; // @[MemPrimitives.scala 110:228:@13582.4]
  assign _T_1370 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13584.4]
  assign _T_1373 = _T_1370 & _T_628; // @[MemPrimitives.scala 110:228:@13586.4]
  assign _T_1376 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13588.4]
  assign _T_1379 = _T_1376 & _T_634; // @[MemPrimitives.scala 110:228:@13590.4]
  assign _T_1382 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13592.4]
  assign _T_1385 = _T_1382 & _T_640; // @[MemPrimitives.scala 110:228:@13594.4]
  assign _T_1388 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13596.4]
  assign _T_1391 = _T_1388 & _T_646; // @[MemPrimitives.scala 110:228:@13598.4]
  assign _T_1394 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13600.4]
  assign _T_1397 = _T_1394 & _T_652; // @[MemPrimitives.scala 110:228:@13602.4]
  assign _T_1399 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 126:35:@13613.4]
  assign _T_1400 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 126:35:@13614.4]
  assign _T_1401 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 126:35:@13615.4]
  assign _T_1402 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 126:35:@13616.4]
  assign _T_1403 = StickySelects_12_io_outs_4; // @[MemPrimitives.scala 126:35:@13617.4]
  assign _T_1404 = StickySelects_12_io_outs_5; // @[MemPrimitives.scala 126:35:@13618.4]
  assign _T_1406 = {_T_1399,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13620.4]
  assign _T_1408 = {_T_1400,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13622.4]
  assign _T_1410 = {_T_1401,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13624.4]
  assign _T_1412 = {_T_1402,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13626.4]
  assign _T_1414 = {_T_1403,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13628.4]
  assign _T_1416 = {_T_1404,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13630.4]
  assign _T_1417 = _T_1403 ? _T_1414 : _T_1416; // @[Mux.scala 31:69:@13631.4]
  assign _T_1418 = _T_1402 ? _T_1412 : _T_1417; // @[Mux.scala 31:69:@13632.4]
  assign _T_1419 = _T_1401 ? _T_1410 : _T_1418; // @[Mux.scala 31:69:@13633.4]
  assign _T_1420 = _T_1400 ? _T_1408 : _T_1419; // @[Mux.scala 31:69:@13634.4]
  assign _T_1421 = _T_1399 ? _T_1406 : _T_1420; // @[Mux.scala 31:69:@13635.4]
  assign _T_1426 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13642.4]
  assign _T_1429 = _T_1426 & _T_684; // @[MemPrimitives.scala 110:228:@13644.4]
  assign _T_1432 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13646.4]
  assign _T_1435 = _T_1432 & _T_690; // @[MemPrimitives.scala 110:228:@13648.4]
  assign _T_1438 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13650.4]
  assign _T_1441 = _T_1438 & _T_696; // @[MemPrimitives.scala 110:228:@13652.4]
  assign _T_1444 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13654.4]
  assign _T_1447 = _T_1444 & _T_702; // @[MemPrimitives.scala 110:228:@13656.4]
  assign _T_1450 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13658.4]
  assign _T_1453 = _T_1450 & _T_708; // @[MemPrimitives.scala 110:228:@13660.4]
  assign _T_1456 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13662.4]
  assign _T_1459 = _T_1456 & _T_714; // @[MemPrimitives.scala 110:228:@13664.4]
  assign _T_1461 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 126:35:@13675.4]
  assign _T_1462 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 126:35:@13676.4]
  assign _T_1463 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 126:35:@13677.4]
  assign _T_1464 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 126:35:@13678.4]
  assign _T_1465 = StickySelects_13_io_outs_4; // @[MemPrimitives.scala 126:35:@13679.4]
  assign _T_1466 = StickySelects_13_io_outs_5; // @[MemPrimitives.scala 126:35:@13680.4]
  assign _T_1468 = {_T_1461,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13682.4]
  assign _T_1470 = {_T_1462,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13684.4]
  assign _T_1472 = {_T_1463,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13686.4]
  assign _T_1474 = {_T_1464,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13688.4]
  assign _T_1476 = {_T_1465,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13690.4]
  assign _T_1478 = {_T_1466,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13692.4]
  assign _T_1479 = _T_1465 ? _T_1476 : _T_1478; // @[Mux.scala 31:69:@13693.4]
  assign _T_1480 = _T_1464 ? _T_1474 : _T_1479; // @[Mux.scala 31:69:@13694.4]
  assign _T_1481 = _T_1463 ? _T_1472 : _T_1480; // @[Mux.scala 31:69:@13695.4]
  assign _T_1482 = _T_1462 ? _T_1470 : _T_1481; // @[Mux.scala 31:69:@13696.4]
  assign _T_1483 = _T_1461 ? _T_1468 : _T_1482; // @[Mux.scala 31:69:@13697.4]
  assign _T_1491 = _T_1364 & _T_746; // @[MemPrimitives.scala 110:228:@13706.4]
  assign _T_1497 = _T_1370 & _T_752; // @[MemPrimitives.scala 110:228:@13710.4]
  assign _T_1503 = _T_1376 & _T_758; // @[MemPrimitives.scala 110:228:@13714.4]
  assign _T_1509 = _T_1382 & _T_764; // @[MemPrimitives.scala 110:228:@13718.4]
  assign _T_1515 = _T_1388 & _T_770; // @[MemPrimitives.scala 110:228:@13722.4]
  assign _T_1521 = _T_1394 & _T_776; // @[MemPrimitives.scala 110:228:@13726.4]
  assign _T_1523 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 126:35:@13737.4]
  assign _T_1524 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 126:35:@13738.4]
  assign _T_1525 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 126:35:@13739.4]
  assign _T_1526 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 126:35:@13740.4]
  assign _T_1527 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 126:35:@13741.4]
  assign _T_1528 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 126:35:@13742.4]
  assign _T_1530 = {_T_1523,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13744.4]
  assign _T_1532 = {_T_1524,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13746.4]
  assign _T_1534 = {_T_1525,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13748.4]
  assign _T_1536 = {_T_1526,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13750.4]
  assign _T_1538 = {_T_1527,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13752.4]
  assign _T_1540 = {_T_1528,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13754.4]
  assign _T_1541 = _T_1527 ? _T_1538 : _T_1540; // @[Mux.scala 31:69:@13755.4]
  assign _T_1542 = _T_1526 ? _T_1536 : _T_1541; // @[Mux.scala 31:69:@13756.4]
  assign _T_1543 = _T_1525 ? _T_1534 : _T_1542; // @[Mux.scala 31:69:@13757.4]
  assign _T_1544 = _T_1524 ? _T_1532 : _T_1543; // @[Mux.scala 31:69:@13758.4]
  assign _T_1545 = _T_1523 ? _T_1530 : _T_1544; // @[Mux.scala 31:69:@13759.4]
  assign _T_1553 = _T_1426 & _T_808; // @[MemPrimitives.scala 110:228:@13768.4]
  assign _T_1559 = _T_1432 & _T_814; // @[MemPrimitives.scala 110:228:@13772.4]
  assign _T_1565 = _T_1438 & _T_820; // @[MemPrimitives.scala 110:228:@13776.4]
  assign _T_1571 = _T_1444 & _T_826; // @[MemPrimitives.scala 110:228:@13780.4]
  assign _T_1577 = _T_1450 & _T_832; // @[MemPrimitives.scala 110:228:@13784.4]
  assign _T_1583 = _T_1456 & _T_838; // @[MemPrimitives.scala 110:228:@13788.4]
  assign _T_1585 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 126:35:@13799.4]
  assign _T_1586 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 126:35:@13800.4]
  assign _T_1587 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 126:35:@13801.4]
  assign _T_1588 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 126:35:@13802.4]
  assign _T_1589 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 126:35:@13803.4]
  assign _T_1590 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 126:35:@13804.4]
  assign _T_1592 = {_T_1585,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13806.4]
  assign _T_1594 = {_T_1586,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13808.4]
  assign _T_1596 = {_T_1587,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13810.4]
  assign _T_1598 = {_T_1588,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13812.4]
  assign _T_1600 = {_T_1589,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13814.4]
  assign _T_1602 = {_T_1590,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13816.4]
  assign _T_1603 = _T_1589 ? _T_1600 : _T_1602; // @[Mux.scala 31:69:@13817.4]
  assign _T_1604 = _T_1588 ? _T_1598 : _T_1603; // @[Mux.scala 31:69:@13818.4]
  assign _T_1605 = _T_1587 ? _T_1596 : _T_1604; // @[Mux.scala 31:69:@13819.4]
  assign _T_1606 = _T_1586 ? _T_1594 : _T_1605; // @[Mux.scala 31:69:@13820.4]
  assign _T_1607 = _T_1585 ? _T_1592 : _T_1606; // @[Mux.scala 31:69:@13821.4]
  assign _T_1671 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@13906.4 package.scala 96:25:@13907.4]
  assign _T_1675 = _T_1671 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@13916.4]
  assign _T_1668 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@13898.4 package.scala 96:25:@13899.4]
  assign _T_1676 = _T_1668 ? Mem1D_10_io_output : _T_1675; // @[Mux.scala 31:69:@13917.4]
  assign _T_1665 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@13890.4 package.scala 96:25:@13891.4]
  assign _T_1677 = _T_1665 ? Mem1D_8_io_output : _T_1676; // @[Mux.scala 31:69:@13918.4]
  assign _T_1662 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@13882.4 package.scala 96:25:@13883.4]
  assign _T_1678 = _T_1662 ? Mem1D_6_io_output : _T_1677; // @[Mux.scala 31:69:@13919.4]
  assign _T_1659 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@13874.4 package.scala 96:25:@13875.4]
  assign _T_1679 = _T_1659 ? Mem1D_4_io_output : _T_1678; // @[Mux.scala 31:69:@13920.4]
  assign _T_1656 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@13866.4 package.scala 96:25:@13867.4]
  assign _T_1680 = _T_1656 ? Mem1D_2_io_output : _T_1679; // @[Mux.scala 31:69:@13921.4]
  assign _T_1653 = RetimeWrapper_io_out; // @[package.scala 96:25:@13858.4 package.scala 96:25:@13859.4]
  assign _T_1742 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@14002.4 package.scala 96:25:@14003.4]
  assign _T_1746 = _T_1742 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14012.4]
  assign _T_1739 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@13994.4 package.scala 96:25:@13995.4]
  assign _T_1747 = _T_1739 ? Mem1D_11_io_output : _T_1746; // @[Mux.scala 31:69:@14013.4]
  assign _T_1736 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@13986.4 package.scala 96:25:@13987.4]
  assign _T_1748 = _T_1736 ? Mem1D_9_io_output : _T_1747; // @[Mux.scala 31:69:@14014.4]
  assign _T_1733 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@13978.4 package.scala 96:25:@13979.4]
  assign _T_1749 = _T_1733 ? Mem1D_7_io_output : _T_1748; // @[Mux.scala 31:69:@14015.4]
  assign _T_1730 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@13970.4 package.scala 96:25:@13971.4]
  assign _T_1750 = _T_1730 ? Mem1D_5_io_output : _T_1749; // @[Mux.scala 31:69:@14016.4]
  assign _T_1727 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@13962.4 package.scala 96:25:@13963.4]
  assign _T_1751 = _T_1727 ? Mem1D_3_io_output : _T_1750; // @[Mux.scala 31:69:@14017.4]
  assign _T_1724 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@13954.4 package.scala 96:25:@13955.4]
  assign _T_1813 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@14098.4 package.scala 96:25:@14099.4]
  assign _T_1817 = _T_1813 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14108.4]
  assign _T_1810 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@14090.4 package.scala 96:25:@14091.4]
  assign _T_1818 = _T_1810 ? Mem1D_11_io_output : _T_1817; // @[Mux.scala 31:69:@14109.4]
  assign _T_1807 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@14082.4 package.scala 96:25:@14083.4]
  assign _T_1819 = _T_1807 ? Mem1D_9_io_output : _T_1818; // @[Mux.scala 31:69:@14110.4]
  assign _T_1804 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@14074.4 package.scala 96:25:@14075.4]
  assign _T_1820 = _T_1804 ? Mem1D_7_io_output : _T_1819; // @[Mux.scala 31:69:@14111.4]
  assign _T_1801 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@14066.4 package.scala 96:25:@14067.4]
  assign _T_1821 = _T_1801 ? Mem1D_5_io_output : _T_1820; // @[Mux.scala 31:69:@14112.4]
  assign _T_1798 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@14058.4 package.scala 96:25:@14059.4]
  assign _T_1822 = _T_1798 ? Mem1D_3_io_output : _T_1821; // @[Mux.scala 31:69:@14113.4]
  assign _T_1795 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@14050.4 package.scala 96:25:@14051.4]
  assign _T_1884 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@14194.4 package.scala 96:25:@14195.4]
  assign _T_1888 = _T_1884 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14204.4]
  assign _T_1881 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@14186.4 package.scala 96:25:@14187.4]
  assign _T_1889 = _T_1881 ? Mem1D_10_io_output : _T_1888; // @[Mux.scala 31:69:@14205.4]
  assign _T_1878 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@14178.4 package.scala 96:25:@14179.4]
  assign _T_1890 = _T_1878 ? Mem1D_8_io_output : _T_1889; // @[Mux.scala 31:69:@14206.4]
  assign _T_1875 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@14170.4 package.scala 96:25:@14171.4]
  assign _T_1891 = _T_1875 ? Mem1D_6_io_output : _T_1890; // @[Mux.scala 31:69:@14207.4]
  assign _T_1872 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@14162.4 package.scala 96:25:@14163.4]
  assign _T_1892 = _T_1872 ? Mem1D_4_io_output : _T_1891; // @[Mux.scala 31:69:@14208.4]
  assign _T_1869 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@14154.4 package.scala 96:25:@14155.4]
  assign _T_1893 = _T_1869 ? Mem1D_2_io_output : _T_1892; // @[Mux.scala 31:69:@14209.4]
  assign _T_1866 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@14146.4 package.scala 96:25:@14147.4]
  assign _T_1955 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@14290.4 package.scala 96:25:@14291.4]
  assign _T_1959 = _T_1955 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14300.4]
  assign _T_1952 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@14282.4 package.scala 96:25:@14283.4]
  assign _T_1960 = _T_1952 ? Mem1D_10_io_output : _T_1959; // @[Mux.scala 31:69:@14301.4]
  assign _T_1949 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@14274.4 package.scala 96:25:@14275.4]
  assign _T_1961 = _T_1949 ? Mem1D_8_io_output : _T_1960; // @[Mux.scala 31:69:@14302.4]
  assign _T_1946 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@14266.4 package.scala 96:25:@14267.4]
  assign _T_1962 = _T_1946 ? Mem1D_6_io_output : _T_1961; // @[Mux.scala 31:69:@14303.4]
  assign _T_1943 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@14258.4 package.scala 96:25:@14259.4]
  assign _T_1963 = _T_1943 ? Mem1D_4_io_output : _T_1962; // @[Mux.scala 31:69:@14304.4]
  assign _T_1940 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@14250.4 package.scala 96:25:@14251.4]
  assign _T_1964 = _T_1940 ? Mem1D_2_io_output : _T_1963; // @[Mux.scala 31:69:@14305.4]
  assign _T_1937 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@14242.4 package.scala 96:25:@14243.4]
  assign _T_2026 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@14386.4 package.scala 96:25:@14387.4]
  assign _T_2030 = _T_2026 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14396.4]
  assign _T_2023 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@14378.4 package.scala 96:25:@14379.4]
  assign _T_2031 = _T_2023 ? Mem1D_11_io_output : _T_2030; // @[Mux.scala 31:69:@14397.4]
  assign _T_2020 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@14370.4 package.scala 96:25:@14371.4]
  assign _T_2032 = _T_2020 ? Mem1D_9_io_output : _T_2031; // @[Mux.scala 31:69:@14398.4]
  assign _T_2017 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@14362.4 package.scala 96:25:@14363.4]
  assign _T_2033 = _T_2017 ? Mem1D_7_io_output : _T_2032; // @[Mux.scala 31:69:@14399.4]
  assign _T_2014 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@14354.4 package.scala 96:25:@14355.4]
  assign _T_2034 = _T_2014 ? Mem1D_5_io_output : _T_2033; // @[Mux.scala 31:69:@14400.4]
  assign _T_2011 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@14346.4 package.scala 96:25:@14347.4]
  assign _T_2035 = _T_2011 ? Mem1D_3_io_output : _T_2034; // @[Mux.scala 31:69:@14401.4]
  assign _T_2008 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@14338.4 package.scala 96:25:@14339.4]
  assign _T_2097 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@14482.4 package.scala 96:25:@14483.4]
  assign _T_2101 = _T_2097 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14492.4]
  assign _T_2094 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@14474.4 package.scala 96:25:@14475.4]
  assign _T_2102 = _T_2094 ? Mem1D_10_io_output : _T_2101; // @[Mux.scala 31:69:@14493.4]
  assign _T_2091 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@14466.4 package.scala 96:25:@14467.4]
  assign _T_2103 = _T_2091 ? Mem1D_8_io_output : _T_2102; // @[Mux.scala 31:69:@14494.4]
  assign _T_2088 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@14458.4 package.scala 96:25:@14459.4]
  assign _T_2104 = _T_2088 ? Mem1D_6_io_output : _T_2103; // @[Mux.scala 31:69:@14495.4]
  assign _T_2085 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@14450.4 package.scala 96:25:@14451.4]
  assign _T_2105 = _T_2085 ? Mem1D_4_io_output : _T_2104; // @[Mux.scala 31:69:@14496.4]
  assign _T_2082 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@14442.4 package.scala 96:25:@14443.4]
  assign _T_2106 = _T_2082 ? Mem1D_2_io_output : _T_2105; // @[Mux.scala 31:69:@14497.4]
  assign _T_2079 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@14434.4 package.scala 96:25:@14435.4]
  assign _T_2168 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@14578.4 package.scala 96:25:@14579.4]
  assign _T_2172 = _T_2168 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14588.4]
  assign _T_2165 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@14570.4 package.scala 96:25:@14571.4]
  assign _T_2173 = _T_2165 ? Mem1D_11_io_output : _T_2172; // @[Mux.scala 31:69:@14589.4]
  assign _T_2162 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@14562.4 package.scala 96:25:@14563.4]
  assign _T_2174 = _T_2162 ? Mem1D_9_io_output : _T_2173; // @[Mux.scala 31:69:@14590.4]
  assign _T_2159 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@14554.4 package.scala 96:25:@14555.4]
  assign _T_2175 = _T_2159 ? Mem1D_7_io_output : _T_2174; // @[Mux.scala 31:69:@14591.4]
  assign _T_2156 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@14546.4 package.scala 96:25:@14547.4]
  assign _T_2176 = _T_2156 ? Mem1D_5_io_output : _T_2175; // @[Mux.scala 31:69:@14592.4]
  assign _T_2153 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@14538.4 package.scala 96:25:@14539.4]
  assign _T_2177 = _T_2153 ? Mem1D_3_io_output : _T_2176; // @[Mux.scala 31:69:@14593.4]
  assign _T_2150 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@14530.4 package.scala 96:25:@14531.4]
  assign _T_2239 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@14674.4 package.scala 96:25:@14675.4]
  assign _T_2243 = _T_2239 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14684.4]
  assign _T_2236 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@14666.4 package.scala 96:25:@14667.4]
  assign _T_2244 = _T_2236 ? Mem1D_11_io_output : _T_2243; // @[Mux.scala 31:69:@14685.4]
  assign _T_2233 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@14658.4 package.scala 96:25:@14659.4]
  assign _T_2245 = _T_2233 ? Mem1D_9_io_output : _T_2244; // @[Mux.scala 31:69:@14686.4]
  assign _T_2230 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@14650.4 package.scala 96:25:@14651.4]
  assign _T_2246 = _T_2230 ? Mem1D_7_io_output : _T_2245; // @[Mux.scala 31:69:@14687.4]
  assign _T_2227 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@14642.4 package.scala 96:25:@14643.4]
  assign _T_2247 = _T_2227 ? Mem1D_5_io_output : _T_2246; // @[Mux.scala 31:69:@14688.4]
  assign _T_2224 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@14634.4 package.scala 96:25:@14635.4]
  assign _T_2248 = _T_2224 ? Mem1D_3_io_output : _T_2247; // @[Mux.scala 31:69:@14689.4]
  assign _T_2221 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@14626.4 package.scala 96:25:@14627.4]
  assign _T_2310 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@14770.4 package.scala 96:25:@14771.4]
  assign _T_2314 = _T_2310 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14780.4]
  assign _T_2307 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@14762.4 package.scala 96:25:@14763.4]
  assign _T_2315 = _T_2307 ? Mem1D_10_io_output : _T_2314; // @[Mux.scala 31:69:@14781.4]
  assign _T_2304 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@14754.4 package.scala 96:25:@14755.4]
  assign _T_2316 = _T_2304 ? Mem1D_8_io_output : _T_2315; // @[Mux.scala 31:69:@14782.4]
  assign _T_2301 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@14746.4 package.scala 96:25:@14747.4]
  assign _T_2317 = _T_2301 ? Mem1D_6_io_output : _T_2316; // @[Mux.scala 31:69:@14783.4]
  assign _T_2298 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@14738.4 package.scala 96:25:@14739.4]
  assign _T_2318 = _T_2298 ? Mem1D_4_io_output : _T_2317; // @[Mux.scala 31:69:@14784.4]
  assign _T_2295 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@14730.4 package.scala 96:25:@14731.4]
  assign _T_2319 = _T_2295 ? Mem1D_2_io_output : _T_2318; // @[Mux.scala 31:69:@14785.4]
  assign _T_2292 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@14722.4 package.scala 96:25:@14723.4]
  assign _T_2381 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@14866.4 package.scala 96:25:@14867.4]
  assign _T_2385 = _T_2381 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14876.4]
  assign _T_2378 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@14858.4 package.scala 96:25:@14859.4]
  assign _T_2386 = _T_2378 ? Mem1D_10_io_output : _T_2385; // @[Mux.scala 31:69:@14877.4]
  assign _T_2375 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@14850.4 package.scala 96:25:@14851.4]
  assign _T_2387 = _T_2375 ? Mem1D_8_io_output : _T_2386; // @[Mux.scala 31:69:@14878.4]
  assign _T_2372 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@14842.4 package.scala 96:25:@14843.4]
  assign _T_2388 = _T_2372 ? Mem1D_6_io_output : _T_2387; // @[Mux.scala 31:69:@14879.4]
  assign _T_2369 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@14834.4 package.scala 96:25:@14835.4]
  assign _T_2389 = _T_2369 ? Mem1D_4_io_output : _T_2388; // @[Mux.scala 31:69:@14880.4]
  assign _T_2366 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@14826.4 package.scala 96:25:@14827.4]
  assign _T_2390 = _T_2366 ? Mem1D_2_io_output : _T_2389; // @[Mux.scala 31:69:@14881.4]
  assign _T_2363 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@14818.4 package.scala 96:25:@14819.4]
  assign _T_2452 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@14962.4 package.scala 96:25:@14963.4]
  assign _T_2456 = _T_2452 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14972.4]
  assign _T_2449 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@14954.4 package.scala 96:25:@14955.4]
  assign _T_2457 = _T_2449 ? Mem1D_11_io_output : _T_2456; // @[Mux.scala 31:69:@14973.4]
  assign _T_2446 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@14946.4 package.scala 96:25:@14947.4]
  assign _T_2458 = _T_2446 ? Mem1D_9_io_output : _T_2457; // @[Mux.scala 31:69:@14974.4]
  assign _T_2443 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@14938.4 package.scala 96:25:@14939.4]
  assign _T_2459 = _T_2443 ? Mem1D_7_io_output : _T_2458; // @[Mux.scala 31:69:@14975.4]
  assign _T_2440 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@14930.4 package.scala 96:25:@14931.4]
  assign _T_2460 = _T_2440 ? Mem1D_5_io_output : _T_2459; // @[Mux.scala 31:69:@14976.4]
  assign _T_2437 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@14922.4 package.scala 96:25:@14923.4]
  assign _T_2461 = _T_2437 ? Mem1D_3_io_output : _T_2460; // @[Mux.scala 31:69:@14977.4]
  assign _T_2434 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@14914.4 package.scala 96:25:@14915.4]
  assign io_rPort_11_output_0 = _T_2434 ? Mem1D_1_io_output : _T_2461; // @[MemPrimitives.scala 152:13:@14979.4]
  assign io_rPort_10_output_0 = _T_2363 ? Mem1D_io_output : _T_2390; // @[MemPrimitives.scala 152:13:@14883.4]
  assign io_rPort_9_output_0 = _T_2292 ? Mem1D_io_output : _T_2319; // @[MemPrimitives.scala 152:13:@14787.4]
  assign io_rPort_8_output_0 = _T_2221 ? Mem1D_1_io_output : _T_2248; // @[MemPrimitives.scala 152:13:@14691.4]
  assign io_rPort_7_output_0 = _T_2150 ? Mem1D_1_io_output : _T_2177; // @[MemPrimitives.scala 152:13:@14595.4]
  assign io_rPort_6_output_0 = _T_2079 ? Mem1D_io_output : _T_2106; // @[MemPrimitives.scala 152:13:@14499.4]
  assign io_rPort_5_output_0 = _T_2008 ? Mem1D_1_io_output : _T_2035; // @[MemPrimitives.scala 152:13:@14403.4]
  assign io_rPort_4_output_0 = _T_1937 ? Mem1D_io_output : _T_1964; // @[MemPrimitives.scala 152:13:@14307.4]
  assign io_rPort_3_output_0 = _T_1866 ? Mem1D_io_output : _T_1893; // @[MemPrimitives.scala 152:13:@14211.4]
  assign io_rPort_2_output_0 = _T_1795 ? Mem1D_1_io_output : _T_1822; // @[MemPrimitives.scala 152:13:@14115.4]
  assign io_rPort_1_output_0 = _T_1724 ? Mem1D_1_io_output : _T_1751; // @[MemPrimitives.scala 152:13:@14019.4]
  assign io_rPort_0_output_0 = _T_1653 ? Mem1D_io_output : _T_1680; // @[MemPrimitives.scala 152:13:@13923.4]
  assign Mem1D_clock = clock; // @[:@12389.4]
  assign Mem1D_reset = reset; // @[:@12390.4]
  assign Mem1D_io_r_ofs_0 = _T_677[8:0]; // @[MemPrimitives.scala 131:28:@12895.4]
  assign Mem1D_io_r_backpressure = _T_677[9]; // @[MemPrimitives.scala 132:32:@12896.4]
  assign Mem1D_io_w_ofs_0 = _T_450[8:0]; // @[MemPrimitives.scala 94:28:@12653.4]
  assign Mem1D_io_w_data_0 = _T_450[40:9]; // @[MemPrimitives.scala 95:29:@12654.4]
  assign Mem1D_io_w_en_0 = _T_450[41]; // @[MemPrimitives.scala 96:27:@12655.4]
  assign Mem1D_1_clock = clock; // @[:@12405.4]
  assign Mem1D_1_reset = reset; // @[:@12406.4]
  assign Mem1D_1_io_r_ofs_0 = _T_739[8:0]; // @[MemPrimitives.scala 131:28:@12957.4]
  assign Mem1D_1_io_r_backpressure = _T_739[9]; // @[MemPrimitives.scala 132:32:@12958.4]
  assign Mem1D_1_io_w_ofs_0 = _T_461[8:0]; // @[MemPrimitives.scala 94:28:@12665.4]
  assign Mem1D_1_io_w_data_0 = _T_461[40:9]; // @[MemPrimitives.scala 95:29:@12666.4]
  assign Mem1D_1_io_w_en_0 = _T_461[41]; // @[MemPrimitives.scala 96:27:@12667.4]
  assign Mem1D_2_clock = clock; // @[:@12421.4]
  assign Mem1D_2_reset = reset; // @[:@12422.4]
  assign Mem1D_2_io_r_ofs_0 = _T_801[8:0]; // @[MemPrimitives.scala 131:28:@13019.4]
  assign Mem1D_2_io_r_backpressure = _T_801[9]; // @[MemPrimitives.scala 132:32:@13020.4]
  assign Mem1D_2_io_w_ofs_0 = _T_472[8:0]; // @[MemPrimitives.scala 94:28:@12677.4]
  assign Mem1D_2_io_w_data_0 = _T_472[40:9]; // @[MemPrimitives.scala 95:29:@12678.4]
  assign Mem1D_2_io_w_en_0 = _T_472[41]; // @[MemPrimitives.scala 96:27:@12679.4]
  assign Mem1D_3_clock = clock; // @[:@12437.4]
  assign Mem1D_3_reset = reset; // @[:@12438.4]
  assign Mem1D_3_io_r_ofs_0 = _T_863[8:0]; // @[MemPrimitives.scala 131:28:@13081.4]
  assign Mem1D_3_io_r_backpressure = _T_863[9]; // @[MemPrimitives.scala 132:32:@13082.4]
  assign Mem1D_3_io_w_ofs_0 = _T_483[8:0]; // @[MemPrimitives.scala 94:28:@12689.4]
  assign Mem1D_3_io_w_data_0 = _T_483[40:9]; // @[MemPrimitives.scala 95:29:@12690.4]
  assign Mem1D_3_io_w_en_0 = _T_483[41]; // @[MemPrimitives.scala 96:27:@12691.4]
  assign Mem1D_4_clock = clock; // @[:@12453.4]
  assign Mem1D_4_reset = reset; // @[:@12454.4]
  assign Mem1D_4_io_r_ofs_0 = _T_925[8:0]; // @[MemPrimitives.scala 131:28:@13143.4]
  assign Mem1D_4_io_r_backpressure = _T_925[9]; // @[MemPrimitives.scala 132:32:@13144.4]
  assign Mem1D_4_io_w_ofs_0 = _T_494[8:0]; // @[MemPrimitives.scala 94:28:@12701.4]
  assign Mem1D_4_io_w_data_0 = _T_494[40:9]; // @[MemPrimitives.scala 95:29:@12702.4]
  assign Mem1D_4_io_w_en_0 = _T_494[41]; // @[MemPrimitives.scala 96:27:@12703.4]
  assign Mem1D_5_clock = clock; // @[:@12469.4]
  assign Mem1D_5_reset = reset; // @[:@12470.4]
  assign Mem1D_5_io_r_ofs_0 = _T_987[8:0]; // @[MemPrimitives.scala 131:28:@13205.4]
  assign Mem1D_5_io_r_backpressure = _T_987[9]; // @[MemPrimitives.scala 132:32:@13206.4]
  assign Mem1D_5_io_w_ofs_0 = _T_505[8:0]; // @[MemPrimitives.scala 94:28:@12713.4]
  assign Mem1D_5_io_w_data_0 = _T_505[40:9]; // @[MemPrimitives.scala 95:29:@12714.4]
  assign Mem1D_5_io_w_en_0 = _T_505[41]; // @[MemPrimitives.scala 96:27:@12715.4]
  assign Mem1D_6_clock = clock; // @[:@12485.4]
  assign Mem1D_6_reset = reset; // @[:@12486.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1049[8:0]; // @[MemPrimitives.scala 131:28:@13267.4]
  assign Mem1D_6_io_r_backpressure = _T_1049[9]; // @[MemPrimitives.scala 132:32:@13268.4]
  assign Mem1D_6_io_w_ofs_0 = _T_516[8:0]; // @[MemPrimitives.scala 94:28:@12725.4]
  assign Mem1D_6_io_w_data_0 = _T_516[40:9]; // @[MemPrimitives.scala 95:29:@12726.4]
  assign Mem1D_6_io_w_en_0 = _T_516[41]; // @[MemPrimitives.scala 96:27:@12727.4]
  assign Mem1D_7_clock = clock; // @[:@12501.4]
  assign Mem1D_7_reset = reset; // @[:@12502.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1111[8:0]; // @[MemPrimitives.scala 131:28:@13329.4]
  assign Mem1D_7_io_r_backpressure = _T_1111[9]; // @[MemPrimitives.scala 132:32:@13330.4]
  assign Mem1D_7_io_w_ofs_0 = _T_527[8:0]; // @[MemPrimitives.scala 94:28:@12737.4]
  assign Mem1D_7_io_w_data_0 = _T_527[40:9]; // @[MemPrimitives.scala 95:29:@12738.4]
  assign Mem1D_7_io_w_en_0 = _T_527[41]; // @[MemPrimitives.scala 96:27:@12739.4]
  assign Mem1D_8_clock = clock; // @[:@12517.4]
  assign Mem1D_8_reset = reset; // @[:@12518.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1173[8:0]; // @[MemPrimitives.scala 131:28:@13391.4]
  assign Mem1D_8_io_r_backpressure = _T_1173[9]; // @[MemPrimitives.scala 132:32:@13392.4]
  assign Mem1D_8_io_w_ofs_0 = _T_538[8:0]; // @[MemPrimitives.scala 94:28:@12749.4]
  assign Mem1D_8_io_w_data_0 = _T_538[40:9]; // @[MemPrimitives.scala 95:29:@12750.4]
  assign Mem1D_8_io_w_en_0 = _T_538[41]; // @[MemPrimitives.scala 96:27:@12751.4]
  assign Mem1D_9_clock = clock; // @[:@12533.4]
  assign Mem1D_9_reset = reset; // @[:@12534.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1235[8:0]; // @[MemPrimitives.scala 131:28:@13453.4]
  assign Mem1D_9_io_r_backpressure = _T_1235[9]; // @[MemPrimitives.scala 132:32:@13454.4]
  assign Mem1D_9_io_w_ofs_0 = _T_549[8:0]; // @[MemPrimitives.scala 94:28:@12761.4]
  assign Mem1D_9_io_w_data_0 = _T_549[40:9]; // @[MemPrimitives.scala 95:29:@12762.4]
  assign Mem1D_9_io_w_en_0 = _T_549[41]; // @[MemPrimitives.scala 96:27:@12763.4]
  assign Mem1D_10_clock = clock; // @[:@12549.4]
  assign Mem1D_10_reset = reset; // @[:@12550.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1297[8:0]; // @[MemPrimitives.scala 131:28:@13515.4]
  assign Mem1D_10_io_r_backpressure = _T_1297[9]; // @[MemPrimitives.scala 132:32:@13516.4]
  assign Mem1D_10_io_w_ofs_0 = _T_560[8:0]; // @[MemPrimitives.scala 94:28:@12773.4]
  assign Mem1D_10_io_w_data_0 = _T_560[40:9]; // @[MemPrimitives.scala 95:29:@12774.4]
  assign Mem1D_10_io_w_en_0 = _T_560[41]; // @[MemPrimitives.scala 96:27:@12775.4]
  assign Mem1D_11_clock = clock; // @[:@12565.4]
  assign Mem1D_11_reset = reset; // @[:@12566.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1359[8:0]; // @[MemPrimitives.scala 131:28:@13577.4]
  assign Mem1D_11_io_r_backpressure = _T_1359[9]; // @[MemPrimitives.scala 132:32:@13578.4]
  assign Mem1D_11_io_w_ofs_0 = _T_571[8:0]; // @[MemPrimitives.scala 94:28:@12785.4]
  assign Mem1D_11_io_w_data_0 = _T_571[40:9]; // @[MemPrimitives.scala 95:29:@12786.4]
  assign Mem1D_11_io_w_en_0 = _T_571[41]; // @[MemPrimitives.scala 96:27:@12787.4]
  assign Mem1D_12_clock = clock; // @[:@12581.4]
  assign Mem1D_12_reset = reset; // @[:@12582.4]
  assign Mem1D_12_io_r_ofs_0 = _T_1421[8:0]; // @[MemPrimitives.scala 131:28:@13639.4]
  assign Mem1D_12_io_r_backpressure = _T_1421[9]; // @[MemPrimitives.scala 132:32:@13640.4]
  assign Mem1D_12_io_w_ofs_0 = _T_582[8:0]; // @[MemPrimitives.scala 94:28:@12797.4]
  assign Mem1D_12_io_w_data_0 = _T_582[40:9]; // @[MemPrimitives.scala 95:29:@12798.4]
  assign Mem1D_12_io_w_en_0 = _T_582[41]; // @[MemPrimitives.scala 96:27:@12799.4]
  assign Mem1D_13_clock = clock; // @[:@12597.4]
  assign Mem1D_13_reset = reset; // @[:@12598.4]
  assign Mem1D_13_io_r_ofs_0 = _T_1483[8:0]; // @[MemPrimitives.scala 131:28:@13701.4]
  assign Mem1D_13_io_r_backpressure = _T_1483[9]; // @[MemPrimitives.scala 132:32:@13702.4]
  assign Mem1D_13_io_w_ofs_0 = _T_593[8:0]; // @[MemPrimitives.scala 94:28:@12809.4]
  assign Mem1D_13_io_w_data_0 = _T_593[40:9]; // @[MemPrimitives.scala 95:29:@12810.4]
  assign Mem1D_13_io_w_en_0 = _T_593[41]; // @[MemPrimitives.scala 96:27:@12811.4]
  assign Mem1D_14_clock = clock; // @[:@12613.4]
  assign Mem1D_14_reset = reset; // @[:@12614.4]
  assign Mem1D_14_io_r_ofs_0 = _T_1545[8:0]; // @[MemPrimitives.scala 131:28:@13763.4]
  assign Mem1D_14_io_r_backpressure = _T_1545[9]; // @[MemPrimitives.scala 132:32:@13764.4]
  assign Mem1D_14_io_w_ofs_0 = _T_604[8:0]; // @[MemPrimitives.scala 94:28:@12821.4]
  assign Mem1D_14_io_w_data_0 = _T_604[40:9]; // @[MemPrimitives.scala 95:29:@12822.4]
  assign Mem1D_14_io_w_en_0 = _T_604[41]; // @[MemPrimitives.scala 96:27:@12823.4]
  assign Mem1D_15_clock = clock; // @[:@12629.4]
  assign Mem1D_15_reset = reset; // @[:@12630.4]
  assign Mem1D_15_io_r_ofs_0 = _T_1607[8:0]; // @[MemPrimitives.scala 131:28:@13825.4]
  assign Mem1D_15_io_r_backpressure = _T_1607[9]; // @[MemPrimitives.scala 132:32:@13826.4]
  assign Mem1D_15_io_w_ofs_0 = _T_615[8:0]; // @[MemPrimitives.scala 94:28:@12833.4]
  assign Mem1D_15_io_w_data_0 = _T_615[40:9]; // @[MemPrimitives.scala 95:29:@12834.4]
  assign Mem1D_15_io_w_en_0 = _T_615[41]; // @[MemPrimitives.scala 96:27:@12835.4]
  assign StickySelects_clock = clock; // @[:@12861.4]
  assign StickySelects_reset = reset; // @[:@12862.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0 & _T_623; // @[MemPrimitives.scala 125:64:@12863.4]
  assign StickySelects_io_ins_1 = io_rPort_3_en_0 & _T_629; // @[MemPrimitives.scala 125:64:@12864.4]
  assign StickySelects_io_ins_2 = io_rPort_4_en_0 & _T_635; // @[MemPrimitives.scala 125:64:@12865.4]
  assign StickySelects_io_ins_3 = io_rPort_6_en_0 & _T_641; // @[MemPrimitives.scala 125:64:@12866.4]
  assign StickySelects_io_ins_4 = io_rPort_9_en_0 & _T_647; // @[MemPrimitives.scala 125:64:@12867.4]
  assign StickySelects_io_ins_5 = io_rPort_10_en_0 & _T_653; // @[MemPrimitives.scala 125:64:@12868.4]
  assign StickySelects_1_clock = clock; // @[:@12923.4]
  assign StickySelects_1_reset = reset; // @[:@12924.4]
  assign StickySelects_1_io_ins_0 = io_rPort_1_en_0 & _T_685; // @[MemPrimitives.scala 125:64:@12925.4]
  assign StickySelects_1_io_ins_1 = io_rPort_2_en_0 & _T_691; // @[MemPrimitives.scala 125:64:@12926.4]
  assign StickySelects_1_io_ins_2 = io_rPort_5_en_0 & _T_697; // @[MemPrimitives.scala 125:64:@12927.4]
  assign StickySelects_1_io_ins_3 = io_rPort_7_en_0 & _T_703; // @[MemPrimitives.scala 125:64:@12928.4]
  assign StickySelects_1_io_ins_4 = io_rPort_8_en_0 & _T_709; // @[MemPrimitives.scala 125:64:@12929.4]
  assign StickySelects_1_io_ins_5 = io_rPort_11_en_0 & _T_715; // @[MemPrimitives.scala 125:64:@12930.4]
  assign StickySelects_2_clock = clock; // @[:@12985.4]
  assign StickySelects_2_reset = reset; // @[:@12986.4]
  assign StickySelects_2_io_ins_0 = io_rPort_0_en_0 & _T_747; // @[MemPrimitives.scala 125:64:@12987.4]
  assign StickySelects_2_io_ins_1 = io_rPort_3_en_0 & _T_753; // @[MemPrimitives.scala 125:64:@12988.4]
  assign StickySelects_2_io_ins_2 = io_rPort_4_en_0 & _T_759; // @[MemPrimitives.scala 125:64:@12989.4]
  assign StickySelects_2_io_ins_3 = io_rPort_6_en_0 & _T_765; // @[MemPrimitives.scala 125:64:@12990.4]
  assign StickySelects_2_io_ins_4 = io_rPort_9_en_0 & _T_771; // @[MemPrimitives.scala 125:64:@12991.4]
  assign StickySelects_2_io_ins_5 = io_rPort_10_en_0 & _T_777; // @[MemPrimitives.scala 125:64:@12992.4]
  assign StickySelects_3_clock = clock; // @[:@13047.4]
  assign StickySelects_3_reset = reset; // @[:@13048.4]
  assign StickySelects_3_io_ins_0 = io_rPort_1_en_0 & _T_809; // @[MemPrimitives.scala 125:64:@13049.4]
  assign StickySelects_3_io_ins_1 = io_rPort_2_en_0 & _T_815; // @[MemPrimitives.scala 125:64:@13050.4]
  assign StickySelects_3_io_ins_2 = io_rPort_5_en_0 & _T_821; // @[MemPrimitives.scala 125:64:@13051.4]
  assign StickySelects_3_io_ins_3 = io_rPort_7_en_0 & _T_827; // @[MemPrimitives.scala 125:64:@13052.4]
  assign StickySelects_3_io_ins_4 = io_rPort_8_en_0 & _T_833; // @[MemPrimitives.scala 125:64:@13053.4]
  assign StickySelects_3_io_ins_5 = io_rPort_11_en_0 & _T_839; // @[MemPrimitives.scala 125:64:@13054.4]
  assign StickySelects_4_clock = clock; // @[:@13109.4]
  assign StickySelects_4_reset = reset; // @[:@13110.4]
  assign StickySelects_4_io_ins_0 = io_rPort_0_en_0 & _T_871; // @[MemPrimitives.scala 125:64:@13111.4]
  assign StickySelects_4_io_ins_1 = io_rPort_3_en_0 & _T_877; // @[MemPrimitives.scala 125:64:@13112.4]
  assign StickySelects_4_io_ins_2 = io_rPort_4_en_0 & _T_883; // @[MemPrimitives.scala 125:64:@13113.4]
  assign StickySelects_4_io_ins_3 = io_rPort_6_en_0 & _T_889; // @[MemPrimitives.scala 125:64:@13114.4]
  assign StickySelects_4_io_ins_4 = io_rPort_9_en_0 & _T_895; // @[MemPrimitives.scala 125:64:@13115.4]
  assign StickySelects_4_io_ins_5 = io_rPort_10_en_0 & _T_901; // @[MemPrimitives.scala 125:64:@13116.4]
  assign StickySelects_5_clock = clock; // @[:@13171.4]
  assign StickySelects_5_reset = reset; // @[:@13172.4]
  assign StickySelects_5_io_ins_0 = io_rPort_1_en_0 & _T_933; // @[MemPrimitives.scala 125:64:@13173.4]
  assign StickySelects_5_io_ins_1 = io_rPort_2_en_0 & _T_939; // @[MemPrimitives.scala 125:64:@13174.4]
  assign StickySelects_5_io_ins_2 = io_rPort_5_en_0 & _T_945; // @[MemPrimitives.scala 125:64:@13175.4]
  assign StickySelects_5_io_ins_3 = io_rPort_7_en_0 & _T_951; // @[MemPrimitives.scala 125:64:@13176.4]
  assign StickySelects_5_io_ins_4 = io_rPort_8_en_0 & _T_957; // @[MemPrimitives.scala 125:64:@13177.4]
  assign StickySelects_5_io_ins_5 = io_rPort_11_en_0 & _T_963; // @[MemPrimitives.scala 125:64:@13178.4]
  assign StickySelects_6_clock = clock; // @[:@13233.4]
  assign StickySelects_6_reset = reset; // @[:@13234.4]
  assign StickySelects_6_io_ins_0 = io_rPort_0_en_0 & _T_995; // @[MemPrimitives.scala 125:64:@13235.4]
  assign StickySelects_6_io_ins_1 = io_rPort_3_en_0 & _T_1001; // @[MemPrimitives.scala 125:64:@13236.4]
  assign StickySelects_6_io_ins_2 = io_rPort_4_en_0 & _T_1007; // @[MemPrimitives.scala 125:64:@13237.4]
  assign StickySelects_6_io_ins_3 = io_rPort_6_en_0 & _T_1013; // @[MemPrimitives.scala 125:64:@13238.4]
  assign StickySelects_6_io_ins_4 = io_rPort_9_en_0 & _T_1019; // @[MemPrimitives.scala 125:64:@13239.4]
  assign StickySelects_6_io_ins_5 = io_rPort_10_en_0 & _T_1025; // @[MemPrimitives.scala 125:64:@13240.4]
  assign StickySelects_7_clock = clock; // @[:@13295.4]
  assign StickySelects_7_reset = reset; // @[:@13296.4]
  assign StickySelects_7_io_ins_0 = io_rPort_1_en_0 & _T_1057; // @[MemPrimitives.scala 125:64:@13297.4]
  assign StickySelects_7_io_ins_1 = io_rPort_2_en_0 & _T_1063; // @[MemPrimitives.scala 125:64:@13298.4]
  assign StickySelects_7_io_ins_2 = io_rPort_5_en_0 & _T_1069; // @[MemPrimitives.scala 125:64:@13299.4]
  assign StickySelects_7_io_ins_3 = io_rPort_7_en_0 & _T_1075; // @[MemPrimitives.scala 125:64:@13300.4]
  assign StickySelects_7_io_ins_4 = io_rPort_8_en_0 & _T_1081; // @[MemPrimitives.scala 125:64:@13301.4]
  assign StickySelects_7_io_ins_5 = io_rPort_11_en_0 & _T_1087; // @[MemPrimitives.scala 125:64:@13302.4]
  assign StickySelects_8_clock = clock; // @[:@13357.4]
  assign StickySelects_8_reset = reset; // @[:@13358.4]
  assign StickySelects_8_io_ins_0 = io_rPort_0_en_0 & _T_1119; // @[MemPrimitives.scala 125:64:@13359.4]
  assign StickySelects_8_io_ins_1 = io_rPort_3_en_0 & _T_1125; // @[MemPrimitives.scala 125:64:@13360.4]
  assign StickySelects_8_io_ins_2 = io_rPort_4_en_0 & _T_1131; // @[MemPrimitives.scala 125:64:@13361.4]
  assign StickySelects_8_io_ins_3 = io_rPort_6_en_0 & _T_1137; // @[MemPrimitives.scala 125:64:@13362.4]
  assign StickySelects_8_io_ins_4 = io_rPort_9_en_0 & _T_1143; // @[MemPrimitives.scala 125:64:@13363.4]
  assign StickySelects_8_io_ins_5 = io_rPort_10_en_0 & _T_1149; // @[MemPrimitives.scala 125:64:@13364.4]
  assign StickySelects_9_clock = clock; // @[:@13419.4]
  assign StickySelects_9_reset = reset; // @[:@13420.4]
  assign StickySelects_9_io_ins_0 = io_rPort_1_en_0 & _T_1181; // @[MemPrimitives.scala 125:64:@13421.4]
  assign StickySelects_9_io_ins_1 = io_rPort_2_en_0 & _T_1187; // @[MemPrimitives.scala 125:64:@13422.4]
  assign StickySelects_9_io_ins_2 = io_rPort_5_en_0 & _T_1193; // @[MemPrimitives.scala 125:64:@13423.4]
  assign StickySelects_9_io_ins_3 = io_rPort_7_en_0 & _T_1199; // @[MemPrimitives.scala 125:64:@13424.4]
  assign StickySelects_9_io_ins_4 = io_rPort_8_en_0 & _T_1205; // @[MemPrimitives.scala 125:64:@13425.4]
  assign StickySelects_9_io_ins_5 = io_rPort_11_en_0 & _T_1211; // @[MemPrimitives.scala 125:64:@13426.4]
  assign StickySelects_10_clock = clock; // @[:@13481.4]
  assign StickySelects_10_reset = reset; // @[:@13482.4]
  assign StickySelects_10_io_ins_0 = io_rPort_0_en_0 & _T_1243; // @[MemPrimitives.scala 125:64:@13483.4]
  assign StickySelects_10_io_ins_1 = io_rPort_3_en_0 & _T_1249; // @[MemPrimitives.scala 125:64:@13484.4]
  assign StickySelects_10_io_ins_2 = io_rPort_4_en_0 & _T_1255; // @[MemPrimitives.scala 125:64:@13485.4]
  assign StickySelects_10_io_ins_3 = io_rPort_6_en_0 & _T_1261; // @[MemPrimitives.scala 125:64:@13486.4]
  assign StickySelects_10_io_ins_4 = io_rPort_9_en_0 & _T_1267; // @[MemPrimitives.scala 125:64:@13487.4]
  assign StickySelects_10_io_ins_5 = io_rPort_10_en_0 & _T_1273; // @[MemPrimitives.scala 125:64:@13488.4]
  assign StickySelects_11_clock = clock; // @[:@13543.4]
  assign StickySelects_11_reset = reset; // @[:@13544.4]
  assign StickySelects_11_io_ins_0 = io_rPort_1_en_0 & _T_1305; // @[MemPrimitives.scala 125:64:@13545.4]
  assign StickySelects_11_io_ins_1 = io_rPort_2_en_0 & _T_1311; // @[MemPrimitives.scala 125:64:@13546.4]
  assign StickySelects_11_io_ins_2 = io_rPort_5_en_0 & _T_1317; // @[MemPrimitives.scala 125:64:@13547.4]
  assign StickySelects_11_io_ins_3 = io_rPort_7_en_0 & _T_1323; // @[MemPrimitives.scala 125:64:@13548.4]
  assign StickySelects_11_io_ins_4 = io_rPort_8_en_0 & _T_1329; // @[MemPrimitives.scala 125:64:@13549.4]
  assign StickySelects_11_io_ins_5 = io_rPort_11_en_0 & _T_1335; // @[MemPrimitives.scala 125:64:@13550.4]
  assign StickySelects_12_clock = clock; // @[:@13605.4]
  assign StickySelects_12_reset = reset; // @[:@13606.4]
  assign StickySelects_12_io_ins_0 = io_rPort_0_en_0 & _T_1367; // @[MemPrimitives.scala 125:64:@13607.4]
  assign StickySelects_12_io_ins_1 = io_rPort_3_en_0 & _T_1373; // @[MemPrimitives.scala 125:64:@13608.4]
  assign StickySelects_12_io_ins_2 = io_rPort_4_en_0 & _T_1379; // @[MemPrimitives.scala 125:64:@13609.4]
  assign StickySelects_12_io_ins_3 = io_rPort_6_en_0 & _T_1385; // @[MemPrimitives.scala 125:64:@13610.4]
  assign StickySelects_12_io_ins_4 = io_rPort_9_en_0 & _T_1391; // @[MemPrimitives.scala 125:64:@13611.4]
  assign StickySelects_12_io_ins_5 = io_rPort_10_en_0 & _T_1397; // @[MemPrimitives.scala 125:64:@13612.4]
  assign StickySelects_13_clock = clock; // @[:@13667.4]
  assign StickySelects_13_reset = reset; // @[:@13668.4]
  assign StickySelects_13_io_ins_0 = io_rPort_1_en_0 & _T_1429; // @[MemPrimitives.scala 125:64:@13669.4]
  assign StickySelects_13_io_ins_1 = io_rPort_2_en_0 & _T_1435; // @[MemPrimitives.scala 125:64:@13670.4]
  assign StickySelects_13_io_ins_2 = io_rPort_5_en_0 & _T_1441; // @[MemPrimitives.scala 125:64:@13671.4]
  assign StickySelects_13_io_ins_3 = io_rPort_7_en_0 & _T_1447; // @[MemPrimitives.scala 125:64:@13672.4]
  assign StickySelects_13_io_ins_4 = io_rPort_8_en_0 & _T_1453; // @[MemPrimitives.scala 125:64:@13673.4]
  assign StickySelects_13_io_ins_5 = io_rPort_11_en_0 & _T_1459; // @[MemPrimitives.scala 125:64:@13674.4]
  assign StickySelects_14_clock = clock; // @[:@13729.4]
  assign StickySelects_14_reset = reset; // @[:@13730.4]
  assign StickySelects_14_io_ins_0 = io_rPort_0_en_0 & _T_1491; // @[MemPrimitives.scala 125:64:@13731.4]
  assign StickySelects_14_io_ins_1 = io_rPort_3_en_0 & _T_1497; // @[MemPrimitives.scala 125:64:@13732.4]
  assign StickySelects_14_io_ins_2 = io_rPort_4_en_0 & _T_1503; // @[MemPrimitives.scala 125:64:@13733.4]
  assign StickySelects_14_io_ins_3 = io_rPort_6_en_0 & _T_1509; // @[MemPrimitives.scala 125:64:@13734.4]
  assign StickySelects_14_io_ins_4 = io_rPort_9_en_0 & _T_1515; // @[MemPrimitives.scala 125:64:@13735.4]
  assign StickySelects_14_io_ins_5 = io_rPort_10_en_0 & _T_1521; // @[MemPrimitives.scala 125:64:@13736.4]
  assign StickySelects_15_clock = clock; // @[:@13791.4]
  assign StickySelects_15_reset = reset; // @[:@13792.4]
  assign StickySelects_15_io_ins_0 = io_rPort_1_en_0 & _T_1553; // @[MemPrimitives.scala 125:64:@13793.4]
  assign StickySelects_15_io_ins_1 = io_rPort_2_en_0 & _T_1559; // @[MemPrimitives.scala 125:64:@13794.4]
  assign StickySelects_15_io_ins_2 = io_rPort_5_en_0 & _T_1565; // @[MemPrimitives.scala 125:64:@13795.4]
  assign StickySelects_15_io_ins_3 = io_rPort_7_en_0 & _T_1571; // @[MemPrimitives.scala 125:64:@13796.4]
  assign StickySelects_15_io_ins_4 = io_rPort_8_en_0 & _T_1577; // @[MemPrimitives.scala 125:64:@13797.4]
  assign StickySelects_15_io_ins_5 = io_rPort_11_en_0 & _T_1583; // @[MemPrimitives.scala 125:64:@13798.4]
  assign RetimeWrapper_clock = clock; // @[:@13854.4]
  assign RetimeWrapper_reset = reset; // @[:@13855.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13857.4]
  assign RetimeWrapper_io_in = _T_623 & io_rPort_0_en_0; // @[package.scala 94:16:@13856.4]
  assign RetimeWrapper_1_clock = clock; // @[:@13862.4]
  assign RetimeWrapper_1_reset = reset; // @[:@13863.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13865.4]
  assign RetimeWrapper_1_io_in = _T_747 & io_rPort_0_en_0; // @[package.scala 94:16:@13864.4]
  assign RetimeWrapper_2_clock = clock; // @[:@13870.4]
  assign RetimeWrapper_2_reset = reset; // @[:@13871.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13873.4]
  assign RetimeWrapper_2_io_in = _T_871 & io_rPort_0_en_0; // @[package.scala 94:16:@13872.4]
  assign RetimeWrapper_3_clock = clock; // @[:@13878.4]
  assign RetimeWrapper_3_reset = reset; // @[:@13879.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13881.4]
  assign RetimeWrapper_3_io_in = _T_995 & io_rPort_0_en_0; // @[package.scala 94:16:@13880.4]
  assign RetimeWrapper_4_clock = clock; // @[:@13886.4]
  assign RetimeWrapper_4_reset = reset; // @[:@13887.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13889.4]
  assign RetimeWrapper_4_io_in = _T_1119 & io_rPort_0_en_0; // @[package.scala 94:16:@13888.4]
  assign RetimeWrapper_5_clock = clock; // @[:@13894.4]
  assign RetimeWrapper_5_reset = reset; // @[:@13895.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13897.4]
  assign RetimeWrapper_5_io_in = _T_1243 & io_rPort_0_en_0; // @[package.scala 94:16:@13896.4]
  assign RetimeWrapper_6_clock = clock; // @[:@13902.4]
  assign RetimeWrapper_6_reset = reset; // @[:@13903.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13905.4]
  assign RetimeWrapper_6_io_in = _T_1367 & io_rPort_0_en_0; // @[package.scala 94:16:@13904.4]
  assign RetimeWrapper_7_clock = clock; // @[:@13910.4]
  assign RetimeWrapper_7_reset = reset; // @[:@13911.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@13913.4]
  assign RetimeWrapper_7_io_in = _T_1491 & io_rPort_0_en_0; // @[package.scala 94:16:@13912.4]
  assign RetimeWrapper_8_clock = clock; // @[:@13950.4]
  assign RetimeWrapper_8_reset = reset; // @[:@13951.4]
  assign RetimeWrapper_8_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13953.4]
  assign RetimeWrapper_8_io_in = _T_685 & io_rPort_1_en_0; // @[package.scala 94:16:@13952.4]
  assign RetimeWrapper_9_clock = clock; // @[:@13958.4]
  assign RetimeWrapper_9_reset = reset; // @[:@13959.4]
  assign RetimeWrapper_9_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13961.4]
  assign RetimeWrapper_9_io_in = _T_809 & io_rPort_1_en_0; // @[package.scala 94:16:@13960.4]
  assign RetimeWrapper_10_clock = clock; // @[:@13966.4]
  assign RetimeWrapper_10_reset = reset; // @[:@13967.4]
  assign RetimeWrapper_10_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13969.4]
  assign RetimeWrapper_10_io_in = _T_933 & io_rPort_1_en_0; // @[package.scala 94:16:@13968.4]
  assign RetimeWrapper_11_clock = clock; // @[:@13974.4]
  assign RetimeWrapper_11_reset = reset; // @[:@13975.4]
  assign RetimeWrapper_11_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13977.4]
  assign RetimeWrapper_11_io_in = _T_1057 & io_rPort_1_en_0; // @[package.scala 94:16:@13976.4]
  assign RetimeWrapper_12_clock = clock; // @[:@13982.4]
  assign RetimeWrapper_12_reset = reset; // @[:@13983.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13985.4]
  assign RetimeWrapper_12_io_in = _T_1181 & io_rPort_1_en_0; // @[package.scala 94:16:@13984.4]
  assign RetimeWrapper_13_clock = clock; // @[:@13990.4]
  assign RetimeWrapper_13_reset = reset; // @[:@13991.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@13993.4]
  assign RetimeWrapper_13_io_in = _T_1305 & io_rPort_1_en_0; // @[package.scala 94:16:@13992.4]
  assign RetimeWrapper_14_clock = clock; // @[:@13998.4]
  assign RetimeWrapper_14_reset = reset; // @[:@13999.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14001.4]
  assign RetimeWrapper_14_io_in = _T_1429 & io_rPort_1_en_0; // @[package.scala 94:16:@14000.4]
  assign RetimeWrapper_15_clock = clock; // @[:@14006.4]
  assign RetimeWrapper_15_reset = reset; // @[:@14007.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14009.4]
  assign RetimeWrapper_15_io_in = _T_1553 & io_rPort_1_en_0; // @[package.scala 94:16:@14008.4]
  assign RetimeWrapper_16_clock = clock; // @[:@14046.4]
  assign RetimeWrapper_16_reset = reset; // @[:@14047.4]
  assign RetimeWrapper_16_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14049.4]
  assign RetimeWrapper_16_io_in = _T_691 & io_rPort_2_en_0; // @[package.scala 94:16:@14048.4]
  assign RetimeWrapper_17_clock = clock; // @[:@14054.4]
  assign RetimeWrapper_17_reset = reset; // @[:@14055.4]
  assign RetimeWrapper_17_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14057.4]
  assign RetimeWrapper_17_io_in = _T_815 & io_rPort_2_en_0; // @[package.scala 94:16:@14056.4]
  assign RetimeWrapper_18_clock = clock; // @[:@14062.4]
  assign RetimeWrapper_18_reset = reset; // @[:@14063.4]
  assign RetimeWrapper_18_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14065.4]
  assign RetimeWrapper_18_io_in = _T_939 & io_rPort_2_en_0; // @[package.scala 94:16:@14064.4]
  assign RetimeWrapper_19_clock = clock; // @[:@14070.4]
  assign RetimeWrapper_19_reset = reset; // @[:@14071.4]
  assign RetimeWrapper_19_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14073.4]
  assign RetimeWrapper_19_io_in = _T_1063 & io_rPort_2_en_0; // @[package.scala 94:16:@14072.4]
  assign RetimeWrapper_20_clock = clock; // @[:@14078.4]
  assign RetimeWrapper_20_reset = reset; // @[:@14079.4]
  assign RetimeWrapper_20_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14081.4]
  assign RetimeWrapper_20_io_in = _T_1187 & io_rPort_2_en_0; // @[package.scala 94:16:@14080.4]
  assign RetimeWrapper_21_clock = clock; // @[:@14086.4]
  assign RetimeWrapper_21_reset = reset; // @[:@14087.4]
  assign RetimeWrapper_21_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14089.4]
  assign RetimeWrapper_21_io_in = _T_1311 & io_rPort_2_en_0; // @[package.scala 94:16:@14088.4]
  assign RetimeWrapper_22_clock = clock; // @[:@14094.4]
  assign RetimeWrapper_22_reset = reset; // @[:@14095.4]
  assign RetimeWrapper_22_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14097.4]
  assign RetimeWrapper_22_io_in = _T_1435 & io_rPort_2_en_0; // @[package.scala 94:16:@14096.4]
  assign RetimeWrapper_23_clock = clock; // @[:@14102.4]
  assign RetimeWrapper_23_reset = reset; // @[:@14103.4]
  assign RetimeWrapper_23_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14105.4]
  assign RetimeWrapper_23_io_in = _T_1559 & io_rPort_2_en_0; // @[package.scala 94:16:@14104.4]
  assign RetimeWrapper_24_clock = clock; // @[:@14142.4]
  assign RetimeWrapper_24_reset = reset; // @[:@14143.4]
  assign RetimeWrapper_24_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14145.4]
  assign RetimeWrapper_24_io_in = _T_629 & io_rPort_3_en_0; // @[package.scala 94:16:@14144.4]
  assign RetimeWrapper_25_clock = clock; // @[:@14150.4]
  assign RetimeWrapper_25_reset = reset; // @[:@14151.4]
  assign RetimeWrapper_25_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14153.4]
  assign RetimeWrapper_25_io_in = _T_753 & io_rPort_3_en_0; // @[package.scala 94:16:@14152.4]
  assign RetimeWrapper_26_clock = clock; // @[:@14158.4]
  assign RetimeWrapper_26_reset = reset; // @[:@14159.4]
  assign RetimeWrapper_26_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14161.4]
  assign RetimeWrapper_26_io_in = _T_877 & io_rPort_3_en_0; // @[package.scala 94:16:@14160.4]
  assign RetimeWrapper_27_clock = clock; // @[:@14166.4]
  assign RetimeWrapper_27_reset = reset; // @[:@14167.4]
  assign RetimeWrapper_27_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14169.4]
  assign RetimeWrapper_27_io_in = _T_1001 & io_rPort_3_en_0; // @[package.scala 94:16:@14168.4]
  assign RetimeWrapper_28_clock = clock; // @[:@14174.4]
  assign RetimeWrapper_28_reset = reset; // @[:@14175.4]
  assign RetimeWrapper_28_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14177.4]
  assign RetimeWrapper_28_io_in = _T_1125 & io_rPort_3_en_0; // @[package.scala 94:16:@14176.4]
  assign RetimeWrapper_29_clock = clock; // @[:@14182.4]
  assign RetimeWrapper_29_reset = reset; // @[:@14183.4]
  assign RetimeWrapper_29_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14185.4]
  assign RetimeWrapper_29_io_in = _T_1249 & io_rPort_3_en_0; // @[package.scala 94:16:@14184.4]
  assign RetimeWrapper_30_clock = clock; // @[:@14190.4]
  assign RetimeWrapper_30_reset = reset; // @[:@14191.4]
  assign RetimeWrapper_30_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14193.4]
  assign RetimeWrapper_30_io_in = _T_1373 & io_rPort_3_en_0; // @[package.scala 94:16:@14192.4]
  assign RetimeWrapper_31_clock = clock; // @[:@14198.4]
  assign RetimeWrapper_31_reset = reset; // @[:@14199.4]
  assign RetimeWrapper_31_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14201.4]
  assign RetimeWrapper_31_io_in = _T_1497 & io_rPort_3_en_0; // @[package.scala 94:16:@14200.4]
  assign RetimeWrapper_32_clock = clock; // @[:@14238.4]
  assign RetimeWrapper_32_reset = reset; // @[:@14239.4]
  assign RetimeWrapper_32_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14241.4]
  assign RetimeWrapper_32_io_in = _T_635 & io_rPort_4_en_0; // @[package.scala 94:16:@14240.4]
  assign RetimeWrapper_33_clock = clock; // @[:@14246.4]
  assign RetimeWrapper_33_reset = reset; // @[:@14247.4]
  assign RetimeWrapper_33_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14249.4]
  assign RetimeWrapper_33_io_in = _T_759 & io_rPort_4_en_0; // @[package.scala 94:16:@14248.4]
  assign RetimeWrapper_34_clock = clock; // @[:@14254.4]
  assign RetimeWrapper_34_reset = reset; // @[:@14255.4]
  assign RetimeWrapper_34_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14257.4]
  assign RetimeWrapper_34_io_in = _T_883 & io_rPort_4_en_0; // @[package.scala 94:16:@14256.4]
  assign RetimeWrapper_35_clock = clock; // @[:@14262.4]
  assign RetimeWrapper_35_reset = reset; // @[:@14263.4]
  assign RetimeWrapper_35_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14265.4]
  assign RetimeWrapper_35_io_in = _T_1007 & io_rPort_4_en_0; // @[package.scala 94:16:@14264.4]
  assign RetimeWrapper_36_clock = clock; // @[:@14270.4]
  assign RetimeWrapper_36_reset = reset; // @[:@14271.4]
  assign RetimeWrapper_36_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14273.4]
  assign RetimeWrapper_36_io_in = _T_1131 & io_rPort_4_en_0; // @[package.scala 94:16:@14272.4]
  assign RetimeWrapper_37_clock = clock; // @[:@14278.4]
  assign RetimeWrapper_37_reset = reset; // @[:@14279.4]
  assign RetimeWrapper_37_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14281.4]
  assign RetimeWrapper_37_io_in = _T_1255 & io_rPort_4_en_0; // @[package.scala 94:16:@14280.4]
  assign RetimeWrapper_38_clock = clock; // @[:@14286.4]
  assign RetimeWrapper_38_reset = reset; // @[:@14287.4]
  assign RetimeWrapper_38_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14289.4]
  assign RetimeWrapper_38_io_in = _T_1379 & io_rPort_4_en_0; // @[package.scala 94:16:@14288.4]
  assign RetimeWrapper_39_clock = clock; // @[:@14294.4]
  assign RetimeWrapper_39_reset = reset; // @[:@14295.4]
  assign RetimeWrapper_39_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14297.4]
  assign RetimeWrapper_39_io_in = _T_1503 & io_rPort_4_en_0; // @[package.scala 94:16:@14296.4]
  assign RetimeWrapper_40_clock = clock; // @[:@14334.4]
  assign RetimeWrapper_40_reset = reset; // @[:@14335.4]
  assign RetimeWrapper_40_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14337.4]
  assign RetimeWrapper_40_io_in = _T_697 & io_rPort_5_en_0; // @[package.scala 94:16:@14336.4]
  assign RetimeWrapper_41_clock = clock; // @[:@14342.4]
  assign RetimeWrapper_41_reset = reset; // @[:@14343.4]
  assign RetimeWrapper_41_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14345.4]
  assign RetimeWrapper_41_io_in = _T_821 & io_rPort_5_en_0; // @[package.scala 94:16:@14344.4]
  assign RetimeWrapper_42_clock = clock; // @[:@14350.4]
  assign RetimeWrapper_42_reset = reset; // @[:@14351.4]
  assign RetimeWrapper_42_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14353.4]
  assign RetimeWrapper_42_io_in = _T_945 & io_rPort_5_en_0; // @[package.scala 94:16:@14352.4]
  assign RetimeWrapper_43_clock = clock; // @[:@14358.4]
  assign RetimeWrapper_43_reset = reset; // @[:@14359.4]
  assign RetimeWrapper_43_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14361.4]
  assign RetimeWrapper_43_io_in = _T_1069 & io_rPort_5_en_0; // @[package.scala 94:16:@14360.4]
  assign RetimeWrapper_44_clock = clock; // @[:@14366.4]
  assign RetimeWrapper_44_reset = reset; // @[:@14367.4]
  assign RetimeWrapper_44_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14369.4]
  assign RetimeWrapper_44_io_in = _T_1193 & io_rPort_5_en_0; // @[package.scala 94:16:@14368.4]
  assign RetimeWrapper_45_clock = clock; // @[:@14374.4]
  assign RetimeWrapper_45_reset = reset; // @[:@14375.4]
  assign RetimeWrapper_45_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14377.4]
  assign RetimeWrapper_45_io_in = _T_1317 & io_rPort_5_en_0; // @[package.scala 94:16:@14376.4]
  assign RetimeWrapper_46_clock = clock; // @[:@14382.4]
  assign RetimeWrapper_46_reset = reset; // @[:@14383.4]
  assign RetimeWrapper_46_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14385.4]
  assign RetimeWrapper_46_io_in = _T_1441 & io_rPort_5_en_0; // @[package.scala 94:16:@14384.4]
  assign RetimeWrapper_47_clock = clock; // @[:@14390.4]
  assign RetimeWrapper_47_reset = reset; // @[:@14391.4]
  assign RetimeWrapper_47_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14393.4]
  assign RetimeWrapper_47_io_in = _T_1565 & io_rPort_5_en_0; // @[package.scala 94:16:@14392.4]
  assign RetimeWrapper_48_clock = clock; // @[:@14430.4]
  assign RetimeWrapper_48_reset = reset; // @[:@14431.4]
  assign RetimeWrapper_48_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14433.4]
  assign RetimeWrapper_48_io_in = _T_641 & io_rPort_6_en_0; // @[package.scala 94:16:@14432.4]
  assign RetimeWrapper_49_clock = clock; // @[:@14438.4]
  assign RetimeWrapper_49_reset = reset; // @[:@14439.4]
  assign RetimeWrapper_49_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14441.4]
  assign RetimeWrapper_49_io_in = _T_765 & io_rPort_6_en_0; // @[package.scala 94:16:@14440.4]
  assign RetimeWrapper_50_clock = clock; // @[:@14446.4]
  assign RetimeWrapper_50_reset = reset; // @[:@14447.4]
  assign RetimeWrapper_50_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14449.4]
  assign RetimeWrapper_50_io_in = _T_889 & io_rPort_6_en_0; // @[package.scala 94:16:@14448.4]
  assign RetimeWrapper_51_clock = clock; // @[:@14454.4]
  assign RetimeWrapper_51_reset = reset; // @[:@14455.4]
  assign RetimeWrapper_51_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14457.4]
  assign RetimeWrapper_51_io_in = _T_1013 & io_rPort_6_en_0; // @[package.scala 94:16:@14456.4]
  assign RetimeWrapper_52_clock = clock; // @[:@14462.4]
  assign RetimeWrapper_52_reset = reset; // @[:@14463.4]
  assign RetimeWrapper_52_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14465.4]
  assign RetimeWrapper_52_io_in = _T_1137 & io_rPort_6_en_0; // @[package.scala 94:16:@14464.4]
  assign RetimeWrapper_53_clock = clock; // @[:@14470.4]
  assign RetimeWrapper_53_reset = reset; // @[:@14471.4]
  assign RetimeWrapper_53_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14473.4]
  assign RetimeWrapper_53_io_in = _T_1261 & io_rPort_6_en_0; // @[package.scala 94:16:@14472.4]
  assign RetimeWrapper_54_clock = clock; // @[:@14478.4]
  assign RetimeWrapper_54_reset = reset; // @[:@14479.4]
  assign RetimeWrapper_54_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14481.4]
  assign RetimeWrapper_54_io_in = _T_1385 & io_rPort_6_en_0; // @[package.scala 94:16:@14480.4]
  assign RetimeWrapper_55_clock = clock; // @[:@14486.4]
  assign RetimeWrapper_55_reset = reset; // @[:@14487.4]
  assign RetimeWrapper_55_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14489.4]
  assign RetimeWrapper_55_io_in = _T_1509 & io_rPort_6_en_0; // @[package.scala 94:16:@14488.4]
  assign RetimeWrapper_56_clock = clock; // @[:@14526.4]
  assign RetimeWrapper_56_reset = reset; // @[:@14527.4]
  assign RetimeWrapper_56_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14529.4]
  assign RetimeWrapper_56_io_in = _T_703 & io_rPort_7_en_0; // @[package.scala 94:16:@14528.4]
  assign RetimeWrapper_57_clock = clock; // @[:@14534.4]
  assign RetimeWrapper_57_reset = reset; // @[:@14535.4]
  assign RetimeWrapper_57_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14537.4]
  assign RetimeWrapper_57_io_in = _T_827 & io_rPort_7_en_0; // @[package.scala 94:16:@14536.4]
  assign RetimeWrapper_58_clock = clock; // @[:@14542.4]
  assign RetimeWrapper_58_reset = reset; // @[:@14543.4]
  assign RetimeWrapper_58_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14545.4]
  assign RetimeWrapper_58_io_in = _T_951 & io_rPort_7_en_0; // @[package.scala 94:16:@14544.4]
  assign RetimeWrapper_59_clock = clock; // @[:@14550.4]
  assign RetimeWrapper_59_reset = reset; // @[:@14551.4]
  assign RetimeWrapper_59_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14553.4]
  assign RetimeWrapper_59_io_in = _T_1075 & io_rPort_7_en_0; // @[package.scala 94:16:@14552.4]
  assign RetimeWrapper_60_clock = clock; // @[:@14558.4]
  assign RetimeWrapper_60_reset = reset; // @[:@14559.4]
  assign RetimeWrapper_60_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14561.4]
  assign RetimeWrapper_60_io_in = _T_1199 & io_rPort_7_en_0; // @[package.scala 94:16:@14560.4]
  assign RetimeWrapper_61_clock = clock; // @[:@14566.4]
  assign RetimeWrapper_61_reset = reset; // @[:@14567.4]
  assign RetimeWrapper_61_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14569.4]
  assign RetimeWrapper_61_io_in = _T_1323 & io_rPort_7_en_0; // @[package.scala 94:16:@14568.4]
  assign RetimeWrapper_62_clock = clock; // @[:@14574.4]
  assign RetimeWrapper_62_reset = reset; // @[:@14575.4]
  assign RetimeWrapper_62_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14577.4]
  assign RetimeWrapper_62_io_in = _T_1447 & io_rPort_7_en_0; // @[package.scala 94:16:@14576.4]
  assign RetimeWrapper_63_clock = clock; // @[:@14582.4]
  assign RetimeWrapper_63_reset = reset; // @[:@14583.4]
  assign RetimeWrapper_63_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14585.4]
  assign RetimeWrapper_63_io_in = _T_1571 & io_rPort_7_en_0; // @[package.scala 94:16:@14584.4]
  assign RetimeWrapper_64_clock = clock; // @[:@14622.4]
  assign RetimeWrapper_64_reset = reset; // @[:@14623.4]
  assign RetimeWrapper_64_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14625.4]
  assign RetimeWrapper_64_io_in = _T_709 & io_rPort_8_en_0; // @[package.scala 94:16:@14624.4]
  assign RetimeWrapper_65_clock = clock; // @[:@14630.4]
  assign RetimeWrapper_65_reset = reset; // @[:@14631.4]
  assign RetimeWrapper_65_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14633.4]
  assign RetimeWrapper_65_io_in = _T_833 & io_rPort_8_en_0; // @[package.scala 94:16:@14632.4]
  assign RetimeWrapper_66_clock = clock; // @[:@14638.4]
  assign RetimeWrapper_66_reset = reset; // @[:@14639.4]
  assign RetimeWrapper_66_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14641.4]
  assign RetimeWrapper_66_io_in = _T_957 & io_rPort_8_en_0; // @[package.scala 94:16:@14640.4]
  assign RetimeWrapper_67_clock = clock; // @[:@14646.4]
  assign RetimeWrapper_67_reset = reset; // @[:@14647.4]
  assign RetimeWrapper_67_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14649.4]
  assign RetimeWrapper_67_io_in = _T_1081 & io_rPort_8_en_0; // @[package.scala 94:16:@14648.4]
  assign RetimeWrapper_68_clock = clock; // @[:@14654.4]
  assign RetimeWrapper_68_reset = reset; // @[:@14655.4]
  assign RetimeWrapper_68_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14657.4]
  assign RetimeWrapper_68_io_in = _T_1205 & io_rPort_8_en_0; // @[package.scala 94:16:@14656.4]
  assign RetimeWrapper_69_clock = clock; // @[:@14662.4]
  assign RetimeWrapper_69_reset = reset; // @[:@14663.4]
  assign RetimeWrapper_69_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14665.4]
  assign RetimeWrapper_69_io_in = _T_1329 & io_rPort_8_en_0; // @[package.scala 94:16:@14664.4]
  assign RetimeWrapper_70_clock = clock; // @[:@14670.4]
  assign RetimeWrapper_70_reset = reset; // @[:@14671.4]
  assign RetimeWrapper_70_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14673.4]
  assign RetimeWrapper_70_io_in = _T_1453 & io_rPort_8_en_0; // @[package.scala 94:16:@14672.4]
  assign RetimeWrapper_71_clock = clock; // @[:@14678.4]
  assign RetimeWrapper_71_reset = reset; // @[:@14679.4]
  assign RetimeWrapper_71_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@14681.4]
  assign RetimeWrapper_71_io_in = _T_1577 & io_rPort_8_en_0; // @[package.scala 94:16:@14680.4]
  assign RetimeWrapper_72_clock = clock; // @[:@14718.4]
  assign RetimeWrapper_72_reset = reset; // @[:@14719.4]
  assign RetimeWrapper_72_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14721.4]
  assign RetimeWrapper_72_io_in = _T_647 & io_rPort_9_en_0; // @[package.scala 94:16:@14720.4]
  assign RetimeWrapper_73_clock = clock; // @[:@14726.4]
  assign RetimeWrapper_73_reset = reset; // @[:@14727.4]
  assign RetimeWrapper_73_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14729.4]
  assign RetimeWrapper_73_io_in = _T_771 & io_rPort_9_en_0; // @[package.scala 94:16:@14728.4]
  assign RetimeWrapper_74_clock = clock; // @[:@14734.4]
  assign RetimeWrapper_74_reset = reset; // @[:@14735.4]
  assign RetimeWrapper_74_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14737.4]
  assign RetimeWrapper_74_io_in = _T_895 & io_rPort_9_en_0; // @[package.scala 94:16:@14736.4]
  assign RetimeWrapper_75_clock = clock; // @[:@14742.4]
  assign RetimeWrapper_75_reset = reset; // @[:@14743.4]
  assign RetimeWrapper_75_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14745.4]
  assign RetimeWrapper_75_io_in = _T_1019 & io_rPort_9_en_0; // @[package.scala 94:16:@14744.4]
  assign RetimeWrapper_76_clock = clock; // @[:@14750.4]
  assign RetimeWrapper_76_reset = reset; // @[:@14751.4]
  assign RetimeWrapper_76_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14753.4]
  assign RetimeWrapper_76_io_in = _T_1143 & io_rPort_9_en_0; // @[package.scala 94:16:@14752.4]
  assign RetimeWrapper_77_clock = clock; // @[:@14758.4]
  assign RetimeWrapper_77_reset = reset; // @[:@14759.4]
  assign RetimeWrapper_77_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14761.4]
  assign RetimeWrapper_77_io_in = _T_1267 & io_rPort_9_en_0; // @[package.scala 94:16:@14760.4]
  assign RetimeWrapper_78_clock = clock; // @[:@14766.4]
  assign RetimeWrapper_78_reset = reset; // @[:@14767.4]
  assign RetimeWrapper_78_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14769.4]
  assign RetimeWrapper_78_io_in = _T_1391 & io_rPort_9_en_0; // @[package.scala 94:16:@14768.4]
  assign RetimeWrapper_79_clock = clock; // @[:@14774.4]
  assign RetimeWrapper_79_reset = reset; // @[:@14775.4]
  assign RetimeWrapper_79_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@14777.4]
  assign RetimeWrapper_79_io_in = _T_1515 & io_rPort_9_en_0; // @[package.scala 94:16:@14776.4]
  assign RetimeWrapper_80_clock = clock; // @[:@14814.4]
  assign RetimeWrapper_80_reset = reset; // @[:@14815.4]
  assign RetimeWrapper_80_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@14817.4]
  assign RetimeWrapper_80_io_in = _T_653 & io_rPort_10_en_0; // @[package.scala 94:16:@14816.4]
  assign RetimeWrapper_81_clock = clock; // @[:@14822.4]
  assign RetimeWrapper_81_reset = reset; // @[:@14823.4]
  assign RetimeWrapper_81_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@14825.4]
  assign RetimeWrapper_81_io_in = _T_777 & io_rPort_10_en_0; // @[package.scala 94:16:@14824.4]
  assign RetimeWrapper_82_clock = clock; // @[:@14830.4]
  assign RetimeWrapper_82_reset = reset; // @[:@14831.4]
  assign RetimeWrapper_82_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@14833.4]
  assign RetimeWrapper_82_io_in = _T_901 & io_rPort_10_en_0; // @[package.scala 94:16:@14832.4]
  assign RetimeWrapper_83_clock = clock; // @[:@14838.4]
  assign RetimeWrapper_83_reset = reset; // @[:@14839.4]
  assign RetimeWrapper_83_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@14841.4]
  assign RetimeWrapper_83_io_in = _T_1025 & io_rPort_10_en_0; // @[package.scala 94:16:@14840.4]
  assign RetimeWrapper_84_clock = clock; // @[:@14846.4]
  assign RetimeWrapper_84_reset = reset; // @[:@14847.4]
  assign RetimeWrapper_84_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@14849.4]
  assign RetimeWrapper_84_io_in = _T_1149 & io_rPort_10_en_0; // @[package.scala 94:16:@14848.4]
  assign RetimeWrapper_85_clock = clock; // @[:@14854.4]
  assign RetimeWrapper_85_reset = reset; // @[:@14855.4]
  assign RetimeWrapper_85_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@14857.4]
  assign RetimeWrapper_85_io_in = _T_1273 & io_rPort_10_en_0; // @[package.scala 94:16:@14856.4]
  assign RetimeWrapper_86_clock = clock; // @[:@14862.4]
  assign RetimeWrapper_86_reset = reset; // @[:@14863.4]
  assign RetimeWrapper_86_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@14865.4]
  assign RetimeWrapper_86_io_in = _T_1397 & io_rPort_10_en_0; // @[package.scala 94:16:@14864.4]
  assign RetimeWrapper_87_clock = clock; // @[:@14870.4]
  assign RetimeWrapper_87_reset = reset; // @[:@14871.4]
  assign RetimeWrapper_87_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@14873.4]
  assign RetimeWrapper_87_io_in = _T_1521 & io_rPort_10_en_0; // @[package.scala 94:16:@14872.4]
  assign RetimeWrapper_88_clock = clock; // @[:@14910.4]
  assign RetimeWrapper_88_reset = reset; // @[:@14911.4]
  assign RetimeWrapper_88_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@14913.4]
  assign RetimeWrapper_88_io_in = _T_715 & io_rPort_11_en_0; // @[package.scala 94:16:@14912.4]
  assign RetimeWrapper_89_clock = clock; // @[:@14918.4]
  assign RetimeWrapper_89_reset = reset; // @[:@14919.4]
  assign RetimeWrapper_89_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@14921.4]
  assign RetimeWrapper_89_io_in = _T_839 & io_rPort_11_en_0; // @[package.scala 94:16:@14920.4]
  assign RetimeWrapper_90_clock = clock; // @[:@14926.4]
  assign RetimeWrapper_90_reset = reset; // @[:@14927.4]
  assign RetimeWrapper_90_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@14929.4]
  assign RetimeWrapper_90_io_in = _T_963 & io_rPort_11_en_0; // @[package.scala 94:16:@14928.4]
  assign RetimeWrapper_91_clock = clock; // @[:@14934.4]
  assign RetimeWrapper_91_reset = reset; // @[:@14935.4]
  assign RetimeWrapper_91_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@14937.4]
  assign RetimeWrapper_91_io_in = _T_1087 & io_rPort_11_en_0; // @[package.scala 94:16:@14936.4]
  assign RetimeWrapper_92_clock = clock; // @[:@14942.4]
  assign RetimeWrapper_92_reset = reset; // @[:@14943.4]
  assign RetimeWrapper_92_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@14945.4]
  assign RetimeWrapper_92_io_in = _T_1211 & io_rPort_11_en_0; // @[package.scala 94:16:@14944.4]
  assign RetimeWrapper_93_clock = clock; // @[:@14950.4]
  assign RetimeWrapper_93_reset = reset; // @[:@14951.4]
  assign RetimeWrapper_93_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@14953.4]
  assign RetimeWrapper_93_io_in = _T_1335 & io_rPort_11_en_0; // @[package.scala 94:16:@14952.4]
  assign RetimeWrapper_94_clock = clock; // @[:@14958.4]
  assign RetimeWrapper_94_reset = reset; // @[:@14959.4]
  assign RetimeWrapper_94_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@14961.4]
  assign RetimeWrapper_94_io_in = _T_1459 & io_rPort_11_en_0; // @[package.scala 94:16:@14960.4]
  assign RetimeWrapper_95_clock = clock; // @[:@14966.4]
  assign RetimeWrapper_95_reset = reset; // @[:@14967.4]
  assign RetimeWrapper_95_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@14969.4]
  assign RetimeWrapper_95_io_in = _T_1583 & io_rPort_11_en_0; // @[package.scala 94:16:@14968.4]
endmodule
module StickySelects_17( // @[:@16693.2]
  input   clock, // @[:@16694.4]
  input   reset, // @[:@16695.4]
  input   io_ins_0, // @[:@16696.4]
  input   io_ins_1, // @[:@16696.4]
  output  io_outs_0, // @[:@16696.4]
  output  io_outs_1 // @[:@16696.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@16698.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@16699.4]
  reg [31:0] _RAND_1;
  wire  _T_23; // @[StickySelects.scala 49:53:@16700.4]
  wire  _T_24; // @[StickySelects.scala 49:21:@16701.4]
  wire  _T_25; // @[StickySelects.scala 49:53:@16703.4]
  wire  _T_26; // @[StickySelects.scala 49:21:@16704.4]
  assign _T_23 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@16700.4]
  assign _T_24 = io_ins_1 ? io_ins_0 : _T_23; // @[StickySelects.scala 49:21:@16701.4]
  assign _T_25 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@16703.4]
  assign _T_26 = io_ins_0 ? io_ins_1 : _T_25; // @[StickySelects.scala 49:21:@16704.4]
  assign io_outs_0 = io_ins_1 ? io_ins_0 : _T_23; // @[StickySelects.scala 53:57:@16706.4]
  assign io_outs_1 = io_ins_0 ? io_ins_1 : _T_25; // @[StickySelects.scala 53:57:@16707.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (io_ins_1) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_23;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (io_ins_0) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_25;
      end
    end
  end
endmodule
module StickySelects_18( // @[:@16709.2]
  input   clock, // @[:@16710.4]
  input   reset, // @[:@16711.4]
  input   io_ins_0, // @[:@16712.4]
  input   io_ins_1, // @[:@16712.4]
  input   io_ins_2, // @[:@16712.4]
  input   io_ins_3, // @[:@16712.4]
  output  io_outs_0, // @[:@16712.4]
  output  io_outs_1, // @[:@16712.4]
  output  io_outs_2, // @[:@16712.4]
  output  io_outs_3 // @[:@16712.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@16714.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@16715.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@16716.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@16717.4]
  reg [31:0] _RAND_3;
  wire  _T_29; // @[StickySelects.scala 47:46:@16718.4]
  wire  _T_30; // @[StickySelects.scala 47:46:@16719.4]
  wire  _T_31; // @[StickySelects.scala 49:53:@16720.4]
  wire  _T_32; // @[StickySelects.scala 49:21:@16721.4]
  wire  _T_33; // @[StickySelects.scala 47:46:@16723.4]
  wire  _T_34; // @[StickySelects.scala 47:46:@16724.4]
  wire  _T_35; // @[StickySelects.scala 49:53:@16725.4]
  wire  _T_36; // @[StickySelects.scala 49:21:@16726.4]
  wire  _T_37; // @[StickySelects.scala 47:46:@16728.4]
  wire  _T_38; // @[StickySelects.scala 47:46:@16729.4]
  wire  _T_39; // @[StickySelects.scala 49:53:@16730.4]
  wire  _T_40; // @[StickySelects.scala 49:21:@16731.4]
  wire  _T_42; // @[StickySelects.scala 47:46:@16734.4]
  wire  _T_43; // @[StickySelects.scala 49:53:@16735.4]
  wire  _T_44; // @[StickySelects.scala 49:21:@16736.4]
  assign _T_29 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@16718.4]
  assign _T_30 = _T_29 | io_ins_3; // @[StickySelects.scala 47:46:@16719.4]
  assign _T_31 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@16720.4]
  assign _T_32 = _T_30 ? io_ins_0 : _T_31; // @[StickySelects.scala 49:21:@16721.4]
  assign _T_33 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@16723.4]
  assign _T_34 = _T_33 | io_ins_3; // @[StickySelects.scala 47:46:@16724.4]
  assign _T_35 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@16725.4]
  assign _T_36 = _T_34 ? io_ins_1 : _T_35; // @[StickySelects.scala 49:21:@16726.4]
  assign _T_37 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@16728.4]
  assign _T_38 = _T_37 | io_ins_3; // @[StickySelects.scala 47:46:@16729.4]
  assign _T_39 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@16730.4]
  assign _T_40 = _T_38 ? io_ins_2 : _T_39; // @[StickySelects.scala 49:21:@16731.4]
  assign _T_42 = _T_37 | io_ins_2; // @[StickySelects.scala 47:46:@16734.4]
  assign _T_43 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@16735.4]
  assign _T_44 = _T_42 ? io_ins_3 : _T_43; // @[StickySelects.scala 49:21:@16736.4]
  assign io_outs_0 = _T_30 ? io_ins_0 : _T_31; // @[StickySelects.scala 53:57:@16738.4]
  assign io_outs_1 = _T_34 ? io_ins_1 : _T_35; // @[StickySelects.scala 53:57:@16739.4]
  assign io_outs_2 = _T_38 ? io_ins_2 : _T_39; // @[StickySelects.scala 53:57:@16740.4]
  assign io_outs_3 = _T_42 ? io_ins_3 : _T_43; // @[StickySelects.scala 53:57:@16741.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_30) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_31;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_34) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_35;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_38) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_39;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_42) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_43;
      end
    end
  end
endmodule
module x286_lb2_0( // @[:@18629.2]
  input         clock, // @[:@18630.4]
  input         reset, // @[:@18631.4]
  input  [2:0]  io_rPort_5_banks_1, // @[:@18632.4]
  input  [2:0]  io_rPort_5_banks_0, // @[:@18632.4]
  input  [8:0]  io_rPort_5_ofs_0, // @[:@18632.4]
  input         io_rPort_5_en_0, // @[:@18632.4]
  input         io_rPort_5_backpressure, // @[:@18632.4]
  output [31:0] io_rPort_5_output_0, // @[:@18632.4]
  input  [2:0]  io_rPort_4_banks_1, // @[:@18632.4]
  input  [2:0]  io_rPort_4_banks_0, // @[:@18632.4]
  input  [8:0]  io_rPort_4_ofs_0, // @[:@18632.4]
  input         io_rPort_4_en_0, // @[:@18632.4]
  input         io_rPort_4_backpressure, // @[:@18632.4]
  output [31:0] io_rPort_4_output_0, // @[:@18632.4]
  input  [2:0]  io_rPort_3_banks_1, // @[:@18632.4]
  input  [2:0]  io_rPort_3_banks_0, // @[:@18632.4]
  input  [8:0]  io_rPort_3_ofs_0, // @[:@18632.4]
  input         io_rPort_3_en_0, // @[:@18632.4]
  input         io_rPort_3_backpressure, // @[:@18632.4]
  output [31:0] io_rPort_3_output_0, // @[:@18632.4]
  input  [2:0]  io_rPort_2_banks_1, // @[:@18632.4]
  input  [2:0]  io_rPort_2_banks_0, // @[:@18632.4]
  input  [8:0]  io_rPort_2_ofs_0, // @[:@18632.4]
  input         io_rPort_2_en_0, // @[:@18632.4]
  input         io_rPort_2_backpressure, // @[:@18632.4]
  output [31:0] io_rPort_2_output_0, // @[:@18632.4]
  input  [2:0]  io_rPort_1_banks_1, // @[:@18632.4]
  input  [2:0]  io_rPort_1_banks_0, // @[:@18632.4]
  input  [8:0]  io_rPort_1_ofs_0, // @[:@18632.4]
  input         io_rPort_1_en_0, // @[:@18632.4]
  input         io_rPort_1_backpressure, // @[:@18632.4]
  output [31:0] io_rPort_1_output_0, // @[:@18632.4]
  input  [2:0]  io_rPort_0_banks_1, // @[:@18632.4]
  input  [2:0]  io_rPort_0_banks_0, // @[:@18632.4]
  input  [8:0]  io_rPort_0_ofs_0, // @[:@18632.4]
  input         io_rPort_0_en_0, // @[:@18632.4]
  input         io_rPort_0_backpressure, // @[:@18632.4]
  output [31:0] io_rPort_0_output_0, // @[:@18632.4]
  input  [2:0]  io_wPort_1_banks_1, // @[:@18632.4]
  input  [2:0]  io_wPort_1_banks_0, // @[:@18632.4]
  input  [8:0]  io_wPort_1_ofs_0, // @[:@18632.4]
  input  [31:0] io_wPort_1_data_0, // @[:@18632.4]
  input         io_wPort_1_en_0, // @[:@18632.4]
  input  [2:0]  io_wPort_0_banks_1, // @[:@18632.4]
  input  [2:0]  io_wPort_0_banks_0, // @[:@18632.4]
  input  [8:0]  io_wPort_0_ofs_0, // @[:@18632.4]
  input  [31:0] io_wPort_0_data_0, // @[:@18632.4]
  input         io_wPort_0_en_0 // @[:@18632.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@18687.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@18687.4]
  wire [8:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18687.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18687.4]
  wire [8:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18687.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@18687.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@18687.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@18687.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@18703.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@18703.4]
  wire [8:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18703.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18703.4]
  wire [8:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18703.4]
  wire [31:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@18703.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@18703.4]
  wire [31:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@18703.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@18719.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@18719.4]
  wire [8:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18719.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18719.4]
  wire [8:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18719.4]
  wire [31:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@18719.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@18719.4]
  wire [31:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@18719.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@18735.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@18735.4]
  wire [8:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18735.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18735.4]
  wire [8:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18735.4]
  wire [31:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@18735.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@18735.4]
  wire [31:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@18735.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@18751.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@18751.4]
  wire [8:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18751.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18751.4]
  wire [8:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18751.4]
  wire [31:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@18751.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@18751.4]
  wire [31:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@18751.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@18767.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@18767.4]
  wire [8:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18767.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18767.4]
  wire [8:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18767.4]
  wire [31:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@18767.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@18767.4]
  wire [31:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@18767.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@18783.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@18783.4]
  wire [8:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18783.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18783.4]
  wire [8:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18783.4]
  wire [31:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@18783.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@18783.4]
  wire [31:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@18783.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@18799.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@18799.4]
  wire [8:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18799.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18799.4]
  wire [8:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18799.4]
  wire [31:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@18799.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@18799.4]
  wire [31:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@18799.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@18815.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@18815.4]
  wire [8:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18815.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18815.4]
  wire [8:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18815.4]
  wire [31:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@18815.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@18815.4]
  wire [31:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@18815.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@18831.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@18831.4]
  wire [8:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18831.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18831.4]
  wire [8:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18831.4]
  wire [31:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@18831.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@18831.4]
  wire [31:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@18831.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@18847.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@18847.4]
  wire [8:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18847.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18847.4]
  wire [8:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18847.4]
  wire [31:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@18847.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@18847.4]
  wire [31:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@18847.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@18863.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@18863.4]
  wire [8:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18863.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18863.4]
  wire [8:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18863.4]
  wire [31:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@18863.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@18863.4]
  wire [31:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@18863.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@18879.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@18879.4]
  wire [8:0] Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18879.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18879.4]
  wire [8:0] Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18879.4]
  wire [31:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@18879.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@18879.4]
  wire [31:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@18879.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@18895.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@18895.4]
  wire [8:0] Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18895.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18895.4]
  wire [8:0] Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18895.4]
  wire [31:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@18895.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@18895.4]
  wire [31:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@18895.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@18911.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@18911.4]
  wire [8:0] Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18911.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18911.4]
  wire [8:0] Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18911.4]
  wire [31:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@18911.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@18911.4]
  wire [31:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@18911.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@18927.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@18927.4]
  wire [8:0] Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@18927.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@18927.4]
  wire [8:0] Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@18927.4]
  wire [31:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@18927.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@18927.4]
  wire [31:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@18927.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@19143.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@19143.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@19143.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@19143.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@19143.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@19143.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 124:33:@19177.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 124:33:@19213.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 124:33:@19213.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 124:33:@19213.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 124:33:@19213.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 124:33:@19213.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 124:33:@19213.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 124:33:@19247.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 124:33:@19283.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 124:33:@19283.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 124:33:@19283.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 124:33:@19283.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 124:33:@19283.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 124:33:@19283.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 124:33:@19317.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 124:33:@19353.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 124:33:@19353.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 124:33:@19353.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 124:33:@19353.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 124:33:@19353.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 124:33:@19353.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 124:33:@19387.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 124:33:@19423.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 124:33:@19423.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 124:33:@19423.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 124:33:@19423.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 124:33:@19423.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 124:33:@19423.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 124:33:@19457.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 124:33:@19493.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 124:33:@19493.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 124:33:@19493.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 124:33:@19493.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 124:33:@19493.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 124:33:@19493.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 124:33:@19527.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 124:33:@19563.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 124:33:@19563.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 124:33:@19563.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 124:33:@19563.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 124:33:@19563.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 124:33:@19563.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 124:33:@19597.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 124:33:@19633.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 124:33:@19633.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 124:33:@19633.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 124:33:@19633.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 124:33:@19633.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 124:33:@19633.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 124:33:@19667.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@19720.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@19720.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@19720.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@19720.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@19720.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@19728.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@19728.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@19728.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@19728.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@19728.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@19736.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@19736.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@19736.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@19736.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@19736.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@19744.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@19744.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@19744.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@19744.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@19744.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@19752.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@19752.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@19752.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@19752.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@19752.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@19760.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@19760.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@19760.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@19760.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@19760.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@19768.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@19768.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@19768.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@19768.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@19768.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@19776.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@19776.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@19776.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@19776.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@19776.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@19816.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@19816.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@19816.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@19816.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@19816.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@19824.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@19824.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@19824.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@19824.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@19824.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@19832.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@19832.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@19832.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@19832.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@19832.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@19840.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@19840.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@19840.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@19840.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@19840.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@19848.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@19848.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@19848.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@19848.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@19848.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@19856.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@19856.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@19856.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@19856.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@19856.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@19864.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@19864.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@19864.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@19864.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@19864.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@19872.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@19872.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@19872.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@19872.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@19872.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@19912.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@19912.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@19912.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@19912.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@19912.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@19920.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@19920.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@19920.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@19920.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@19920.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@19928.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@19928.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@19928.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@19928.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@19928.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@19936.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@19936.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@19936.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@19936.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@19936.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@19944.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@19944.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@19944.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@19944.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@19944.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@19952.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@19952.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@19952.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@19952.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@19952.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@19960.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@19960.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@19960.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@19960.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@19960.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@19968.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@19968.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@19968.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@19968.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@19968.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@20008.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@20008.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@20008.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@20008.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@20008.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@20016.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@20016.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@20016.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@20016.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@20016.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@20024.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@20024.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@20024.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@20024.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@20024.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@20032.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@20032.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@20032.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@20032.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@20032.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@20040.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@20040.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@20040.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@20040.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@20040.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@20048.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@20048.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@20048.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@20048.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@20048.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@20056.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@20056.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@20056.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@20056.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@20056.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@20064.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@20064.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@20064.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@20064.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@20064.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@20104.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@20104.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@20104.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@20104.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@20104.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@20112.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@20112.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@20112.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@20112.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@20112.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@20120.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@20120.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@20120.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@20120.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@20120.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@20128.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@20128.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@20128.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@20128.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@20128.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@20136.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@20136.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@20136.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@20136.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@20136.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@20144.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@20144.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@20144.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@20144.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@20144.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@20152.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@20152.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@20152.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@20152.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@20152.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@20160.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@20160.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@20160.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@20160.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@20160.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@20200.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@20200.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@20200.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@20200.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@20200.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@20208.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@20208.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@20208.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@20208.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@20208.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@20216.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@20216.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@20216.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@20216.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@20216.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@20224.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@20224.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@20224.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@20224.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@20224.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@20232.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@20232.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@20232.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@20232.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@20232.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@20240.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@20240.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@20240.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@20240.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@20240.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@20248.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@20248.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@20248.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@20248.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@20248.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@20256.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@20256.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@20256.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@20256.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@20256.4]
  wire  _T_264; // @[MemPrimitives.scala 82:210:@18943.4]
  wire  _T_266; // @[MemPrimitives.scala 82:210:@18944.4]
  wire  _T_267; // @[MemPrimitives.scala 82:228:@18945.4]
  wire  _T_268; // @[MemPrimitives.scala 83:102:@18946.4]
  wire [41:0] _T_270; // @[Cat.scala 30:58:@18948.4]
  wire  _T_275; // @[MemPrimitives.scala 82:210:@18955.4]
  wire  _T_277; // @[MemPrimitives.scala 82:210:@18956.4]
  wire  _T_278; // @[MemPrimitives.scala 82:228:@18957.4]
  wire  _T_279; // @[MemPrimitives.scala 83:102:@18958.4]
  wire [41:0] _T_281; // @[Cat.scala 30:58:@18960.4]
  wire  _T_288; // @[MemPrimitives.scala 82:210:@18968.4]
  wire  _T_289; // @[MemPrimitives.scala 82:228:@18969.4]
  wire  _T_290; // @[MemPrimitives.scala 83:102:@18970.4]
  wire [41:0] _T_292; // @[Cat.scala 30:58:@18972.4]
  wire  _T_299; // @[MemPrimitives.scala 82:210:@18980.4]
  wire  _T_300; // @[MemPrimitives.scala 82:228:@18981.4]
  wire  _T_301; // @[MemPrimitives.scala 83:102:@18982.4]
  wire [41:0] _T_303; // @[Cat.scala 30:58:@18984.4]
  wire  _T_308; // @[MemPrimitives.scala 82:210:@18991.4]
  wire  _T_311; // @[MemPrimitives.scala 82:228:@18993.4]
  wire  _T_312; // @[MemPrimitives.scala 83:102:@18994.4]
  wire [41:0] _T_314; // @[Cat.scala 30:58:@18996.4]
  wire  _T_319; // @[MemPrimitives.scala 82:210:@19003.4]
  wire  _T_322; // @[MemPrimitives.scala 82:228:@19005.4]
  wire  _T_323; // @[MemPrimitives.scala 83:102:@19006.4]
  wire [41:0] _T_325; // @[Cat.scala 30:58:@19008.4]
  wire  _T_333; // @[MemPrimitives.scala 82:228:@19017.4]
  wire  _T_334; // @[MemPrimitives.scala 83:102:@19018.4]
  wire [41:0] _T_336; // @[Cat.scala 30:58:@19020.4]
  wire  _T_344; // @[MemPrimitives.scala 82:228:@19029.4]
  wire  _T_345; // @[MemPrimitives.scala 83:102:@19030.4]
  wire [41:0] _T_347; // @[Cat.scala 30:58:@19032.4]
  wire  _T_352; // @[MemPrimitives.scala 82:210:@19039.4]
  wire  _T_355; // @[MemPrimitives.scala 82:228:@19041.4]
  wire  _T_356; // @[MemPrimitives.scala 83:102:@19042.4]
  wire [41:0] _T_358; // @[Cat.scala 30:58:@19044.4]
  wire  _T_363; // @[MemPrimitives.scala 82:210:@19051.4]
  wire  _T_366; // @[MemPrimitives.scala 82:228:@19053.4]
  wire  _T_367; // @[MemPrimitives.scala 83:102:@19054.4]
  wire [41:0] _T_369; // @[Cat.scala 30:58:@19056.4]
  wire  _T_377; // @[MemPrimitives.scala 82:228:@19065.4]
  wire  _T_378; // @[MemPrimitives.scala 83:102:@19066.4]
  wire [41:0] _T_380; // @[Cat.scala 30:58:@19068.4]
  wire  _T_388; // @[MemPrimitives.scala 82:228:@19077.4]
  wire  _T_389; // @[MemPrimitives.scala 83:102:@19078.4]
  wire [41:0] _T_391; // @[Cat.scala 30:58:@19080.4]
  wire  _T_396; // @[MemPrimitives.scala 82:210:@19087.4]
  wire  _T_399; // @[MemPrimitives.scala 82:228:@19089.4]
  wire  _T_400; // @[MemPrimitives.scala 83:102:@19090.4]
  wire [41:0] _T_402; // @[Cat.scala 30:58:@19092.4]
  wire  _T_407; // @[MemPrimitives.scala 82:210:@19099.4]
  wire  _T_410; // @[MemPrimitives.scala 82:228:@19101.4]
  wire  _T_411; // @[MemPrimitives.scala 83:102:@19102.4]
  wire [41:0] _T_413; // @[Cat.scala 30:58:@19104.4]
  wire  _T_421; // @[MemPrimitives.scala 82:228:@19113.4]
  wire  _T_422; // @[MemPrimitives.scala 83:102:@19114.4]
  wire [41:0] _T_424; // @[Cat.scala 30:58:@19116.4]
  wire  _T_432; // @[MemPrimitives.scala 82:228:@19125.4]
  wire  _T_433; // @[MemPrimitives.scala 83:102:@19126.4]
  wire [41:0] _T_435; // @[Cat.scala 30:58:@19128.4]
  wire  _T_440; // @[MemPrimitives.scala 110:210:@19135.4]
  wire  _T_442; // @[MemPrimitives.scala 110:210:@19136.4]
  wire  _T_443; // @[MemPrimitives.scala 110:228:@19137.4]
  wire  _T_446; // @[MemPrimitives.scala 110:210:@19139.4]
  wire  _T_448; // @[MemPrimitives.scala 110:210:@19140.4]
  wire  _T_449; // @[MemPrimitives.scala 110:228:@19141.4]
  wire  _T_451; // @[MemPrimitives.scala 126:35:@19148.4]
  wire  _T_452; // @[MemPrimitives.scala 126:35:@19149.4]
  wire [10:0] _T_454; // @[Cat.scala 30:58:@19151.4]
  wire [10:0] _T_456; // @[Cat.scala 30:58:@19153.4]
  wire [10:0] _T_457; // @[Mux.scala 31:69:@19154.4]
  wire  _T_462; // @[MemPrimitives.scala 110:210:@19161.4]
  wire  _T_464; // @[MemPrimitives.scala 110:210:@19162.4]
  wire  _T_465; // @[MemPrimitives.scala 110:228:@19163.4]
  wire  _T_468; // @[MemPrimitives.scala 110:210:@19165.4]
  wire  _T_470; // @[MemPrimitives.scala 110:210:@19166.4]
  wire  _T_471; // @[MemPrimitives.scala 110:228:@19167.4]
  wire  _T_474; // @[MemPrimitives.scala 110:210:@19169.4]
  wire  _T_476; // @[MemPrimitives.scala 110:210:@19170.4]
  wire  _T_477; // @[MemPrimitives.scala 110:228:@19171.4]
  wire  _T_480; // @[MemPrimitives.scala 110:210:@19173.4]
  wire  _T_482; // @[MemPrimitives.scala 110:210:@19174.4]
  wire  _T_483; // @[MemPrimitives.scala 110:228:@19175.4]
  wire  _T_485; // @[MemPrimitives.scala 126:35:@19184.4]
  wire  _T_486; // @[MemPrimitives.scala 126:35:@19185.4]
  wire  _T_487; // @[MemPrimitives.scala 126:35:@19186.4]
  wire  _T_488; // @[MemPrimitives.scala 126:35:@19187.4]
  wire [10:0] _T_490; // @[Cat.scala 30:58:@19189.4]
  wire [10:0] _T_492; // @[Cat.scala 30:58:@19191.4]
  wire [10:0] _T_494; // @[Cat.scala 30:58:@19193.4]
  wire [10:0] _T_496; // @[Cat.scala 30:58:@19195.4]
  wire [10:0] _T_497; // @[Mux.scala 31:69:@19196.4]
  wire [10:0] _T_498; // @[Mux.scala 31:69:@19197.4]
  wire [10:0] _T_499; // @[Mux.scala 31:69:@19198.4]
  wire  _T_506; // @[MemPrimitives.scala 110:210:@19206.4]
  wire  _T_507; // @[MemPrimitives.scala 110:228:@19207.4]
  wire  _T_512; // @[MemPrimitives.scala 110:210:@19210.4]
  wire  _T_513; // @[MemPrimitives.scala 110:228:@19211.4]
  wire  _T_515; // @[MemPrimitives.scala 126:35:@19218.4]
  wire  _T_516; // @[MemPrimitives.scala 126:35:@19219.4]
  wire [10:0] _T_518; // @[Cat.scala 30:58:@19221.4]
  wire [10:0] _T_520; // @[Cat.scala 30:58:@19223.4]
  wire [10:0] _T_521; // @[Mux.scala 31:69:@19224.4]
  wire  _T_528; // @[MemPrimitives.scala 110:210:@19232.4]
  wire  _T_529; // @[MemPrimitives.scala 110:228:@19233.4]
  wire  _T_534; // @[MemPrimitives.scala 110:210:@19236.4]
  wire  _T_535; // @[MemPrimitives.scala 110:228:@19237.4]
  wire  _T_540; // @[MemPrimitives.scala 110:210:@19240.4]
  wire  _T_541; // @[MemPrimitives.scala 110:228:@19241.4]
  wire  _T_546; // @[MemPrimitives.scala 110:210:@19244.4]
  wire  _T_547; // @[MemPrimitives.scala 110:228:@19245.4]
  wire  _T_549; // @[MemPrimitives.scala 126:35:@19254.4]
  wire  _T_550; // @[MemPrimitives.scala 126:35:@19255.4]
  wire  _T_551; // @[MemPrimitives.scala 126:35:@19256.4]
  wire  _T_552; // @[MemPrimitives.scala 126:35:@19257.4]
  wire [10:0] _T_554; // @[Cat.scala 30:58:@19259.4]
  wire [10:0] _T_556; // @[Cat.scala 30:58:@19261.4]
  wire [10:0] _T_558; // @[Cat.scala 30:58:@19263.4]
  wire [10:0] _T_560; // @[Cat.scala 30:58:@19265.4]
  wire [10:0] _T_561; // @[Mux.scala 31:69:@19266.4]
  wire [10:0] _T_562; // @[Mux.scala 31:69:@19267.4]
  wire [10:0] _T_563; // @[Mux.scala 31:69:@19268.4]
  wire  _T_568; // @[MemPrimitives.scala 110:210:@19275.4]
  wire  _T_571; // @[MemPrimitives.scala 110:228:@19277.4]
  wire  _T_574; // @[MemPrimitives.scala 110:210:@19279.4]
  wire  _T_577; // @[MemPrimitives.scala 110:228:@19281.4]
  wire  _T_579; // @[MemPrimitives.scala 126:35:@19288.4]
  wire  _T_580; // @[MemPrimitives.scala 126:35:@19289.4]
  wire [10:0] _T_582; // @[Cat.scala 30:58:@19291.4]
  wire [10:0] _T_584; // @[Cat.scala 30:58:@19293.4]
  wire [10:0] _T_585; // @[Mux.scala 31:69:@19294.4]
  wire  _T_590; // @[MemPrimitives.scala 110:210:@19301.4]
  wire  _T_593; // @[MemPrimitives.scala 110:228:@19303.4]
  wire  _T_596; // @[MemPrimitives.scala 110:210:@19305.4]
  wire  _T_599; // @[MemPrimitives.scala 110:228:@19307.4]
  wire  _T_602; // @[MemPrimitives.scala 110:210:@19309.4]
  wire  _T_605; // @[MemPrimitives.scala 110:228:@19311.4]
  wire  _T_608; // @[MemPrimitives.scala 110:210:@19313.4]
  wire  _T_611; // @[MemPrimitives.scala 110:228:@19315.4]
  wire  _T_613; // @[MemPrimitives.scala 126:35:@19324.4]
  wire  _T_614; // @[MemPrimitives.scala 126:35:@19325.4]
  wire  _T_615; // @[MemPrimitives.scala 126:35:@19326.4]
  wire  _T_616; // @[MemPrimitives.scala 126:35:@19327.4]
  wire [10:0] _T_618; // @[Cat.scala 30:58:@19329.4]
  wire [10:0] _T_620; // @[Cat.scala 30:58:@19331.4]
  wire [10:0] _T_622; // @[Cat.scala 30:58:@19333.4]
  wire [10:0] _T_624; // @[Cat.scala 30:58:@19335.4]
  wire [10:0] _T_625; // @[Mux.scala 31:69:@19336.4]
  wire [10:0] _T_626; // @[Mux.scala 31:69:@19337.4]
  wire [10:0] _T_627; // @[Mux.scala 31:69:@19338.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@19347.4]
  wire  _T_641; // @[MemPrimitives.scala 110:228:@19351.4]
  wire  _T_643; // @[MemPrimitives.scala 126:35:@19358.4]
  wire  _T_644; // @[MemPrimitives.scala 126:35:@19359.4]
  wire [10:0] _T_646; // @[Cat.scala 30:58:@19361.4]
  wire [10:0] _T_648; // @[Cat.scala 30:58:@19363.4]
  wire [10:0] _T_649; // @[Mux.scala 31:69:@19364.4]
  wire  _T_657; // @[MemPrimitives.scala 110:228:@19373.4]
  wire  _T_663; // @[MemPrimitives.scala 110:228:@19377.4]
  wire  _T_669; // @[MemPrimitives.scala 110:228:@19381.4]
  wire  _T_675; // @[MemPrimitives.scala 110:228:@19385.4]
  wire  _T_677; // @[MemPrimitives.scala 126:35:@19394.4]
  wire  _T_678; // @[MemPrimitives.scala 126:35:@19395.4]
  wire  _T_679; // @[MemPrimitives.scala 126:35:@19396.4]
  wire  _T_680; // @[MemPrimitives.scala 126:35:@19397.4]
  wire [10:0] _T_682; // @[Cat.scala 30:58:@19399.4]
  wire [10:0] _T_684; // @[Cat.scala 30:58:@19401.4]
  wire [10:0] _T_686; // @[Cat.scala 30:58:@19403.4]
  wire [10:0] _T_688; // @[Cat.scala 30:58:@19405.4]
  wire [10:0] _T_689; // @[Mux.scala 31:69:@19406.4]
  wire [10:0] _T_690; // @[Mux.scala 31:69:@19407.4]
  wire [10:0] _T_691; // @[Mux.scala 31:69:@19408.4]
  wire  _T_696; // @[MemPrimitives.scala 110:210:@19415.4]
  wire  _T_699; // @[MemPrimitives.scala 110:228:@19417.4]
  wire  _T_702; // @[MemPrimitives.scala 110:210:@19419.4]
  wire  _T_705; // @[MemPrimitives.scala 110:228:@19421.4]
  wire  _T_707; // @[MemPrimitives.scala 126:35:@19428.4]
  wire  _T_708; // @[MemPrimitives.scala 126:35:@19429.4]
  wire [10:0] _T_710; // @[Cat.scala 30:58:@19431.4]
  wire [10:0] _T_712; // @[Cat.scala 30:58:@19433.4]
  wire [10:0] _T_713; // @[Mux.scala 31:69:@19434.4]
  wire  _T_718; // @[MemPrimitives.scala 110:210:@19441.4]
  wire  _T_721; // @[MemPrimitives.scala 110:228:@19443.4]
  wire  _T_724; // @[MemPrimitives.scala 110:210:@19445.4]
  wire  _T_727; // @[MemPrimitives.scala 110:228:@19447.4]
  wire  _T_730; // @[MemPrimitives.scala 110:210:@19449.4]
  wire  _T_733; // @[MemPrimitives.scala 110:228:@19451.4]
  wire  _T_736; // @[MemPrimitives.scala 110:210:@19453.4]
  wire  _T_739; // @[MemPrimitives.scala 110:228:@19455.4]
  wire  _T_741; // @[MemPrimitives.scala 126:35:@19464.4]
  wire  _T_742; // @[MemPrimitives.scala 126:35:@19465.4]
  wire  _T_743; // @[MemPrimitives.scala 126:35:@19466.4]
  wire  _T_744; // @[MemPrimitives.scala 126:35:@19467.4]
  wire [10:0] _T_746; // @[Cat.scala 30:58:@19469.4]
  wire [10:0] _T_748; // @[Cat.scala 30:58:@19471.4]
  wire [10:0] _T_750; // @[Cat.scala 30:58:@19473.4]
  wire [10:0] _T_752; // @[Cat.scala 30:58:@19475.4]
  wire [10:0] _T_753; // @[Mux.scala 31:69:@19476.4]
  wire [10:0] _T_754; // @[Mux.scala 31:69:@19477.4]
  wire [10:0] _T_755; // @[Mux.scala 31:69:@19478.4]
  wire  _T_763; // @[MemPrimitives.scala 110:228:@19487.4]
  wire  _T_769; // @[MemPrimitives.scala 110:228:@19491.4]
  wire  _T_771; // @[MemPrimitives.scala 126:35:@19498.4]
  wire  _T_772; // @[MemPrimitives.scala 126:35:@19499.4]
  wire [10:0] _T_774; // @[Cat.scala 30:58:@19501.4]
  wire [10:0] _T_776; // @[Cat.scala 30:58:@19503.4]
  wire [10:0] _T_777; // @[Mux.scala 31:69:@19504.4]
  wire  _T_785; // @[MemPrimitives.scala 110:228:@19513.4]
  wire  _T_791; // @[MemPrimitives.scala 110:228:@19517.4]
  wire  _T_797; // @[MemPrimitives.scala 110:228:@19521.4]
  wire  _T_803; // @[MemPrimitives.scala 110:228:@19525.4]
  wire  _T_805; // @[MemPrimitives.scala 126:35:@19534.4]
  wire  _T_806; // @[MemPrimitives.scala 126:35:@19535.4]
  wire  _T_807; // @[MemPrimitives.scala 126:35:@19536.4]
  wire  _T_808; // @[MemPrimitives.scala 126:35:@19537.4]
  wire [10:0] _T_810; // @[Cat.scala 30:58:@19539.4]
  wire [10:0] _T_812; // @[Cat.scala 30:58:@19541.4]
  wire [10:0] _T_814; // @[Cat.scala 30:58:@19543.4]
  wire [10:0] _T_816; // @[Cat.scala 30:58:@19545.4]
  wire [10:0] _T_817; // @[Mux.scala 31:69:@19546.4]
  wire [10:0] _T_818; // @[Mux.scala 31:69:@19547.4]
  wire [10:0] _T_819; // @[Mux.scala 31:69:@19548.4]
  wire  _T_824; // @[MemPrimitives.scala 110:210:@19555.4]
  wire  _T_827; // @[MemPrimitives.scala 110:228:@19557.4]
  wire  _T_830; // @[MemPrimitives.scala 110:210:@19559.4]
  wire  _T_833; // @[MemPrimitives.scala 110:228:@19561.4]
  wire  _T_835; // @[MemPrimitives.scala 126:35:@19568.4]
  wire  _T_836; // @[MemPrimitives.scala 126:35:@19569.4]
  wire [10:0] _T_838; // @[Cat.scala 30:58:@19571.4]
  wire [10:0] _T_840; // @[Cat.scala 30:58:@19573.4]
  wire [10:0] _T_841; // @[Mux.scala 31:69:@19574.4]
  wire  _T_846; // @[MemPrimitives.scala 110:210:@19581.4]
  wire  _T_849; // @[MemPrimitives.scala 110:228:@19583.4]
  wire  _T_852; // @[MemPrimitives.scala 110:210:@19585.4]
  wire  _T_855; // @[MemPrimitives.scala 110:228:@19587.4]
  wire  _T_858; // @[MemPrimitives.scala 110:210:@19589.4]
  wire  _T_861; // @[MemPrimitives.scala 110:228:@19591.4]
  wire  _T_864; // @[MemPrimitives.scala 110:210:@19593.4]
  wire  _T_867; // @[MemPrimitives.scala 110:228:@19595.4]
  wire  _T_869; // @[MemPrimitives.scala 126:35:@19604.4]
  wire  _T_870; // @[MemPrimitives.scala 126:35:@19605.4]
  wire  _T_871; // @[MemPrimitives.scala 126:35:@19606.4]
  wire  _T_872; // @[MemPrimitives.scala 126:35:@19607.4]
  wire [10:0] _T_874; // @[Cat.scala 30:58:@19609.4]
  wire [10:0] _T_876; // @[Cat.scala 30:58:@19611.4]
  wire [10:0] _T_878; // @[Cat.scala 30:58:@19613.4]
  wire [10:0] _T_880; // @[Cat.scala 30:58:@19615.4]
  wire [10:0] _T_881; // @[Mux.scala 31:69:@19616.4]
  wire [10:0] _T_882; // @[Mux.scala 31:69:@19617.4]
  wire [10:0] _T_883; // @[Mux.scala 31:69:@19618.4]
  wire  _T_891; // @[MemPrimitives.scala 110:228:@19627.4]
  wire  _T_897; // @[MemPrimitives.scala 110:228:@19631.4]
  wire  _T_899; // @[MemPrimitives.scala 126:35:@19638.4]
  wire  _T_900; // @[MemPrimitives.scala 126:35:@19639.4]
  wire [10:0] _T_902; // @[Cat.scala 30:58:@19641.4]
  wire [10:0] _T_904; // @[Cat.scala 30:58:@19643.4]
  wire [10:0] _T_905; // @[Mux.scala 31:69:@19644.4]
  wire  _T_913; // @[MemPrimitives.scala 110:228:@19653.4]
  wire  _T_919; // @[MemPrimitives.scala 110:228:@19657.4]
  wire  _T_925; // @[MemPrimitives.scala 110:228:@19661.4]
  wire  _T_931; // @[MemPrimitives.scala 110:228:@19665.4]
  wire  _T_933; // @[MemPrimitives.scala 126:35:@19674.4]
  wire  _T_934; // @[MemPrimitives.scala 126:35:@19675.4]
  wire  _T_935; // @[MemPrimitives.scala 126:35:@19676.4]
  wire  _T_936; // @[MemPrimitives.scala 126:35:@19677.4]
  wire [10:0] _T_938; // @[Cat.scala 30:58:@19679.4]
  wire [10:0] _T_940; // @[Cat.scala 30:58:@19681.4]
  wire [10:0] _T_942; // @[Cat.scala 30:58:@19683.4]
  wire [10:0] _T_944; // @[Cat.scala 30:58:@19685.4]
  wire [10:0] _T_945; // @[Mux.scala 31:69:@19686.4]
  wire [10:0] _T_946; // @[Mux.scala 31:69:@19687.4]
  wire [10:0] _T_947; // @[Mux.scala 31:69:@19688.4]
  wire  _T_1011; // @[package.scala 96:25:@19773.4 package.scala 96:25:@19774.4]
  wire [31:0] _T_1015; // @[Mux.scala 31:69:@19783.4]
  wire  _T_1008; // @[package.scala 96:25:@19765.4 package.scala 96:25:@19766.4]
  wire [31:0] _T_1016; // @[Mux.scala 31:69:@19784.4]
  wire  _T_1005; // @[package.scala 96:25:@19757.4 package.scala 96:25:@19758.4]
  wire [31:0] _T_1017; // @[Mux.scala 31:69:@19785.4]
  wire  _T_1002; // @[package.scala 96:25:@19749.4 package.scala 96:25:@19750.4]
  wire [31:0] _T_1018; // @[Mux.scala 31:69:@19786.4]
  wire  _T_999; // @[package.scala 96:25:@19741.4 package.scala 96:25:@19742.4]
  wire [31:0] _T_1019; // @[Mux.scala 31:69:@19787.4]
  wire  _T_996; // @[package.scala 96:25:@19733.4 package.scala 96:25:@19734.4]
  wire [31:0] _T_1020; // @[Mux.scala 31:69:@19788.4]
  wire  _T_993; // @[package.scala 96:25:@19725.4 package.scala 96:25:@19726.4]
  wire  _T_1082; // @[package.scala 96:25:@19869.4 package.scala 96:25:@19870.4]
  wire [31:0] _T_1086; // @[Mux.scala 31:69:@19879.4]
  wire  _T_1079; // @[package.scala 96:25:@19861.4 package.scala 96:25:@19862.4]
  wire [31:0] _T_1087; // @[Mux.scala 31:69:@19880.4]
  wire  _T_1076; // @[package.scala 96:25:@19853.4 package.scala 96:25:@19854.4]
  wire [31:0] _T_1088; // @[Mux.scala 31:69:@19881.4]
  wire  _T_1073; // @[package.scala 96:25:@19845.4 package.scala 96:25:@19846.4]
  wire [31:0] _T_1089; // @[Mux.scala 31:69:@19882.4]
  wire  _T_1070; // @[package.scala 96:25:@19837.4 package.scala 96:25:@19838.4]
  wire [31:0] _T_1090; // @[Mux.scala 31:69:@19883.4]
  wire  _T_1067; // @[package.scala 96:25:@19829.4 package.scala 96:25:@19830.4]
  wire [31:0] _T_1091; // @[Mux.scala 31:69:@19884.4]
  wire  _T_1064; // @[package.scala 96:25:@19821.4 package.scala 96:25:@19822.4]
  wire  _T_1153; // @[package.scala 96:25:@19965.4 package.scala 96:25:@19966.4]
  wire [31:0] _T_1157; // @[Mux.scala 31:69:@19975.4]
  wire  _T_1150; // @[package.scala 96:25:@19957.4 package.scala 96:25:@19958.4]
  wire [31:0] _T_1158; // @[Mux.scala 31:69:@19976.4]
  wire  _T_1147; // @[package.scala 96:25:@19949.4 package.scala 96:25:@19950.4]
  wire [31:0] _T_1159; // @[Mux.scala 31:69:@19977.4]
  wire  _T_1144; // @[package.scala 96:25:@19941.4 package.scala 96:25:@19942.4]
  wire [31:0] _T_1160; // @[Mux.scala 31:69:@19978.4]
  wire  _T_1141; // @[package.scala 96:25:@19933.4 package.scala 96:25:@19934.4]
  wire [31:0] _T_1161; // @[Mux.scala 31:69:@19979.4]
  wire  _T_1138; // @[package.scala 96:25:@19925.4 package.scala 96:25:@19926.4]
  wire [31:0] _T_1162; // @[Mux.scala 31:69:@19980.4]
  wire  _T_1135; // @[package.scala 96:25:@19917.4 package.scala 96:25:@19918.4]
  wire  _T_1224; // @[package.scala 96:25:@20061.4 package.scala 96:25:@20062.4]
  wire [31:0] _T_1228; // @[Mux.scala 31:69:@20071.4]
  wire  _T_1221; // @[package.scala 96:25:@20053.4 package.scala 96:25:@20054.4]
  wire [31:0] _T_1229; // @[Mux.scala 31:69:@20072.4]
  wire  _T_1218; // @[package.scala 96:25:@20045.4 package.scala 96:25:@20046.4]
  wire [31:0] _T_1230; // @[Mux.scala 31:69:@20073.4]
  wire  _T_1215; // @[package.scala 96:25:@20037.4 package.scala 96:25:@20038.4]
  wire [31:0] _T_1231; // @[Mux.scala 31:69:@20074.4]
  wire  _T_1212; // @[package.scala 96:25:@20029.4 package.scala 96:25:@20030.4]
  wire [31:0] _T_1232; // @[Mux.scala 31:69:@20075.4]
  wire  _T_1209; // @[package.scala 96:25:@20021.4 package.scala 96:25:@20022.4]
  wire [31:0] _T_1233; // @[Mux.scala 31:69:@20076.4]
  wire  _T_1206; // @[package.scala 96:25:@20013.4 package.scala 96:25:@20014.4]
  wire  _T_1295; // @[package.scala 96:25:@20157.4 package.scala 96:25:@20158.4]
  wire [31:0] _T_1299; // @[Mux.scala 31:69:@20167.4]
  wire  _T_1292; // @[package.scala 96:25:@20149.4 package.scala 96:25:@20150.4]
  wire [31:0] _T_1300; // @[Mux.scala 31:69:@20168.4]
  wire  _T_1289; // @[package.scala 96:25:@20141.4 package.scala 96:25:@20142.4]
  wire [31:0] _T_1301; // @[Mux.scala 31:69:@20169.4]
  wire  _T_1286; // @[package.scala 96:25:@20133.4 package.scala 96:25:@20134.4]
  wire [31:0] _T_1302; // @[Mux.scala 31:69:@20170.4]
  wire  _T_1283; // @[package.scala 96:25:@20125.4 package.scala 96:25:@20126.4]
  wire [31:0] _T_1303; // @[Mux.scala 31:69:@20171.4]
  wire  _T_1280; // @[package.scala 96:25:@20117.4 package.scala 96:25:@20118.4]
  wire [31:0] _T_1304; // @[Mux.scala 31:69:@20172.4]
  wire  _T_1277; // @[package.scala 96:25:@20109.4 package.scala 96:25:@20110.4]
  wire  _T_1366; // @[package.scala 96:25:@20253.4 package.scala 96:25:@20254.4]
  wire [31:0] _T_1370; // @[Mux.scala 31:69:@20263.4]
  wire  _T_1363; // @[package.scala 96:25:@20245.4 package.scala 96:25:@20246.4]
  wire [31:0] _T_1371; // @[Mux.scala 31:69:@20264.4]
  wire  _T_1360; // @[package.scala 96:25:@20237.4 package.scala 96:25:@20238.4]
  wire [31:0] _T_1372; // @[Mux.scala 31:69:@20265.4]
  wire  _T_1357; // @[package.scala 96:25:@20229.4 package.scala 96:25:@20230.4]
  wire [31:0] _T_1373; // @[Mux.scala 31:69:@20266.4]
  wire  _T_1354; // @[package.scala 96:25:@20221.4 package.scala 96:25:@20222.4]
  wire [31:0] _T_1374; // @[Mux.scala 31:69:@20267.4]
  wire  _T_1351; // @[package.scala 96:25:@20213.4 package.scala 96:25:@20214.4]
  wire [31:0] _T_1375; // @[Mux.scala 31:69:@20268.4]
  wire  _T_1348; // @[package.scala 96:25:@20205.4 package.scala 96:25:@20206.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@18687.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@18703.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@18719.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@18735.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@18751.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@18767.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@18783.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@18799.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@18815.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@18831.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@18847.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@18863.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_5 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@18879.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_5 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@18895.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_5 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@18911.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_5 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@18927.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects_17 StickySelects ( // @[MemPrimitives.scala 124:33:@19143.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1)
  );
  StickySelects_18 StickySelects_1 ( // @[MemPrimitives.scala 124:33:@19177.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3)
  );
  StickySelects_17 StickySelects_2 ( // @[MemPrimitives.scala 124:33:@19213.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1)
  );
  StickySelects_18 StickySelects_3 ( // @[MemPrimitives.scala 124:33:@19247.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3)
  );
  StickySelects_17 StickySelects_4 ( // @[MemPrimitives.scala 124:33:@19283.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1)
  );
  StickySelects_18 StickySelects_5 ( // @[MemPrimitives.scala 124:33:@19317.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3)
  );
  StickySelects_17 StickySelects_6 ( // @[MemPrimitives.scala 124:33:@19353.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1)
  );
  StickySelects_18 StickySelects_7 ( // @[MemPrimitives.scala 124:33:@19387.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3)
  );
  StickySelects_17 StickySelects_8 ( // @[MemPrimitives.scala 124:33:@19423.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1)
  );
  StickySelects_18 StickySelects_9 ( // @[MemPrimitives.scala 124:33:@19457.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3)
  );
  StickySelects_17 StickySelects_10 ( // @[MemPrimitives.scala 124:33:@19493.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1)
  );
  StickySelects_18 StickySelects_11 ( // @[MemPrimitives.scala 124:33:@19527.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3)
  );
  StickySelects_17 StickySelects_12 ( // @[MemPrimitives.scala 124:33:@19563.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1)
  );
  StickySelects_18 StickySelects_13 ( // @[MemPrimitives.scala 124:33:@19597.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3)
  );
  StickySelects_17 StickySelects_14 ( // @[MemPrimitives.scala 124:33:@19633.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1)
  );
  StickySelects_18 StickySelects_15 ( // @[MemPrimitives.scala 124:33:@19667.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@19720.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@19728.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@19736.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@19744.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@19752.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@19760.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@19768.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@19776.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@19816.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@19824.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@19832.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@19840.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@19848.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@19856.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@19864.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@19872.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@19912.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@19920.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@19928.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@19936.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@19944.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@19952.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@19960.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@19968.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@20008.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@20016.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@20024.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@20032.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@20040.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@20048.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@20056.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@20064.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@20104.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@20112.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@20120.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@20128.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@20136.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@20144.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@20152.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@20160.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@20200.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@20208.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@20216.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@20224.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@20232.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@20240.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@20248.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@20256.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  assign _T_264 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@18943.4]
  assign _T_266 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@18944.4]
  assign _T_267 = _T_264 & _T_266; // @[MemPrimitives.scala 82:228:@18945.4]
  assign _T_268 = io_wPort_0_en_0 & _T_267; // @[MemPrimitives.scala 83:102:@18946.4]
  assign _T_270 = {_T_268,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18948.4]
  assign _T_275 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@18955.4]
  assign _T_277 = io_wPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@18956.4]
  assign _T_278 = _T_275 & _T_277; // @[MemPrimitives.scala 82:228:@18957.4]
  assign _T_279 = io_wPort_1_en_0 & _T_278; // @[MemPrimitives.scala 83:102:@18958.4]
  assign _T_281 = {_T_279,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@18960.4]
  assign _T_288 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@18968.4]
  assign _T_289 = _T_264 & _T_288; // @[MemPrimitives.scala 82:228:@18969.4]
  assign _T_290 = io_wPort_0_en_0 & _T_289; // @[MemPrimitives.scala 83:102:@18970.4]
  assign _T_292 = {_T_290,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18972.4]
  assign _T_299 = io_wPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@18980.4]
  assign _T_300 = _T_275 & _T_299; // @[MemPrimitives.scala 82:228:@18981.4]
  assign _T_301 = io_wPort_1_en_0 & _T_300; // @[MemPrimitives.scala 83:102:@18982.4]
  assign _T_303 = {_T_301,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@18984.4]
  assign _T_308 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@18991.4]
  assign _T_311 = _T_308 & _T_266; // @[MemPrimitives.scala 82:228:@18993.4]
  assign _T_312 = io_wPort_0_en_0 & _T_311; // @[MemPrimitives.scala 83:102:@18994.4]
  assign _T_314 = {_T_312,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@18996.4]
  assign _T_319 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@19003.4]
  assign _T_322 = _T_319 & _T_277; // @[MemPrimitives.scala 82:228:@19005.4]
  assign _T_323 = io_wPort_1_en_0 & _T_322; // @[MemPrimitives.scala 83:102:@19006.4]
  assign _T_325 = {_T_323,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@19008.4]
  assign _T_333 = _T_308 & _T_288; // @[MemPrimitives.scala 82:228:@19017.4]
  assign _T_334 = io_wPort_0_en_0 & _T_333; // @[MemPrimitives.scala 83:102:@19018.4]
  assign _T_336 = {_T_334,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@19020.4]
  assign _T_344 = _T_319 & _T_299; // @[MemPrimitives.scala 82:228:@19029.4]
  assign _T_345 = io_wPort_1_en_0 & _T_344; // @[MemPrimitives.scala 83:102:@19030.4]
  assign _T_347 = {_T_345,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@19032.4]
  assign _T_352 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@19039.4]
  assign _T_355 = _T_352 & _T_266; // @[MemPrimitives.scala 82:228:@19041.4]
  assign _T_356 = io_wPort_0_en_0 & _T_355; // @[MemPrimitives.scala 83:102:@19042.4]
  assign _T_358 = {_T_356,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@19044.4]
  assign _T_363 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@19051.4]
  assign _T_366 = _T_363 & _T_277; // @[MemPrimitives.scala 82:228:@19053.4]
  assign _T_367 = io_wPort_1_en_0 & _T_366; // @[MemPrimitives.scala 83:102:@19054.4]
  assign _T_369 = {_T_367,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@19056.4]
  assign _T_377 = _T_352 & _T_288; // @[MemPrimitives.scala 82:228:@19065.4]
  assign _T_378 = io_wPort_0_en_0 & _T_377; // @[MemPrimitives.scala 83:102:@19066.4]
  assign _T_380 = {_T_378,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@19068.4]
  assign _T_388 = _T_363 & _T_299; // @[MemPrimitives.scala 82:228:@19077.4]
  assign _T_389 = io_wPort_1_en_0 & _T_388; // @[MemPrimitives.scala 83:102:@19078.4]
  assign _T_391 = {_T_389,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@19080.4]
  assign _T_396 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@19087.4]
  assign _T_399 = _T_396 & _T_266; // @[MemPrimitives.scala 82:228:@19089.4]
  assign _T_400 = io_wPort_0_en_0 & _T_399; // @[MemPrimitives.scala 83:102:@19090.4]
  assign _T_402 = {_T_400,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@19092.4]
  assign _T_407 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@19099.4]
  assign _T_410 = _T_407 & _T_277; // @[MemPrimitives.scala 82:228:@19101.4]
  assign _T_411 = io_wPort_1_en_0 & _T_410; // @[MemPrimitives.scala 83:102:@19102.4]
  assign _T_413 = {_T_411,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@19104.4]
  assign _T_421 = _T_396 & _T_288; // @[MemPrimitives.scala 82:228:@19113.4]
  assign _T_422 = io_wPort_0_en_0 & _T_421; // @[MemPrimitives.scala 83:102:@19114.4]
  assign _T_424 = {_T_422,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@19116.4]
  assign _T_432 = _T_407 & _T_299; // @[MemPrimitives.scala 82:228:@19125.4]
  assign _T_433 = io_wPort_1_en_0 & _T_432; // @[MemPrimitives.scala 83:102:@19126.4]
  assign _T_435 = {_T_433,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@19128.4]
  assign _T_440 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@19135.4]
  assign _T_442 = io_rPort_3_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@19136.4]
  assign _T_443 = _T_440 & _T_442; // @[MemPrimitives.scala 110:228:@19137.4]
  assign _T_446 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@19139.4]
  assign _T_448 = io_rPort_5_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@19140.4]
  assign _T_449 = _T_446 & _T_448; // @[MemPrimitives.scala 110:228:@19141.4]
  assign _T_451 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@19148.4]
  assign _T_452 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@19149.4]
  assign _T_454 = {_T_451,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19151.4]
  assign _T_456 = {_T_452,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@19153.4]
  assign _T_457 = _T_451 ? _T_454 : _T_456; // @[Mux.scala 31:69:@19154.4]
  assign _T_462 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@19161.4]
  assign _T_464 = io_rPort_0_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@19162.4]
  assign _T_465 = _T_462 & _T_464; // @[MemPrimitives.scala 110:228:@19163.4]
  assign _T_468 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@19165.4]
  assign _T_470 = io_rPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@19166.4]
  assign _T_471 = _T_468 & _T_470; // @[MemPrimitives.scala 110:228:@19167.4]
  assign _T_474 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@19169.4]
  assign _T_476 = io_rPort_2_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@19170.4]
  assign _T_477 = _T_474 & _T_476; // @[MemPrimitives.scala 110:228:@19171.4]
  assign _T_480 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@19173.4]
  assign _T_482 = io_rPort_4_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@19174.4]
  assign _T_483 = _T_480 & _T_482; // @[MemPrimitives.scala 110:228:@19175.4]
  assign _T_485 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 126:35:@19184.4]
  assign _T_486 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 126:35:@19185.4]
  assign _T_487 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 126:35:@19186.4]
  assign _T_488 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 126:35:@19187.4]
  assign _T_490 = {_T_485,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19189.4]
  assign _T_492 = {_T_486,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19191.4]
  assign _T_494 = {_T_487,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19193.4]
  assign _T_496 = {_T_488,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@19195.4]
  assign _T_497 = _T_487 ? _T_494 : _T_496; // @[Mux.scala 31:69:@19196.4]
  assign _T_498 = _T_486 ? _T_492 : _T_497; // @[Mux.scala 31:69:@19197.4]
  assign _T_499 = _T_485 ? _T_490 : _T_498; // @[Mux.scala 31:69:@19198.4]
  assign _T_506 = io_rPort_3_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@19206.4]
  assign _T_507 = _T_440 & _T_506; // @[MemPrimitives.scala 110:228:@19207.4]
  assign _T_512 = io_rPort_5_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@19210.4]
  assign _T_513 = _T_446 & _T_512; // @[MemPrimitives.scala 110:228:@19211.4]
  assign _T_515 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 126:35:@19218.4]
  assign _T_516 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 126:35:@19219.4]
  assign _T_518 = {_T_515,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19221.4]
  assign _T_520 = {_T_516,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@19223.4]
  assign _T_521 = _T_515 ? _T_518 : _T_520; // @[Mux.scala 31:69:@19224.4]
  assign _T_528 = io_rPort_0_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@19232.4]
  assign _T_529 = _T_462 & _T_528; // @[MemPrimitives.scala 110:228:@19233.4]
  assign _T_534 = io_rPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@19236.4]
  assign _T_535 = _T_468 & _T_534; // @[MemPrimitives.scala 110:228:@19237.4]
  assign _T_540 = io_rPort_2_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@19240.4]
  assign _T_541 = _T_474 & _T_540; // @[MemPrimitives.scala 110:228:@19241.4]
  assign _T_546 = io_rPort_4_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@19244.4]
  assign _T_547 = _T_480 & _T_546; // @[MemPrimitives.scala 110:228:@19245.4]
  assign _T_549 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 126:35:@19254.4]
  assign _T_550 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 126:35:@19255.4]
  assign _T_551 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 126:35:@19256.4]
  assign _T_552 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 126:35:@19257.4]
  assign _T_554 = {_T_549,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19259.4]
  assign _T_556 = {_T_550,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19261.4]
  assign _T_558 = {_T_551,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19263.4]
  assign _T_560 = {_T_552,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@19265.4]
  assign _T_561 = _T_551 ? _T_558 : _T_560; // @[Mux.scala 31:69:@19266.4]
  assign _T_562 = _T_550 ? _T_556 : _T_561; // @[Mux.scala 31:69:@19267.4]
  assign _T_563 = _T_549 ? _T_554 : _T_562; // @[Mux.scala 31:69:@19268.4]
  assign _T_568 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@19275.4]
  assign _T_571 = _T_568 & _T_442; // @[MemPrimitives.scala 110:228:@19277.4]
  assign _T_574 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@19279.4]
  assign _T_577 = _T_574 & _T_448; // @[MemPrimitives.scala 110:228:@19281.4]
  assign _T_579 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 126:35:@19288.4]
  assign _T_580 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 126:35:@19289.4]
  assign _T_582 = {_T_579,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19291.4]
  assign _T_584 = {_T_580,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@19293.4]
  assign _T_585 = _T_579 ? _T_582 : _T_584; // @[Mux.scala 31:69:@19294.4]
  assign _T_590 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@19301.4]
  assign _T_593 = _T_590 & _T_464; // @[MemPrimitives.scala 110:228:@19303.4]
  assign _T_596 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@19305.4]
  assign _T_599 = _T_596 & _T_470; // @[MemPrimitives.scala 110:228:@19307.4]
  assign _T_602 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@19309.4]
  assign _T_605 = _T_602 & _T_476; // @[MemPrimitives.scala 110:228:@19311.4]
  assign _T_608 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@19313.4]
  assign _T_611 = _T_608 & _T_482; // @[MemPrimitives.scala 110:228:@19315.4]
  assign _T_613 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 126:35:@19324.4]
  assign _T_614 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 126:35:@19325.4]
  assign _T_615 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 126:35:@19326.4]
  assign _T_616 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 126:35:@19327.4]
  assign _T_618 = {_T_613,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19329.4]
  assign _T_620 = {_T_614,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19331.4]
  assign _T_622 = {_T_615,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19333.4]
  assign _T_624 = {_T_616,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@19335.4]
  assign _T_625 = _T_615 ? _T_622 : _T_624; // @[Mux.scala 31:69:@19336.4]
  assign _T_626 = _T_614 ? _T_620 : _T_625; // @[Mux.scala 31:69:@19337.4]
  assign _T_627 = _T_613 ? _T_618 : _T_626; // @[Mux.scala 31:69:@19338.4]
  assign _T_635 = _T_568 & _T_506; // @[MemPrimitives.scala 110:228:@19347.4]
  assign _T_641 = _T_574 & _T_512; // @[MemPrimitives.scala 110:228:@19351.4]
  assign _T_643 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 126:35:@19358.4]
  assign _T_644 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 126:35:@19359.4]
  assign _T_646 = {_T_643,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19361.4]
  assign _T_648 = {_T_644,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@19363.4]
  assign _T_649 = _T_643 ? _T_646 : _T_648; // @[Mux.scala 31:69:@19364.4]
  assign _T_657 = _T_590 & _T_528; // @[MemPrimitives.scala 110:228:@19373.4]
  assign _T_663 = _T_596 & _T_534; // @[MemPrimitives.scala 110:228:@19377.4]
  assign _T_669 = _T_602 & _T_540; // @[MemPrimitives.scala 110:228:@19381.4]
  assign _T_675 = _T_608 & _T_546; // @[MemPrimitives.scala 110:228:@19385.4]
  assign _T_677 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 126:35:@19394.4]
  assign _T_678 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 126:35:@19395.4]
  assign _T_679 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 126:35:@19396.4]
  assign _T_680 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 126:35:@19397.4]
  assign _T_682 = {_T_677,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19399.4]
  assign _T_684 = {_T_678,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19401.4]
  assign _T_686 = {_T_679,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19403.4]
  assign _T_688 = {_T_680,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@19405.4]
  assign _T_689 = _T_679 ? _T_686 : _T_688; // @[Mux.scala 31:69:@19406.4]
  assign _T_690 = _T_678 ? _T_684 : _T_689; // @[Mux.scala 31:69:@19407.4]
  assign _T_691 = _T_677 ? _T_682 : _T_690; // @[Mux.scala 31:69:@19408.4]
  assign _T_696 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19415.4]
  assign _T_699 = _T_696 & _T_442; // @[MemPrimitives.scala 110:228:@19417.4]
  assign _T_702 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19419.4]
  assign _T_705 = _T_702 & _T_448; // @[MemPrimitives.scala 110:228:@19421.4]
  assign _T_707 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 126:35:@19428.4]
  assign _T_708 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 126:35:@19429.4]
  assign _T_710 = {_T_707,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19431.4]
  assign _T_712 = {_T_708,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@19433.4]
  assign _T_713 = _T_707 ? _T_710 : _T_712; // @[Mux.scala 31:69:@19434.4]
  assign _T_718 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19441.4]
  assign _T_721 = _T_718 & _T_464; // @[MemPrimitives.scala 110:228:@19443.4]
  assign _T_724 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19445.4]
  assign _T_727 = _T_724 & _T_470; // @[MemPrimitives.scala 110:228:@19447.4]
  assign _T_730 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19449.4]
  assign _T_733 = _T_730 & _T_476; // @[MemPrimitives.scala 110:228:@19451.4]
  assign _T_736 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@19453.4]
  assign _T_739 = _T_736 & _T_482; // @[MemPrimitives.scala 110:228:@19455.4]
  assign _T_741 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 126:35:@19464.4]
  assign _T_742 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 126:35:@19465.4]
  assign _T_743 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 126:35:@19466.4]
  assign _T_744 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 126:35:@19467.4]
  assign _T_746 = {_T_741,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19469.4]
  assign _T_748 = {_T_742,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19471.4]
  assign _T_750 = {_T_743,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19473.4]
  assign _T_752 = {_T_744,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@19475.4]
  assign _T_753 = _T_743 ? _T_750 : _T_752; // @[Mux.scala 31:69:@19476.4]
  assign _T_754 = _T_742 ? _T_748 : _T_753; // @[Mux.scala 31:69:@19477.4]
  assign _T_755 = _T_741 ? _T_746 : _T_754; // @[Mux.scala 31:69:@19478.4]
  assign _T_763 = _T_696 & _T_506; // @[MemPrimitives.scala 110:228:@19487.4]
  assign _T_769 = _T_702 & _T_512; // @[MemPrimitives.scala 110:228:@19491.4]
  assign _T_771 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 126:35:@19498.4]
  assign _T_772 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 126:35:@19499.4]
  assign _T_774 = {_T_771,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19501.4]
  assign _T_776 = {_T_772,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@19503.4]
  assign _T_777 = _T_771 ? _T_774 : _T_776; // @[Mux.scala 31:69:@19504.4]
  assign _T_785 = _T_718 & _T_528; // @[MemPrimitives.scala 110:228:@19513.4]
  assign _T_791 = _T_724 & _T_534; // @[MemPrimitives.scala 110:228:@19517.4]
  assign _T_797 = _T_730 & _T_540; // @[MemPrimitives.scala 110:228:@19521.4]
  assign _T_803 = _T_736 & _T_546; // @[MemPrimitives.scala 110:228:@19525.4]
  assign _T_805 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 126:35:@19534.4]
  assign _T_806 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 126:35:@19535.4]
  assign _T_807 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 126:35:@19536.4]
  assign _T_808 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 126:35:@19537.4]
  assign _T_810 = {_T_805,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19539.4]
  assign _T_812 = {_T_806,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19541.4]
  assign _T_814 = {_T_807,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19543.4]
  assign _T_816 = {_T_808,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@19545.4]
  assign _T_817 = _T_807 ? _T_814 : _T_816; // @[Mux.scala 31:69:@19546.4]
  assign _T_818 = _T_806 ? _T_812 : _T_817; // @[Mux.scala 31:69:@19547.4]
  assign _T_819 = _T_805 ? _T_810 : _T_818; // @[Mux.scala 31:69:@19548.4]
  assign _T_824 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19555.4]
  assign _T_827 = _T_824 & _T_442; // @[MemPrimitives.scala 110:228:@19557.4]
  assign _T_830 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19559.4]
  assign _T_833 = _T_830 & _T_448; // @[MemPrimitives.scala 110:228:@19561.4]
  assign _T_835 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 126:35:@19568.4]
  assign _T_836 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 126:35:@19569.4]
  assign _T_838 = {_T_835,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19571.4]
  assign _T_840 = {_T_836,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@19573.4]
  assign _T_841 = _T_835 ? _T_838 : _T_840; // @[Mux.scala 31:69:@19574.4]
  assign _T_846 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19581.4]
  assign _T_849 = _T_846 & _T_464; // @[MemPrimitives.scala 110:228:@19583.4]
  assign _T_852 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19585.4]
  assign _T_855 = _T_852 & _T_470; // @[MemPrimitives.scala 110:228:@19587.4]
  assign _T_858 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19589.4]
  assign _T_861 = _T_858 & _T_476; // @[MemPrimitives.scala 110:228:@19591.4]
  assign _T_864 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@19593.4]
  assign _T_867 = _T_864 & _T_482; // @[MemPrimitives.scala 110:228:@19595.4]
  assign _T_869 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 126:35:@19604.4]
  assign _T_870 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 126:35:@19605.4]
  assign _T_871 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 126:35:@19606.4]
  assign _T_872 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 126:35:@19607.4]
  assign _T_874 = {_T_869,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19609.4]
  assign _T_876 = {_T_870,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19611.4]
  assign _T_878 = {_T_871,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19613.4]
  assign _T_880 = {_T_872,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@19615.4]
  assign _T_881 = _T_871 ? _T_878 : _T_880; // @[Mux.scala 31:69:@19616.4]
  assign _T_882 = _T_870 ? _T_876 : _T_881; // @[Mux.scala 31:69:@19617.4]
  assign _T_883 = _T_869 ? _T_874 : _T_882; // @[Mux.scala 31:69:@19618.4]
  assign _T_891 = _T_824 & _T_506; // @[MemPrimitives.scala 110:228:@19627.4]
  assign _T_897 = _T_830 & _T_512; // @[MemPrimitives.scala 110:228:@19631.4]
  assign _T_899 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 126:35:@19638.4]
  assign _T_900 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 126:35:@19639.4]
  assign _T_902 = {_T_899,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@19641.4]
  assign _T_904 = {_T_900,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@19643.4]
  assign _T_905 = _T_899 ? _T_902 : _T_904; // @[Mux.scala 31:69:@19644.4]
  assign _T_913 = _T_846 & _T_528; // @[MemPrimitives.scala 110:228:@19653.4]
  assign _T_919 = _T_852 & _T_534; // @[MemPrimitives.scala 110:228:@19657.4]
  assign _T_925 = _T_858 & _T_540; // @[MemPrimitives.scala 110:228:@19661.4]
  assign _T_931 = _T_864 & _T_546; // @[MemPrimitives.scala 110:228:@19665.4]
  assign _T_933 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 126:35:@19674.4]
  assign _T_934 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 126:35:@19675.4]
  assign _T_935 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 126:35:@19676.4]
  assign _T_936 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 126:35:@19677.4]
  assign _T_938 = {_T_933,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@19679.4]
  assign _T_940 = {_T_934,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@19681.4]
  assign _T_942 = {_T_935,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@19683.4]
  assign _T_944 = {_T_936,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@19685.4]
  assign _T_945 = _T_935 ? _T_942 : _T_944; // @[Mux.scala 31:69:@19686.4]
  assign _T_946 = _T_934 ? _T_940 : _T_945; // @[Mux.scala 31:69:@19687.4]
  assign _T_947 = _T_933 ? _T_938 : _T_946; // @[Mux.scala 31:69:@19688.4]
  assign _T_1011 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@19773.4 package.scala 96:25:@19774.4]
  assign _T_1015 = _T_1011 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@19783.4]
  assign _T_1008 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@19765.4 package.scala 96:25:@19766.4]
  assign _T_1016 = _T_1008 ? Mem1D_11_io_output : _T_1015; // @[Mux.scala 31:69:@19784.4]
  assign _T_1005 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@19757.4 package.scala 96:25:@19758.4]
  assign _T_1017 = _T_1005 ? Mem1D_9_io_output : _T_1016; // @[Mux.scala 31:69:@19785.4]
  assign _T_1002 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@19749.4 package.scala 96:25:@19750.4]
  assign _T_1018 = _T_1002 ? Mem1D_7_io_output : _T_1017; // @[Mux.scala 31:69:@19786.4]
  assign _T_999 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@19741.4 package.scala 96:25:@19742.4]
  assign _T_1019 = _T_999 ? Mem1D_5_io_output : _T_1018; // @[Mux.scala 31:69:@19787.4]
  assign _T_996 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@19733.4 package.scala 96:25:@19734.4]
  assign _T_1020 = _T_996 ? Mem1D_3_io_output : _T_1019; // @[Mux.scala 31:69:@19788.4]
  assign _T_993 = RetimeWrapper_io_out; // @[package.scala 96:25:@19725.4 package.scala 96:25:@19726.4]
  assign _T_1082 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@19869.4 package.scala 96:25:@19870.4]
  assign _T_1086 = _T_1082 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@19879.4]
  assign _T_1079 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@19861.4 package.scala 96:25:@19862.4]
  assign _T_1087 = _T_1079 ? Mem1D_11_io_output : _T_1086; // @[Mux.scala 31:69:@19880.4]
  assign _T_1076 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@19853.4 package.scala 96:25:@19854.4]
  assign _T_1088 = _T_1076 ? Mem1D_9_io_output : _T_1087; // @[Mux.scala 31:69:@19881.4]
  assign _T_1073 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@19845.4 package.scala 96:25:@19846.4]
  assign _T_1089 = _T_1073 ? Mem1D_7_io_output : _T_1088; // @[Mux.scala 31:69:@19882.4]
  assign _T_1070 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@19837.4 package.scala 96:25:@19838.4]
  assign _T_1090 = _T_1070 ? Mem1D_5_io_output : _T_1089; // @[Mux.scala 31:69:@19883.4]
  assign _T_1067 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@19829.4 package.scala 96:25:@19830.4]
  assign _T_1091 = _T_1067 ? Mem1D_3_io_output : _T_1090; // @[Mux.scala 31:69:@19884.4]
  assign _T_1064 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@19821.4 package.scala 96:25:@19822.4]
  assign _T_1153 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@19965.4 package.scala 96:25:@19966.4]
  assign _T_1157 = _T_1153 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@19975.4]
  assign _T_1150 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@19957.4 package.scala 96:25:@19958.4]
  assign _T_1158 = _T_1150 ? Mem1D_11_io_output : _T_1157; // @[Mux.scala 31:69:@19976.4]
  assign _T_1147 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@19949.4 package.scala 96:25:@19950.4]
  assign _T_1159 = _T_1147 ? Mem1D_9_io_output : _T_1158; // @[Mux.scala 31:69:@19977.4]
  assign _T_1144 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@19941.4 package.scala 96:25:@19942.4]
  assign _T_1160 = _T_1144 ? Mem1D_7_io_output : _T_1159; // @[Mux.scala 31:69:@19978.4]
  assign _T_1141 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@19933.4 package.scala 96:25:@19934.4]
  assign _T_1161 = _T_1141 ? Mem1D_5_io_output : _T_1160; // @[Mux.scala 31:69:@19979.4]
  assign _T_1138 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@19925.4 package.scala 96:25:@19926.4]
  assign _T_1162 = _T_1138 ? Mem1D_3_io_output : _T_1161; // @[Mux.scala 31:69:@19980.4]
  assign _T_1135 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@19917.4 package.scala 96:25:@19918.4]
  assign _T_1224 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@20061.4 package.scala 96:25:@20062.4]
  assign _T_1228 = _T_1224 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@20071.4]
  assign _T_1221 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@20053.4 package.scala 96:25:@20054.4]
  assign _T_1229 = _T_1221 ? Mem1D_10_io_output : _T_1228; // @[Mux.scala 31:69:@20072.4]
  assign _T_1218 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@20045.4 package.scala 96:25:@20046.4]
  assign _T_1230 = _T_1218 ? Mem1D_8_io_output : _T_1229; // @[Mux.scala 31:69:@20073.4]
  assign _T_1215 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@20037.4 package.scala 96:25:@20038.4]
  assign _T_1231 = _T_1215 ? Mem1D_6_io_output : _T_1230; // @[Mux.scala 31:69:@20074.4]
  assign _T_1212 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@20029.4 package.scala 96:25:@20030.4]
  assign _T_1232 = _T_1212 ? Mem1D_4_io_output : _T_1231; // @[Mux.scala 31:69:@20075.4]
  assign _T_1209 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@20021.4 package.scala 96:25:@20022.4]
  assign _T_1233 = _T_1209 ? Mem1D_2_io_output : _T_1232; // @[Mux.scala 31:69:@20076.4]
  assign _T_1206 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@20013.4 package.scala 96:25:@20014.4]
  assign _T_1295 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@20157.4 package.scala 96:25:@20158.4]
  assign _T_1299 = _T_1295 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@20167.4]
  assign _T_1292 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@20149.4 package.scala 96:25:@20150.4]
  assign _T_1300 = _T_1292 ? Mem1D_11_io_output : _T_1299; // @[Mux.scala 31:69:@20168.4]
  assign _T_1289 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@20141.4 package.scala 96:25:@20142.4]
  assign _T_1301 = _T_1289 ? Mem1D_9_io_output : _T_1300; // @[Mux.scala 31:69:@20169.4]
  assign _T_1286 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@20133.4 package.scala 96:25:@20134.4]
  assign _T_1302 = _T_1286 ? Mem1D_7_io_output : _T_1301; // @[Mux.scala 31:69:@20170.4]
  assign _T_1283 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@20125.4 package.scala 96:25:@20126.4]
  assign _T_1303 = _T_1283 ? Mem1D_5_io_output : _T_1302; // @[Mux.scala 31:69:@20171.4]
  assign _T_1280 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@20117.4 package.scala 96:25:@20118.4]
  assign _T_1304 = _T_1280 ? Mem1D_3_io_output : _T_1303; // @[Mux.scala 31:69:@20172.4]
  assign _T_1277 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@20109.4 package.scala 96:25:@20110.4]
  assign _T_1366 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@20253.4 package.scala 96:25:@20254.4]
  assign _T_1370 = _T_1366 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@20263.4]
  assign _T_1363 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@20245.4 package.scala 96:25:@20246.4]
  assign _T_1371 = _T_1363 ? Mem1D_10_io_output : _T_1370; // @[Mux.scala 31:69:@20264.4]
  assign _T_1360 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@20237.4 package.scala 96:25:@20238.4]
  assign _T_1372 = _T_1360 ? Mem1D_8_io_output : _T_1371; // @[Mux.scala 31:69:@20265.4]
  assign _T_1357 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@20229.4 package.scala 96:25:@20230.4]
  assign _T_1373 = _T_1357 ? Mem1D_6_io_output : _T_1372; // @[Mux.scala 31:69:@20266.4]
  assign _T_1354 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@20221.4 package.scala 96:25:@20222.4]
  assign _T_1374 = _T_1354 ? Mem1D_4_io_output : _T_1373; // @[Mux.scala 31:69:@20267.4]
  assign _T_1351 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@20213.4 package.scala 96:25:@20214.4]
  assign _T_1375 = _T_1351 ? Mem1D_2_io_output : _T_1374; // @[Mux.scala 31:69:@20268.4]
  assign _T_1348 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@20205.4 package.scala 96:25:@20206.4]
  assign io_rPort_5_output_0 = _T_1348 ? Mem1D_io_output : _T_1375; // @[MemPrimitives.scala 152:13:@20270.4]
  assign io_rPort_4_output_0 = _T_1277 ? Mem1D_1_io_output : _T_1304; // @[MemPrimitives.scala 152:13:@20174.4]
  assign io_rPort_3_output_0 = _T_1206 ? Mem1D_io_output : _T_1233; // @[MemPrimitives.scala 152:13:@20078.4]
  assign io_rPort_2_output_0 = _T_1135 ? Mem1D_1_io_output : _T_1162; // @[MemPrimitives.scala 152:13:@19982.4]
  assign io_rPort_1_output_0 = _T_1064 ? Mem1D_1_io_output : _T_1091; // @[MemPrimitives.scala 152:13:@19886.4]
  assign io_rPort_0_output_0 = _T_993 ? Mem1D_1_io_output : _T_1020; // @[MemPrimitives.scala 152:13:@19790.4]
  assign Mem1D_clock = clock; // @[:@18688.4]
  assign Mem1D_reset = reset; // @[:@18689.4]
  assign Mem1D_io_r_ofs_0 = _T_457[8:0]; // @[MemPrimitives.scala 131:28:@19158.4]
  assign Mem1D_io_r_backpressure = _T_457[9]; // @[MemPrimitives.scala 132:32:@19159.4]
  assign Mem1D_io_w_ofs_0 = _T_270[8:0]; // @[MemPrimitives.scala 94:28:@18952.4]
  assign Mem1D_io_w_data_0 = _T_270[40:9]; // @[MemPrimitives.scala 95:29:@18953.4]
  assign Mem1D_io_w_en_0 = _T_270[41]; // @[MemPrimitives.scala 96:27:@18954.4]
  assign Mem1D_1_clock = clock; // @[:@18704.4]
  assign Mem1D_1_reset = reset; // @[:@18705.4]
  assign Mem1D_1_io_r_ofs_0 = _T_499[8:0]; // @[MemPrimitives.scala 131:28:@19202.4]
  assign Mem1D_1_io_r_backpressure = _T_499[9]; // @[MemPrimitives.scala 132:32:@19203.4]
  assign Mem1D_1_io_w_ofs_0 = _T_281[8:0]; // @[MemPrimitives.scala 94:28:@18964.4]
  assign Mem1D_1_io_w_data_0 = _T_281[40:9]; // @[MemPrimitives.scala 95:29:@18965.4]
  assign Mem1D_1_io_w_en_0 = _T_281[41]; // @[MemPrimitives.scala 96:27:@18966.4]
  assign Mem1D_2_clock = clock; // @[:@18720.4]
  assign Mem1D_2_reset = reset; // @[:@18721.4]
  assign Mem1D_2_io_r_ofs_0 = _T_521[8:0]; // @[MemPrimitives.scala 131:28:@19228.4]
  assign Mem1D_2_io_r_backpressure = _T_521[9]; // @[MemPrimitives.scala 132:32:@19229.4]
  assign Mem1D_2_io_w_ofs_0 = _T_292[8:0]; // @[MemPrimitives.scala 94:28:@18976.4]
  assign Mem1D_2_io_w_data_0 = _T_292[40:9]; // @[MemPrimitives.scala 95:29:@18977.4]
  assign Mem1D_2_io_w_en_0 = _T_292[41]; // @[MemPrimitives.scala 96:27:@18978.4]
  assign Mem1D_3_clock = clock; // @[:@18736.4]
  assign Mem1D_3_reset = reset; // @[:@18737.4]
  assign Mem1D_3_io_r_ofs_0 = _T_563[8:0]; // @[MemPrimitives.scala 131:28:@19272.4]
  assign Mem1D_3_io_r_backpressure = _T_563[9]; // @[MemPrimitives.scala 132:32:@19273.4]
  assign Mem1D_3_io_w_ofs_0 = _T_303[8:0]; // @[MemPrimitives.scala 94:28:@18988.4]
  assign Mem1D_3_io_w_data_0 = _T_303[40:9]; // @[MemPrimitives.scala 95:29:@18989.4]
  assign Mem1D_3_io_w_en_0 = _T_303[41]; // @[MemPrimitives.scala 96:27:@18990.4]
  assign Mem1D_4_clock = clock; // @[:@18752.4]
  assign Mem1D_4_reset = reset; // @[:@18753.4]
  assign Mem1D_4_io_r_ofs_0 = _T_585[8:0]; // @[MemPrimitives.scala 131:28:@19298.4]
  assign Mem1D_4_io_r_backpressure = _T_585[9]; // @[MemPrimitives.scala 132:32:@19299.4]
  assign Mem1D_4_io_w_ofs_0 = _T_314[8:0]; // @[MemPrimitives.scala 94:28:@19000.4]
  assign Mem1D_4_io_w_data_0 = _T_314[40:9]; // @[MemPrimitives.scala 95:29:@19001.4]
  assign Mem1D_4_io_w_en_0 = _T_314[41]; // @[MemPrimitives.scala 96:27:@19002.4]
  assign Mem1D_5_clock = clock; // @[:@18768.4]
  assign Mem1D_5_reset = reset; // @[:@18769.4]
  assign Mem1D_5_io_r_ofs_0 = _T_627[8:0]; // @[MemPrimitives.scala 131:28:@19342.4]
  assign Mem1D_5_io_r_backpressure = _T_627[9]; // @[MemPrimitives.scala 132:32:@19343.4]
  assign Mem1D_5_io_w_ofs_0 = _T_325[8:0]; // @[MemPrimitives.scala 94:28:@19012.4]
  assign Mem1D_5_io_w_data_0 = _T_325[40:9]; // @[MemPrimitives.scala 95:29:@19013.4]
  assign Mem1D_5_io_w_en_0 = _T_325[41]; // @[MemPrimitives.scala 96:27:@19014.4]
  assign Mem1D_6_clock = clock; // @[:@18784.4]
  assign Mem1D_6_reset = reset; // @[:@18785.4]
  assign Mem1D_6_io_r_ofs_0 = _T_649[8:0]; // @[MemPrimitives.scala 131:28:@19368.4]
  assign Mem1D_6_io_r_backpressure = _T_649[9]; // @[MemPrimitives.scala 132:32:@19369.4]
  assign Mem1D_6_io_w_ofs_0 = _T_336[8:0]; // @[MemPrimitives.scala 94:28:@19024.4]
  assign Mem1D_6_io_w_data_0 = _T_336[40:9]; // @[MemPrimitives.scala 95:29:@19025.4]
  assign Mem1D_6_io_w_en_0 = _T_336[41]; // @[MemPrimitives.scala 96:27:@19026.4]
  assign Mem1D_7_clock = clock; // @[:@18800.4]
  assign Mem1D_7_reset = reset; // @[:@18801.4]
  assign Mem1D_7_io_r_ofs_0 = _T_691[8:0]; // @[MemPrimitives.scala 131:28:@19412.4]
  assign Mem1D_7_io_r_backpressure = _T_691[9]; // @[MemPrimitives.scala 132:32:@19413.4]
  assign Mem1D_7_io_w_ofs_0 = _T_347[8:0]; // @[MemPrimitives.scala 94:28:@19036.4]
  assign Mem1D_7_io_w_data_0 = _T_347[40:9]; // @[MemPrimitives.scala 95:29:@19037.4]
  assign Mem1D_7_io_w_en_0 = _T_347[41]; // @[MemPrimitives.scala 96:27:@19038.4]
  assign Mem1D_8_clock = clock; // @[:@18816.4]
  assign Mem1D_8_reset = reset; // @[:@18817.4]
  assign Mem1D_8_io_r_ofs_0 = _T_713[8:0]; // @[MemPrimitives.scala 131:28:@19438.4]
  assign Mem1D_8_io_r_backpressure = _T_713[9]; // @[MemPrimitives.scala 132:32:@19439.4]
  assign Mem1D_8_io_w_ofs_0 = _T_358[8:0]; // @[MemPrimitives.scala 94:28:@19048.4]
  assign Mem1D_8_io_w_data_0 = _T_358[40:9]; // @[MemPrimitives.scala 95:29:@19049.4]
  assign Mem1D_8_io_w_en_0 = _T_358[41]; // @[MemPrimitives.scala 96:27:@19050.4]
  assign Mem1D_9_clock = clock; // @[:@18832.4]
  assign Mem1D_9_reset = reset; // @[:@18833.4]
  assign Mem1D_9_io_r_ofs_0 = _T_755[8:0]; // @[MemPrimitives.scala 131:28:@19482.4]
  assign Mem1D_9_io_r_backpressure = _T_755[9]; // @[MemPrimitives.scala 132:32:@19483.4]
  assign Mem1D_9_io_w_ofs_0 = _T_369[8:0]; // @[MemPrimitives.scala 94:28:@19060.4]
  assign Mem1D_9_io_w_data_0 = _T_369[40:9]; // @[MemPrimitives.scala 95:29:@19061.4]
  assign Mem1D_9_io_w_en_0 = _T_369[41]; // @[MemPrimitives.scala 96:27:@19062.4]
  assign Mem1D_10_clock = clock; // @[:@18848.4]
  assign Mem1D_10_reset = reset; // @[:@18849.4]
  assign Mem1D_10_io_r_ofs_0 = _T_777[8:0]; // @[MemPrimitives.scala 131:28:@19508.4]
  assign Mem1D_10_io_r_backpressure = _T_777[9]; // @[MemPrimitives.scala 132:32:@19509.4]
  assign Mem1D_10_io_w_ofs_0 = _T_380[8:0]; // @[MemPrimitives.scala 94:28:@19072.4]
  assign Mem1D_10_io_w_data_0 = _T_380[40:9]; // @[MemPrimitives.scala 95:29:@19073.4]
  assign Mem1D_10_io_w_en_0 = _T_380[41]; // @[MemPrimitives.scala 96:27:@19074.4]
  assign Mem1D_11_clock = clock; // @[:@18864.4]
  assign Mem1D_11_reset = reset; // @[:@18865.4]
  assign Mem1D_11_io_r_ofs_0 = _T_819[8:0]; // @[MemPrimitives.scala 131:28:@19552.4]
  assign Mem1D_11_io_r_backpressure = _T_819[9]; // @[MemPrimitives.scala 132:32:@19553.4]
  assign Mem1D_11_io_w_ofs_0 = _T_391[8:0]; // @[MemPrimitives.scala 94:28:@19084.4]
  assign Mem1D_11_io_w_data_0 = _T_391[40:9]; // @[MemPrimitives.scala 95:29:@19085.4]
  assign Mem1D_11_io_w_en_0 = _T_391[41]; // @[MemPrimitives.scala 96:27:@19086.4]
  assign Mem1D_12_clock = clock; // @[:@18880.4]
  assign Mem1D_12_reset = reset; // @[:@18881.4]
  assign Mem1D_12_io_r_ofs_0 = _T_841[8:0]; // @[MemPrimitives.scala 131:28:@19578.4]
  assign Mem1D_12_io_r_backpressure = _T_841[9]; // @[MemPrimitives.scala 132:32:@19579.4]
  assign Mem1D_12_io_w_ofs_0 = _T_402[8:0]; // @[MemPrimitives.scala 94:28:@19096.4]
  assign Mem1D_12_io_w_data_0 = _T_402[40:9]; // @[MemPrimitives.scala 95:29:@19097.4]
  assign Mem1D_12_io_w_en_0 = _T_402[41]; // @[MemPrimitives.scala 96:27:@19098.4]
  assign Mem1D_13_clock = clock; // @[:@18896.4]
  assign Mem1D_13_reset = reset; // @[:@18897.4]
  assign Mem1D_13_io_r_ofs_0 = _T_883[8:0]; // @[MemPrimitives.scala 131:28:@19622.4]
  assign Mem1D_13_io_r_backpressure = _T_883[9]; // @[MemPrimitives.scala 132:32:@19623.4]
  assign Mem1D_13_io_w_ofs_0 = _T_413[8:0]; // @[MemPrimitives.scala 94:28:@19108.4]
  assign Mem1D_13_io_w_data_0 = _T_413[40:9]; // @[MemPrimitives.scala 95:29:@19109.4]
  assign Mem1D_13_io_w_en_0 = _T_413[41]; // @[MemPrimitives.scala 96:27:@19110.4]
  assign Mem1D_14_clock = clock; // @[:@18912.4]
  assign Mem1D_14_reset = reset; // @[:@18913.4]
  assign Mem1D_14_io_r_ofs_0 = _T_905[8:0]; // @[MemPrimitives.scala 131:28:@19648.4]
  assign Mem1D_14_io_r_backpressure = _T_905[9]; // @[MemPrimitives.scala 132:32:@19649.4]
  assign Mem1D_14_io_w_ofs_0 = _T_424[8:0]; // @[MemPrimitives.scala 94:28:@19120.4]
  assign Mem1D_14_io_w_data_0 = _T_424[40:9]; // @[MemPrimitives.scala 95:29:@19121.4]
  assign Mem1D_14_io_w_en_0 = _T_424[41]; // @[MemPrimitives.scala 96:27:@19122.4]
  assign Mem1D_15_clock = clock; // @[:@18928.4]
  assign Mem1D_15_reset = reset; // @[:@18929.4]
  assign Mem1D_15_io_r_ofs_0 = _T_947[8:0]; // @[MemPrimitives.scala 131:28:@19692.4]
  assign Mem1D_15_io_r_backpressure = _T_947[9]; // @[MemPrimitives.scala 132:32:@19693.4]
  assign Mem1D_15_io_w_ofs_0 = _T_435[8:0]; // @[MemPrimitives.scala 94:28:@19132.4]
  assign Mem1D_15_io_w_data_0 = _T_435[40:9]; // @[MemPrimitives.scala 95:29:@19133.4]
  assign Mem1D_15_io_w_en_0 = _T_435[41]; // @[MemPrimitives.scala 96:27:@19134.4]
  assign StickySelects_clock = clock; // @[:@19144.4]
  assign StickySelects_reset = reset; // @[:@19145.4]
  assign StickySelects_io_ins_0 = io_rPort_3_en_0 & _T_443; // @[MemPrimitives.scala 125:64:@19146.4]
  assign StickySelects_io_ins_1 = io_rPort_5_en_0 & _T_449; // @[MemPrimitives.scala 125:64:@19147.4]
  assign StickySelects_1_clock = clock; // @[:@19178.4]
  assign StickySelects_1_reset = reset; // @[:@19179.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_465; // @[MemPrimitives.scala 125:64:@19180.4]
  assign StickySelects_1_io_ins_1 = io_rPort_1_en_0 & _T_471; // @[MemPrimitives.scala 125:64:@19181.4]
  assign StickySelects_1_io_ins_2 = io_rPort_2_en_0 & _T_477; // @[MemPrimitives.scala 125:64:@19182.4]
  assign StickySelects_1_io_ins_3 = io_rPort_4_en_0 & _T_483; // @[MemPrimitives.scala 125:64:@19183.4]
  assign StickySelects_2_clock = clock; // @[:@19214.4]
  assign StickySelects_2_reset = reset; // @[:@19215.4]
  assign StickySelects_2_io_ins_0 = io_rPort_3_en_0 & _T_507; // @[MemPrimitives.scala 125:64:@19216.4]
  assign StickySelects_2_io_ins_1 = io_rPort_5_en_0 & _T_513; // @[MemPrimitives.scala 125:64:@19217.4]
  assign StickySelects_3_clock = clock; // @[:@19248.4]
  assign StickySelects_3_reset = reset; // @[:@19249.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_529; // @[MemPrimitives.scala 125:64:@19250.4]
  assign StickySelects_3_io_ins_1 = io_rPort_1_en_0 & _T_535; // @[MemPrimitives.scala 125:64:@19251.4]
  assign StickySelects_3_io_ins_2 = io_rPort_2_en_0 & _T_541; // @[MemPrimitives.scala 125:64:@19252.4]
  assign StickySelects_3_io_ins_3 = io_rPort_4_en_0 & _T_547; // @[MemPrimitives.scala 125:64:@19253.4]
  assign StickySelects_4_clock = clock; // @[:@19284.4]
  assign StickySelects_4_reset = reset; // @[:@19285.4]
  assign StickySelects_4_io_ins_0 = io_rPort_3_en_0 & _T_571; // @[MemPrimitives.scala 125:64:@19286.4]
  assign StickySelects_4_io_ins_1 = io_rPort_5_en_0 & _T_577; // @[MemPrimitives.scala 125:64:@19287.4]
  assign StickySelects_5_clock = clock; // @[:@19318.4]
  assign StickySelects_5_reset = reset; // @[:@19319.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_593; // @[MemPrimitives.scala 125:64:@19320.4]
  assign StickySelects_5_io_ins_1 = io_rPort_1_en_0 & _T_599; // @[MemPrimitives.scala 125:64:@19321.4]
  assign StickySelects_5_io_ins_2 = io_rPort_2_en_0 & _T_605; // @[MemPrimitives.scala 125:64:@19322.4]
  assign StickySelects_5_io_ins_3 = io_rPort_4_en_0 & _T_611; // @[MemPrimitives.scala 125:64:@19323.4]
  assign StickySelects_6_clock = clock; // @[:@19354.4]
  assign StickySelects_6_reset = reset; // @[:@19355.4]
  assign StickySelects_6_io_ins_0 = io_rPort_3_en_0 & _T_635; // @[MemPrimitives.scala 125:64:@19356.4]
  assign StickySelects_6_io_ins_1 = io_rPort_5_en_0 & _T_641; // @[MemPrimitives.scala 125:64:@19357.4]
  assign StickySelects_7_clock = clock; // @[:@19388.4]
  assign StickySelects_7_reset = reset; // @[:@19389.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_657; // @[MemPrimitives.scala 125:64:@19390.4]
  assign StickySelects_7_io_ins_1 = io_rPort_1_en_0 & _T_663; // @[MemPrimitives.scala 125:64:@19391.4]
  assign StickySelects_7_io_ins_2 = io_rPort_2_en_0 & _T_669; // @[MemPrimitives.scala 125:64:@19392.4]
  assign StickySelects_7_io_ins_3 = io_rPort_4_en_0 & _T_675; // @[MemPrimitives.scala 125:64:@19393.4]
  assign StickySelects_8_clock = clock; // @[:@19424.4]
  assign StickySelects_8_reset = reset; // @[:@19425.4]
  assign StickySelects_8_io_ins_0 = io_rPort_3_en_0 & _T_699; // @[MemPrimitives.scala 125:64:@19426.4]
  assign StickySelects_8_io_ins_1 = io_rPort_5_en_0 & _T_705; // @[MemPrimitives.scala 125:64:@19427.4]
  assign StickySelects_9_clock = clock; // @[:@19458.4]
  assign StickySelects_9_reset = reset; // @[:@19459.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_721; // @[MemPrimitives.scala 125:64:@19460.4]
  assign StickySelects_9_io_ins_1 = io_rPort_1_en_0 & _T_727; // @[MemPrimitives.scala 125:64:@19461.4]
  assign StickySelects_9_io_ins_2 = io_rPort_2_en_0 & _T_733; // @[MemPrimitives.scala 125:64:@19462.4]
  assign StickySelects_9_io_ins_3 = io_rPort_4_en_0 & _T_739; // @[MemPrimitives.scala 125:64:@19463.4]
  assign StickySelects_10_clock = clock; // @[:@19494.4]
  assign StickySelects_10_reset = reset; // @[:@19495.4]
  assign StickySelects_10_io_ins_0 = io_rPort_3_en_0 & _T_763; // @[MemPrimitives.scala 125:64:@19496.4]
  assign StickySelects_10_io_ins_1 = io_rPort_5_en_0 & _T_769; // @[MemPrimitives.scala 125:64:@19497.4]
  assign StickySelects_11_clock = clock; // @[:@19528.4]
  assign StickySelects_11_reset = reset; // @[:@19529.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_785; // @[MemPrimitives.scala 125:64:@19530.4]
  assign StickySelects_11_io_ins_1 = io_rPort_1_en_0 & _T_791; // @[MemPrimitives.scala 125:64:@19531.4]
  assign StickySelects_11_io_ins_2 = io_rPort_2_en_0 & _T_797; // @[MemPrimitives.scala 125:64:@19532.4]
  assign StickySelects_11_io_ins_3 = io_rPort_4_en_0 & _T_803; // @[MemPrimitives.scala 125:64:@19533.4]
  assign StickySelects_12_clock = clock; // @[:@19564.4]
  assign StickySelects_12_reset = reset; // @[:@19565.4]
  assign StickySelects_12_io_ins_0 = io_rPort_3_en_0 & _T_827; // @[MemPrimitives.scala 125:64:@19566.4]
  assign StickySelects_12_io_ins_1 = io_rPort_5_en_0 & _T_833; // @[MemPrimitives.scala 125:64:@19567.4]
  assign StickySelects_13_clock = clock; // @[:@19598.4]
  assign StickySelects_13_reset = reset; // @[:@19599.4]
  assign StickySelects_13_io_ins_0 = io_rPort_0_en_0 & _T_849; // @[MemPrimitives.scala 125:64:@19600.4]
  assign StickySelects_13_io_ins_1 = io_rPort_1_en_0 & _T_855; // @[MemPrimitives.scala 125:64:@19601.4]
  assign StickySelects_13_io_ins_2 = io_rPort_2_en_0 & _T_861; // @[MemPrimitives.scala 125:64:@19602.4]
  assign StickySelects_13_io_ins_3 = io_rPort_4_en_0 & _T_867; // @[MemPrimitives.scala 125:64:@19603.4]
  assign StickySelects_14_clock = clock; // @[:@19634.4]
  assign StickySelects_14_reset = reset; // @[:@19635.4]
  assign StickySelects_14_io_ins_0 = io_rPort_3_en_0 & _T_891; // @[MemPrimitives.scala 125:64:@19636.4]
  assign StickySelects_14_io_ins_1 = io_rPort_5_en_0 & _T_897; // @[MemPrimitives.scala 125:64:@19637.4]
  assign StickySelects_15_clock = clock; // @[:@19668.4]
  assign StickySelects_15_reset = reset; // @[:@19669.4]
  assign StickySelects_15_io_ins_0 = io_rPort_0_en_0 & _T_913; // @[MemPrimitives.scala 125:64:@19670.4]
  assign StickySelects_15_io_ins_1 = io_rPort_1_en_0 & _T_919; // @[MemPrimitives.scala 125:64:@19671.4]
  assign StickySelects_15_io_ins_2 = io_rPort_2_en_0 & _T_925; // @[MemPrimitives.scala 125:64:@19672.4]
  assign StickySelects_15_io_ins_3 = io_rPort_4_en_0 & _T_931; // @[MemPrimitives.scala 125:64:@19673.4]
  assign RetimeWrapper_clock = clock; // @[:@19721.4]
  assign RetimeWrapper_reset = reset; // @[:@19722.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19724.4]
  assign RetimeWrapper_io_in = _T_465 & io_rPort_0_en_0; // @[package.scala 94:16:@19723.4]
  assign RetimeWrapper_1_clock = clock; // @[:@19729.4]
  assign RetimeWrapper_1_reset = reset; // @[:@19730.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19732.4]
  assign RetimeWrapper_1_io_in = _T_529 & io_rPort_0_en_0; // @[package.scala 94:16:@19731.4]
  assign RetimeWrapper_2_clock = clock; // @[:@19737.4]
  assign RetimeWrapper_2_reset = reset; // @[:@19738.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19740.4]
  assign RetimeWrapper_2_io_in = _T_593 & io_rPort_0_en_0; // @[package.scala 94:16:@19739.4]
  assign RetimeWrapper_3_clock = clock; // @[:@19745.4]
  assign RetimeWrapper_3_reset = reset; // @[:@19746.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19748.4]
  assign RetimeWrapper_3_io_in = _T_657 & io_rPort_0_en_0; // @[package.scala 94:16:@19747.4]
  assign RetimeWrapper_4_clock = clock; // @[:@19753.4]
  assign RetimeWrapper_4_reset = reset; // @[:@19754.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19756.4]
  assign RetimeWrapper_4_io_in = _T_721 & io_rPort_0_en_0; // @[package.scala 94:16:@19755.4]
  assign RetimeWrapper_5_clock = clock; // @[:@19761.4]
  assign RetimeWrapper_5_reset = reset; // @[:@19762.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19764.4]
  assign RetimeWrapper_5_io_in = _T_785 & io_rPort_0_en_0; // @[package.scala 94:16:@19763.4]
  assign RetimeWrapper_6_clock = clock; // @[:@19769.4]
  assign RetimeWrapper_6_reset = reset; // @[:@19770.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19772.4]
  assign RetimeWrapper_6_io_in = _T_849 & io_rPort_0_en_0; // @[package.scala 94:16:@19771.4]
  assign RetimeWrapper_7_clock = clock; // @[:@19777.4]
  assign RetimeWrapper_7_reset = reset; // @[:@19778.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@19780.4]
  assign RetimeWrapper_7_io_in = _T_913 & io_rPort_0_en_0; // @[package.scala 94:16:@19779.4]
  assign RetimeWrapper_8_clock = clock; // @[:@19817.4]
  assign RetimeWrapper_8_reset = reset; // @[:@19818.4]
  assign RetimeWrapper_8_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19820.4]
  assign RetimeWrapper_8_io_in = _T_471 & io_rPort_1_en_0; // @[package.scala 94:16:@19819.4]
  assign RetimeWrapper_9_clock = clock; // @[:@19825.4]
  assign RetimeWrapper_9_reset = reset; // @[:@19826.4]
  assign RetimeWrapper_9_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19828.4]
  assign RetimeWrapper_9_io_in = _T_535 & io_rPort_1_en_0; // @[package.scala 94:16:@19827.4]
  assign RetimeWrapper_10_clock = clock; // @[:@19833.4]
  assign RetimeWrapper_10_reset = reset; // @[:@19834.4]
  assign RetimeWrapper_10_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19836.4]
  assign RetimeWrapper_10_io_in = _T_599 & io_rPort_1_en_0; // @[package.scala 94:16:@19835.4]
  assign RetimeWrapper_11_clock = clock; // @[:@19841.4]
  assign RetimeWrapper_11_reset = reset; // @[:@19842.4]
  assign RetimeWrapper_11_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19844.4]
  assign RetimeWrapper_11_io_in = _T_663 & io_rPort_1_en_0; // @[package.scala 94:16:@19843.4]
  assign RetimeWrapper_12_clock = clock; // @[:@19849.4]
  assign RetimeWrapper_12_reset = reset; // @[:@19850.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19852.4]
  assign RetimeWrapper_12_io_in = _T_727 & io_rPort_1_en_0; // @[package.scala 94:16:@19851.4]
  assign RetimeWrapper_13_clock = clock; // @[:@19857.4]
  assign RetimeWrapper_13_reset = reset; // @[:@19858.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19860.4]
  assign RetimeWrapper_13_io_in = _T_791 & io_rPort_1_en_0; // @[package.scala 94:16:@19859.4]
  assign RetimeWrapper_14_clock = clock; // @[:@19865.4]
  assign RetimeWrapper_14_reset = reset; // @[:@19866.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19868.4]
  assign RetimeWrapper_14_io_in = _T_855 & io_rPort_1_en_0; // @[package.scala 94:16:@19867.4]
  assign RetimeWrapper_15_clock = clock; // @[:@19873.4]
  assign RetimeWrapper_15_reset = reset; // @[:@19874.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@19876.4]
  assign RetimeWrapper_15_io_in = _T_919 & io_rPort_1_en_0; // @[package.scala 94:16:@19875.4]
  assign RetimeWrapper_16_clock = clock; // @[:@19913.4]
  assign RetimeWrapper_16_reset = reset; // @[:@19914.4]
  assign RetimeWrapper_16_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19916.4]
  assign RetimeWrapper_16_io_in = _T_477 & io_rPort_2_en_0; // @[package.scala 94:16:@19915.4]
  assign RetimeWrapper_17_clock = clock; // @[:@19921.4]
  assign RetimeWrapper_17_reset = reset; // @[:@19922.4]
  assign RetimeWrapper_17_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19924.4]
  assign RetimeWrapper_17_io_in = _T_541 & io_rPort_2_en_0; // @[package.scala 94:16:@19923.4]
  assign RetimeWrapper_18_clock = clock; // @[:@19929.4]
  assign RetimeWrapper_18_reset = reset; // @[:@19930.4]
  assign RetimeWrapper_18_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19932.4]
  assign RetimeWrapper_18_io_in = _T_605 & io_rPort_2_en_0; // @[package.scala 94:16:@19931.4]
  assign RetimeWrapper_19_clock = clock; // @[:@19937.4]
  assign RetimeWrapper_19_reset = reset; // @[:@19938.4]
  assign RetimeWrapper_19_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19940.4]
  assign RetimeWrapper_19_io_in = _T_669 & io_rPort_2_en_0; // @[package.scala 94:16:@19939.4]
  assign RetimeWrapper_20_clock = clock; // @[:@19945.4]
  assign RetimeWrapper_20_reset = reset; // @[:@19946.4]
  assign RetimeWrapper_20_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19948.4]
  assign RetimeWrapper_20_io_in = _T_733 & io_rPort_2_en_0; // @[package.scala 94:16:@19947.4]
  assign RetimeWrapper_21_clock = clock; // @[:@19953.4]
  assign RetimeWrapper_21_reset = reset; // @[:@19954.4]
  assign RetimeWrapper_21_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19956.4]
  assign RetimeWrapper_21_io_in = _T_797 & io_rPort_2_en_0; // @[package.scala 94:16:@19955.4]
  assign RetimeWrapper_22_clock = clock; // @[:@19961.4]
  assign RetimeWrapper_22_reset = reset; // @[:@19962.4]
  assign RetimeWrapper_22_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19964.4]
  assign RetimeWrapper_22_io_in = _T_861 & io_rPort_2_en_0; // @[package.scala 94:16:@19963.4]
  assign RetimeWrapper_23_clock = clock; // @[:@19969.4]
  assign RetimeWrapper_23_reset = reset; // @[:@19970.4]
  assign RetimeWrapper_23_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@19972.4]
  assign RetimeWrapper_23_io_in = _T_925 & io_rPort_2_en_0; // @[package.scala 94:16:@19971.4]
  assign RetimeWrapper_24_clock = clock; // @[:@20009.4]
  assign RetimeWrapper_24_reset = reset; // @[:@20010.4]
  assign RetimeWrapper_24_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@20012.4]
  assign RetimeWrapper_24_io_in = _T_443 & io_rPort_3_en_0; // @[package.scala 94:16:@20011.4]
  assign RetimeWrapper_25_clock = clock; // @[:@20017.4]
  assign RetimeWrapper_25_reset = reset; // @[:@20018.4]
  assign RetimeWrapper_25_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@20020.4]
  assign RetimeWrapper_25_io_in = _T_507 & io_rPort_3_en_0; // @[package.scala 94:16:@20019.4]
  assign RetimeWrapper_26_clock = clock; // @[:@20025.4]
  assign RetimeWrapper_26_reset = reset; // @[:@20026.4]
  assign RetimeWrapper_26_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@20028.4]
  assign RetimeWrapper_26_io_in = _T_571 & io_rPort_3_en_0; // @[package.scala 94:16:@20027.4]
  assign RetimeWrapper_27_clock = clock; // @[:@20033.4]
  assign RetimeWrapper_27_reset = reset; // @[:@20034.4]
  assign RetimeWrapper_27_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@20036.4]
  assign RetimeWrapper_27_io_in = _T_635 & io_rPort_3_en_0; // @[package.scala 94:16:@20035.4]
  assign RetimeWrapper_28_clock = clock; // @[:@20041.4]
  assign RetimeWrapper_28_reset = reset; // @[:@20042.4]
  assign RetimeWrapper_28_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@20044.4]
  assign RetimeWrapper_28_io_in = _T_699 & io_rPort_3_en_0; // @[package.scala 94:16:@20043.4]
  assign RetimeWrapper_29_clock = clock; // @[:@20049.4]
  assign RetimeWrapper_29_reset = reset; // @[:@20050.4]
  assign RetimeWrapper_29_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@20052.4]
  assign RetimeWrapper_29_io_in = _T_763 & io_rPort_3_en_0; // @[package.scala 94:16:@20051.4]
  assign RetimeWrapper_30_clock = clock; // @[:@20057.4]
  assign RetimeWrapper_30_reset = reset; // @[:@20058.4]
  assign RetimeWrapper_30_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@20060.4]
  assign RetimeWrapper_30_io_in = _T_827 & io_rPort_3_en_0; // @[package.scala 94:16:@20059.4]
  assign RetimeWrapper_31_clock = clock; // @[:@20065.4]
  assign RetimeWrapper_31_reset = reset; // @[:@20066.4]
  assign RetimeWrapper_31_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@20068.4]
  assign RetimeWrapper_31_io_in = _T_891 & io_rPort_3_en_0; // @[package.scala 94:16:@20067.4]
  assign RetimeWrapper_32_clock = clock; // @[:@20105.4]
  assign RetimeWrapper_32_reset = reset; // @[:@20106.4]
  assign RetimeWrapper_32_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@20108.4]
  assign RetimeWrapper_32_io_in = _T_483 & io_rPort_4_en_0; // @[package.scala 94:16:@20107.4]
  assign RetimeWrapper_33_clock = clock; // @[:@20113.4]
  assign RetimeWrapper_33_reset = reset; // @[:@20114.4]
  assign RetimeWrapper_33_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@20116.4]
  assign RetimeWrapper_33_io_in = _T_547 & io_rPort_4_en_0; // @[package.scala 94:16:@20115.4]
  assign RetimeWrapper_34_clock = clock; // @[:@20121.4]
  assign RetimeWrapper_34_reset = reset; // @[:@20122.4]
  assign RetimeWrapper_34_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@20124.4]
  assign RetimeWrapper_34_io_in = _T_611 & io_rPort_4_en_0; // @[package.scala 94:16:@20123.4]
  assign RetimeWrapper_35_clock = clock; // @[:@20129.4]
  assign RetimeWrapper_35_reset = reset; // @[:@20130.4]
  assign RetimeWrapper_35_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@20132.4]
  assign RetimeWrapper_35_io_in = _T_675 & io_rPort_4_en_0; // @[package.scala 94:16:@20131.4]
  assign RetimeWrapper_36_clock = clock; // @[:@20137.4]
  assign RetimeWrapper_36_reset = reset; // @[:@20138.4]
  assign RetimeWrapper_36_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@20140.4]
  assign RetimeWrapper_36_io_in = _T_739 & io_rPort_4_en_0; // @[package.scala 94:16:@20139.4]
  assign RetimeWrapper_37_clock = clock; // @[:@20145.4]
  assign RetimeWrapper_37_reset = reset; // @[:@20146.4]
  assign RetimeWrapper_37_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@20148.4]
  assign RetimeWrapper_37_io_in = _T_803 & io_rPort_4_en_0; // @[package.scala 94:16:@20147.4]
  assign RetimeWrapper_38_clock = clock; // @[:@20153.4]
  assign RetimeWrapper_38_reset = reset; // @[:@20154.4]
  assign RetimeWrapper_38_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@20156.4]
  assign RetimeWrapper_38_io_in = _T_867 & io_rPort_4_en_0; // @[package.scala 94:16:@20155.4]
  assign RetimeWrapper_39_clock = clock; // @[:@20161.4]
  assign RetimeWrapper_39_reset = reset; // @[:@20162.4]
  assign RetimeWrapper_39_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@20164.4]
  assign RetimeWrapper_39_io_in = _T_931 & io_rPort_4_en_0; // @[package.scala 94:16:@20163.4]
  assign RetimeWrapper_40_clock = clock; // @[:@20201.4]
  assign RetimeWrapper_40_reset = reset; // @[:@20202.4]
  assign RetimeWrapper_40_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@20204.4]
  assign RetimeWrapper_40_io_in = _T_449 & io_rPort_5_en_0; // @[package.scala 94:16:@20203.4]
  assign RetimeWrapper_41_clock = clock; // @[:@20209.4]
  assign RetimeWrapper_41_reset = reset; // @[:@20210.4]
  assign RetimeWrapper_41_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@20212.4]
  assign RetimeWrapper_41_io_in = _T_513 & io_rPort_5_en_0; // @[package.scala 94:16:@20211.4]
  assign RetimeWrapper_42_clock = clock; // @[:@20217.4]
  assign RetimeWrapper_42_reset = reset; // @[:@20218.4]
  assign RetimeWrapper_42_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@20220.4]
  assign RetimeWrapper_42_io_in = _T_577 & io_rPort_5_en_0; // @[package.scala 94:16:@20219.4]
  assign RetimeWrapper_43_clock = clock; // @[:@20225.4]
  assign RetimeWrapper_43_reset = reset; // @[:@20226.4]
  assign RetimeWrapper_43_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@20228.4]
  assign RetimeWrapper_43_io_in = _T_641 & io_rPort_5_en_0; // @[package.scala 94:16:@20227.4]
  assign RetimeWrapper_44_clock = clock; // @[:@20233.4]
  assign RetimeWrapper_44_reset = reset; // @[:@20234.4]
  assign RetimeWrapper_44_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@20236.4]
  assign RetimeWrapper_44_io_in = _T_705 & io_rPort_5_en_0; // @[package.scala 94:16:@20235.4]
  assign RetimeWrapper_45_clock = clock; // @[:@20241.4]
  assign RetimeWrapper_45_reset = reset; // @[:@20242.4]
  assign RetimeWrapper_45_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@20244.4]
  assign RetimeWrapper_45_io_in = _T_769 & io_rPort_5_en_0; // @[package.scala 94:16:@20243.4]
  assign RetimeWrapper_46_clock = clock; // @[:@20249.4]
  assign RetimeWrapper_46_reset = reset; // @[:@20250.4]
  assign RetimeWrapper_46_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@20252.4]
  assign RetimeWrapper_46_io_in = _T_833 & io_rPort_5_en_0; // @[package.scala 94:16:@20251.4]
  assign RetimeWrapper_47_clock = clock; // @[:@20257.4]
  assign RetimeWrapper_47_reset = reset; // @[:@20258.4]
  assign RetimeWrapper_47_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@20260.4]
  assign RetimeWrapper_47_io_in = _T_897 & io_rPort_5_en_0; // @[package.scala 94:16:@20259.4]
endmodule
module RetimeWrapper_230( // @[:@20675.2]
  input         clock, // @[:@20676.4]
  input         reset, // @[:@20677.4]
  input         io_flow, // @[:@20678.4]
  input  [31:0] io_in, // @[:@20678.4]
  output [31:0] io_out // @[:@20678.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@20680.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@20680.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@20680.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@20680.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@20680.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@20680.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@20680.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@20693.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@20692.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@20691.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@20690.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@20689.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@20687.4]
endmodule
module RetimeWrapper_232( // @[:@20739.2]
  input         clock, // @[:@20740.4]
  input         reset, // @[:@20741.4]
  input         io_flow, // @[:@20742.4]
  input  [31:0] io_in, // @[:@20742.4]
  output [31:0] io_out // @[:@20742.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@20744.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@20744.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@20744.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@20744.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@20744.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@20744.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@20744.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@20757.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@20756.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@20755.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@20754.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@20753.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@20751.4]
endmodule
module RetimeWrapper_243( // @[:@21385.2]
  input         clock, // @[:@21386.4]
  input         reset, // @[:@21387.4]
  input         io_flow, // @[:@21388.4]
  input  [31:0] io_in, // @[:@21388.4]
  output [31:0] io_out // @[:@21388.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21390.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21390.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21390.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21390.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21390.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21390.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@21390.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21403.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21402.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21401.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21400.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21399.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21397.4]
endmodule
module RetimeWrapper_246( // @[:@21481.2]
  input         clock, // @[:@21482.4]
  input         reset, // @[:@21483.4]
  input         io_flow, // @[:@21484.4]
  input  [31:0] io_in, // @[:@21484.4]
  output [31:0] io_out // @[:@21484.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21486.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21486.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21486.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21486.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21486.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21486.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@21486.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21499.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21498.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21497.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21496.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21495.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21493.4]
endmodule
module RetimeWrapper_248( // @[:@21545.2]
  input   clock, // @[:@21546.4]
  input   reset, // @[:@21547.4]
  input   io_flow, // @[:@21548.4]
  input   io_in, // @[:@21548.4]
  output  io_out // @[:@21548.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@21550.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@21550.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@21550.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21550.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21550.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21550.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(9)) sr ( // @[RetimeShiftRegister.scala 15:20:@21550.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21563.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21562.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@21561.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21560.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21559.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21557.4]
endmodule
module RetimeWrapper_249( // @[:@21577.2]
  input         clock, // @[:@21578.4]
  input         reset, // @[:@21579.4]
  input         io_flow, // @[:@21580.4]
  input  [31:0] io_in, // @[:@21580.4]
  output [31:0] io_out // @[:@21580.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21582.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21582.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21582.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21582.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21582.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21582.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(9)) sr ( // @[RetimeShiftRegister.scala 15:20:@21582.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21595.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21594.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21593.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21592.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21591.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21589.4]
endmodule
module RetimeWrapper_250( // @[:@21609.2]
  input         clock, // @[:@21610.4]
  input         reset, // @[:@21611.4]
  input         io_flow, // @[:@21612.4]
  input  [31:0] io_in, // @[:@21612.4]
  output [31:0] io_out // @[:@21612.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@21614.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@21614.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@21614.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@21614.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@21614.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@21614.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@21614.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@21627.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@21626.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@21625.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@21624.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@21623.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@21621.4]
endmodule
module Multiplier( // @[:@25755.2]
  input         clock, // @[:@25756.4]
  input         io_flow, // @[:@25758.4]
  input  [31:0] io_a, // @[:@25758.4]
  input  [31:0] io_b, // @[:@25758.4]
  output [31:0] io_out // @[:@25758.4]
);
  wire [31:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@25760.4]
  wire [31:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@25760.4]
  wire [31:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@25760.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@25760.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@25760.4]
  mul_32_32_32_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@25760.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@25770.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@25768.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@25767.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@25769.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@25766.4]
endmodule
module x385( // @[:@25790.2]
  input         clock, // @[:@25791.4]
  input  [31:0] io_a, // @[:@25793.4]
  input  [31:0] io_b, // @[:@25793.4]
  input         io_flow, // @[:@25793.4]
  output [31:0] io_result // @[:@25793.4]
);
  wire  x385_clock; // @[BigIPZynq.scala 63:21:@25800.4]
  wire  x385_io_flow; // @[BigIPZynq.scala 63:21:@25800.4]
  wire [31:0] x385_io_a; // @[BigIPZynq.scala 63:21:@25800.4]
  wire [31:0] x385_io_b; // @[BigIPZynq.scala 63:21:@25800.4]
  wire [31:0] x385_io_out; // @[BigIPZynq.scala 63:21:@25800.4]
  wire [31:0] fix2fixBox_io_a; // @[Math.scala 253:30:@25809.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@25809.4]
  Multiplier x385 ( // @[BigIPZynq.scala 63:21:@25800.4]
    .clock(x385_clock),
    .io_flow(x385_io_flow),
    .io_a(x385_io_a),
    .io_b(x385_io_b),
    .io_out(x385_io_out)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 253:30:@25809.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@25817.4]
  assign x385_clock = clock; // @[:@25801.4]
  assign x385_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@25805.4]
  assign x385_io_a = io_a; // @[BigIPZynq.scala 64:14:@25803.4]
  assign x385_io_b = io_b; // @[BigIPZynq.scala 65:14:@25804.4]
  assign fix2fixBox_io_a = x385_io_out; // @[Math.scala 254:23:@25812.4]
endmodule
module fix2fixBox_87( // @[:@26411.2]
  input  [31:0] io_a, // @[:@26414.4]
  output [32:0] io_b // @[:@26414.4]
);
  assign io_b = {1'h0,io_a}; // @[Converter.scala 95:38:@26428.4]
endmodule
module __52( // @[:@26430.2]
  input  [31:0] io_b, // @[:@26433.4]
  output [32:0] io_result // @[:@26433.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@26438.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@26438.4]
  fix2fixBox_87 fix2fixBox ( // @[BigIPZynq.scala 219:30:@26438.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@26446.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@26441.4]
endmodule
module x394_x7( // @[:@26542.2]
  input         clock, // @[:@26543.4]
  input         reset, // @[:@26544.4]
  input  [31:0] io_a, // @[:@26545.4]
  input  [31:0] io_b, // @[:@26545.4]
  input         io_flow, // @[:@26545.4]
  output [31:0] io_result // @[:@26545.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@26553.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@26553.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@26560.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@26560.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@26570.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@26570.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@26570.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@26570.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@26570.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@26558.4 Math.scala 724:14:@26559.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@26565.4 Math.scala 724:14:@26566.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@26567.4]
  __52 _ ( // @[Math.scala 720:24:@26553.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __52 __1 ( // @[Math.scala 720:24:@26560.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@26570.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@26558.4 Math.scala 724:14:@26559.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@26565.4 Math.scala 724:14:@26566.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@26567.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@26578.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@26556.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@26563.4]
  assign fix2fixBox_clock = clock; // @[:@26571.4]
  assign fix2fixBox_reset = reset; // @[:@26572.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@26573.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@26576.4]
endmodule
module fix2fixBox_111( // @[:@27795.2]
  input  [31:0] io_a, // @[:@27798.4]
  output [31:0] io_b // @[:@27798.4]
);
  wire [24:0] new_dec; // @[Converter.scala 63:26:@27808.4]
  assign new_dec = io_a[24:0]; // @[Converter.scala 63:26:@27808.4]
  assign io_b = {new_dec,7'h0}; // @[Converter.scala 94:38:@27811.4]
endmodule
module x402( // @[:@27813.2]
  input  [31:0] io_b, // @[:@27816.4]
  output [31:0] io_result // @[:@27816.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@27821.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@27821.4]
  fix2fixBox_111 fix2fixBox ( // @[BigIPZynq.scala 219:30:@27821.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@27829.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@27824.4]
endmodule
module Multiplier_9( // @[:@27841.2]
  input         clock, // @[:@27842.4]
  input         io_flow, // @[:@27844.4]
  input  [38:0] io_a, // @[:@27844.4]
  input  [38:0] io_b, // @[:@27844.4]
  output [38:0] io_out // @[:@27844.4]
);
  wire [38:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@27846.4]
  wire [38:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@27846.4]
  wire [38:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@27846.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@27846.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@27846.4]
  mul_39_39_39_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@27846.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@27856.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@27854.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@27853.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@27855.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@27852.4]
endmodule
module fix2fixBox_112( // @[:@27858.2]
  input  [38:0] io_a, // @[:@27861.4]
  output [31:0] io_b // @[:@27861.4]
);
  wire [6:0] tmp_frac; // @[Converter.scala 38:42:@27869.4]
  wire [24:0] new_dec; // @[Converter.scala 88:34:@27872.4]
  assign tmp_frac = io_a[13:7]; // @[Converter.scala 38:42:@27869.4]
  assign new_dec = io_a[38:14]; // @[Converter.scala 88:34:@27872.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@27875.4]
endmodule
module x403_mul( // @[:@27877.2]
  input         clock, // @[:@27878.4]
  input  [31:0] io_a, // @[:@27880.4]
  input  [31:0] io_b, // @[:@27880.4]
  input         io_flow, // @[:@27880.4]
  output [31:0] io_result // @[:@27880.4]
);
  wire  x403_mul_clock; // @[BigIPZynq.scala 63:21:@27895.4]
  wire  x403_mul_io_flow; // @[BigIPZynq.scala 63:21:@27895.4]
  wire [38:0] x403_mul_io_a; // @[BigIPZynq.scala 63:21:@27895.4]
  wire [38:0] x403_mul_io_b; // @[BigIPZynq.scala 63:21:@27895.4]
  wire [38:0] x403_mul_io_out; // @[BigIPZynq.scala 63:21:@27895.4]
  wire [38:0] fix2fixBox_io_a; // @[Math.scala 253:30:@27903.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@27903.4]
  wire  _T_16; // @[FixedPoint.scala 50:25:@27887.4]
  wire [6:0] _T_20; // @[Bitwise.scala 72:12:@27889.4]
  wire  _T_22; // @[FixedPoint.scala 50:25:@27891.4]
  wire [6:0] _T_26; // @[Bitwise.scala 72:12:@27893.4]
  Multiplier_9 x403_mul ( // @[BigIPZynq.scala 63:21:@27895.4]
    .clock(x403_mul_clock),
    .io_flow(x403_mul_io_flow),
    .io_a(x403_mul_io_a),
    .io_b(x403_mul_io_b),
    .io_out(x403_mul_io_out)
  );
  fix2fixBox_112 fix2fixBox ( // @[Math.scala 253:30:@27903.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_16 = io_a[31]; // @[FixedPoint.scala 50:25:@27887.4]
  assign _T_20 = _T_16 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@27889.4]
  assign _T_22 = io_b[31]; // @[FixedPoint.scala 50:25:@27891.4]
  assign _T_26 = _T_22 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@27893.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@27911.4]
  assign x403_mul_clock = clock; // @[:@27896.4]
  assign x403_mul_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@27900.4]
  assign x403_mul_io_a = {_T_20,io_a}; // @[BigIPZynq.scala 64:14:@27898.4]
  assign x403_mul_io_b = {_T_26,io_b}; // @[BigIPZynq.scala 65:14:@27899.4]
  assign fix2fixBox_io_a = x403_mul_io_out; // @[Math.scala 254:23:@27906.4]
endmodule
module fix2fixBox_113( // @[:@27913.2]
  input  [31:0] io_a, // @[:@27916.4]
  output [31:0] io_b // @[:@27916.4]
);
  wire [24:0] _T_25; // @[Converter.scala 84:75:@27928.4]
  assign _T_25 = io_a[31:7]; // @[Converter.scala 84:75:@27928.4]
  assign io_b = {7'h0,_T_25}; // @[Converter.scala 95:38:@27931.4]
endmodule
module x404( // @[:@27933.2]
  input  [31:0] io_b, // @[:@27936.4]
  output [31:0] io_result // @[:@27936.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@27941.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@27941.4]
  fix2fixBox_113 fix2fixBox ( // @[BigIPZynq.scala 219:30:@27941.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@27949.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@27944.4]
endmodule
module RetimeWrapper_325( // @[:@30201.2]
  input   clock, // @[:@30202.4]
  input   reset, // @[:@30203.4]
  input   io_flow, // @[:@30204.4]
  input   io_in, // @[:@30204.4]
  output  io_out // @[:@30204.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@30206.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@30206.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@30206.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30206.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30206.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30206.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(28)) sr ( // @[RetimeShiftRegister.scala 15:20:@30206.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30219.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30218.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@30217.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30216.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30215.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30213.4]
endmodule
module RetimeWrapper_326( // @[:@30233.2]
  input         clock, // @[:@30234.4]
  input         reset, // @[:@30235.4]
  input         io_flow, // @[:@30236.4]
  input  [31:0] io_in, // @[:@30236.4]
  output [31:0] io_out // @[:@30236.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@30238.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@30238.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@30238.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30238.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30238.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30238.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(28)) sr ( // @[RetimeShiftRegister.scala 15:20:@30238.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30251.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30250.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30249.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30248.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30247.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30245.4]
endmodule
module RetimeWrapper_328( // @[:@30297.2]
  input         clock, // @[:@30298.4]
  input         reset, // @[:@30299.4]
  input         io_flow, // @[:@30300.4]
  input  [31:0] io_in, // @[:@30300.4]
  output [31:0] io_out // @[:@30300.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@30302.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@30302.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@30302.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30302.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30302.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30302.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(26)) sr ( // @[RetimeShiftRegister.scala 15:20:@30302.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30315.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30314.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30313.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30312.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30311.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30309.4]
endmodule
module RetimeWrapper_333( // @[:@30457.2]
  input         clock, // @[:@30458.4]
  input         reset, // @[:@30459.4]
  input         io_flow, // @[:@30460.4]
  input  [31:0] io_in, // @[:@30460.4]
  output [31:0] io_out // @[:@30460.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@30462.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@30462.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@30462.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30462.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30462.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30462.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(27)) sr ( // @[RetimeShiftRegister.scala 15:20:@30462.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30475.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30474.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30473.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30472.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30471.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30469.4]
endmodule
module RetimeWrapper_336( // @[:@30553.2]
  input   clock, // @[:@30554.4]
  input   reset, // @[:@30555.4]
  input   io_flow, // @[:@30556.4]
  input   io_in, // @[:@30556.4]
  output  io_out // @[:@30556.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@30558.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@30558.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@30558.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30558.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30558.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30558.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(22)) sr ( // @[RetimeShiftRegister.scala 15:20:@30558.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30571.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30570.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@30569.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30568.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30567.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30565.4]
endmodule
module RetimeWrapper_337( // @[:@30585.2]
  input   clock, // @[:@30586.4]
  input   reset, // @[:@30587.4]
  input   io_flow, // @[:@30588.4]
  input   io_in, // @[:@30588.4]
  output  io_out // @[:@30588.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@30590.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@30590.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@30590.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30590.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30590.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30590.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(29)) sr ( // @[RetimeShiftRegister.scala 15:20:@30590.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30603.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30602.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@30601.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30600.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30599.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30597.4]
endmodule
module RetimeWrapper_338( // @[:@30617.2]
  input         clock, // @[:@30618.4]
  input         reset, // @[:@30619.4]
  input         io_flow, // @[:@30620.4]
  input  [31:0] io_in, // @[:@30620.4]
  output [31:0] io_out // @[:@30620.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@30622.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@30622.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@30622.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30622.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30622.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30622.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(29)) sr ( // @[RetimeShiftRegister.scala 15:20:@30622.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30635.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30634.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30633.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30632.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30631.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30629.4]
endmodule
module RetimeWrapper_342( // @[:@30745.2]
  input   clock, // @[:@30746.4]
  input   reset, // @[:@30747.4]
  input   io_flow, // @[:@30748.4]
  input   io_in, // @[:@30748.4]
  output  io_out // @[:@30748.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@30750.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@30750.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@30750.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30750.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30750.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30750.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(23)) sr ( // @[RetimeShiftRegister.scala 15:20:@30750.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30763.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30762.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@30761.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30760.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30759.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30757.4]
endmodule
module RetimeWrapper_346( // @[:@30873.2]
  input         clock, // @[:@30874.4]
  input         reset, // @[:@30875.4]
  input         io_flow, // @[:@30876.4]
  input  [31:0] io_in, // @[:@30876.4]
  output [31:0] io_out // @[:@30876.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@30878.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@30878.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@30878.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30878.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30878.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30878.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@30878.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30891.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30890.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30889.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30888.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30887.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30885.4]
endmodule
module RetimeWrapper_347( // @[:@30905.2]
  input         clock, // @[:@30906.4]
  input         reset, // @[:@30907.4]
  input         io_flow, // @[:@30908.4]
  input  [31:0] io_in, // @[:@30908.4]
  output [31:0] io_out // @[:@30908.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@30910.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@30910.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@30910.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@30910.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@30910.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@30910.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(22)) sr ( // @[RetimeShiftRegister.scala 15:20:@30910.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@30923.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@30922.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@30921.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@30920.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@30919.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@30917.4]
endmodule
module RetimeWrapper_351( // @[:@31033.2]
  input         clock, // @[:@31034.4]
  input         reset, // @[:@31035.4]
  input         io_flow, // @[:@31036.4]
  input  [31:0] io_in, // @[:@31036.4]
  output [31:0] io_out // @[:@31036.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@31038.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@31038.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@31038.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@31038.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@31038.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@31038.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@31038.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@31051.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@31050.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@31049.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@31048.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@31047.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@31045.4]
endmodule
module RetimeWrapper_366( // @[:@33239.2]
  input         clock, // @[:@33240.4]
  input         reset, // @[:@33241.4]
  input         io_flow, // @[:@33242.4]
  input  [63:0] io_in, // @[:@33242.4]
  output [63:0] io_out // @[:@33242.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@33244.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@33244.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@33244.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@33244.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@33244.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@33244.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@33244.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@33257.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@33256.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@33255.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@33254.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@33253.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@33251.4]
endmodule
module RetimeWrapper_367( // @[:@33271.2]
  input   clock, // @[:@33272.4]
  input   reset, // @[:@33273.4]
  input   io_flow, // @[:@33274.4]
  input   io_in, // @[:@33274.4]
  output  io_out // @[:@33274.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@33276.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@33276.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@33276.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@33276.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@33276.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@33276.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(48)) sr ( // @[RetimeShiftRegister.scala 15:20:@33276.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@33289.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@33288.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@33287.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@33286.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@33285.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@33283.4]
endmodule
module x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@33355.2]
  input          clock, // @[:@33356.4]
  input          reset, // @[:@33357.4]
  output         io_in_x251_TVALID, // @[:@33358.4]
  input          io_in_x251_TREADY, // @[:@33358.4]
  output [255:0] io_in_x251_TDATA, // @[:@33358.4]
  output         io_in_x250_TREADY, // @[:@33358.4]
  input  [255:0] io_in_x250_TDATA, // @[:@33358.4]
  input  [7:0]   io_in_x250_TID, // @[:@33358.4]
  input  [7:0]   io_in_x250_TDEST, // @[:@33358.4]
  input          io_sigsIn_backpressure, // @[:@33358.4]
  input          io_sigsIn_datapathEn, // @[:@33358.4]
  input          io_sigsIn_break, // @[:@33358.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@33358.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@33358.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@33358.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@33358.4]
  input          io_rr // @[:@33358.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@33372.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@33372.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@33384.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@33384.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@33407.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@33407.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@33407.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@33407.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@33407.4]
  wire  x285_lb_0_clock; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_reset; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_11_banks_1; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_11_banks_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [8:0] x285_lb_0_io_rPort_11_ofs_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_11_en_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_11_backpressure; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [31:0] x285_lb_0_io_rPort_11_output_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_10_banks_1; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_10_banks_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [8:0] x285_lb_0_io_rPort_10_ofs_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_10_en_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_10_backpressure; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [31:0] x285_lb_0_io_rPort_10_output_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_9_banks_1; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_9_banks_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [8:0] x285_lb_0_io_rPort_9_ofs_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_9_en_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_9_backpressure; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [31:0] x285_lb_0_io_rPort_9_output_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_8_banks_1; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_8_banks_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [8:0] x285_lb_0_io_rPort_8_ofs_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_8_en_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_8_backpressure; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [31:0] x285_lb_0_io_rPort_8_output_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_7_banks_1; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_7_banks_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [8:0] x285_lb_0_io_rPort_7_ofs_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_7_en_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_7_backpressure; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [31:0] x285_lb_0_io_rPort_7_output_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_6_banks_1; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_6_banks_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [8:0] x285_lb_0_io_rPort_6_ofs_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_6_en_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_6_backpressure; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [31:0] x285_lb_0_io_rPort_6_output_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_5_banks_1; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_5_banks_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [8:0] x285_lb_0_io_rPort_5_ofs_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_5_en_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_5_backpressure; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [31:0] x285_lb_0_io_rPort_5_output_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_4_banks_1; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_4_banks_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [8:0] x285_lb_0_io_rPort_4_ofs_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_4_en_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_4_backpressure; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [31:0] x285_lb_0_io_rPort_4_output_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_3_banks_1; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_3_banks_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [8:0] x285_lb_0_io_rPort_3_ofs_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_3_en_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_3_backpressure; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [31:0] x285_lb_0_io_rPort_3_output_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_2_banks_1; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_2_banks_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [8:0] x285_lb_0_io_rPort_2_ofs_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_2_en_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_2_backpressure; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [31:0] x285_lb_0_io_rPort_2_output_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_1_banks_1; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_1_banks_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [8:0] x285_lb_0_io_rPort_1_ofs_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_1_en_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_1_backpressure; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [31:0] x285_lb_0_io_rPort_1_output_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_0_banks_1; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_rPort_0_banks_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [8:0] x285_lb_0_io_rPort_0_ofs_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_0_en_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_rPort_0_backpressure; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [31:0] x285_lb_0_io_rPort_0_output_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_wPort_1_banks_1; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_wPort_1_banks_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [8:0] x285_lb_0_io_wPort_1_ofs_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [31:0] x285_lb_0_io_wPort_1_data_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_wPort_1_en_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_wPort_0_banks_1; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [2:0] x285_lb_0_io_wPort_0_banks_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [8:0] x285_lb_0_io_wPort_0_ofs_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire [31:0] x285_lb_0_io_wPort_0_data_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x285_lb_0_io_wPort_0_en_0; // @[m_x285_lb_0.scala 39:17:@33417.4]
  wire  x286_lb2_0_clock; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire  x286_lb2_0_reset; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [2:0] x286_lb2_0_io_rPort_5_banks_1; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [2:0] x286_lb2_0_io_rPort_5_banks_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [8:0] x286_lb2_0_io_rPort_5_ofs_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire  x286_lb2_0_io_rPort_5_en_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire  x286_lb2_0_io_rPort_5_backpressure; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [31:0] x286_lb2_0_io_rPort_5_output_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [2:0] x286_lb2_0_io_rPort_4_banks_1; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [2:0] x286_lb2_0_io_rPort_4_banks_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [8:0] x286_lb2_0_io_rPort_4_ofs_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire  x286_lb2_0_io_rPort_4_en_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire  x286_lb2_0_io_rPort_4_backpressure; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [31:0] x286_lb2_0_io_rPort_4_output_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [2:0] x286_lb2_0_io_rPort_3_banks_1; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [2:0] x286_lb2_0_io_rPort_3_banks_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [8:0] x286_lb2_0_io_rPort_3_ofs_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire  x286_lb2_0_io_rPort_3_en_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire  x286_lb2_0_io_rPort_3_backpressure; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [31:0] x286_lb2_0_io_rPort_3_output_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [2:0] x286_lb2_0_io_rPort_2_banks_1; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [2:0] x286_lb2_0_io_rPort_2_banks_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [8:0] x286_lb2_0_io_rPort_2_ofs_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire  x286_lb2_0_io_rPort_2_en_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire  x286_lb2_0_io_rPort_2_backpressure; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [31:0] x286_lb2_0_io_rPort_2_output_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [2:0] x286_lb2_0_io_rPort_1_banks_1; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [2:0] x286_lb2_0_io_rPort_1_banks_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [8:0] x286_lb2_0_io_rPort_1_ofs_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire  x286_lb2_0_io_rPort_1_en_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire  x286_lb2_0_io_rPort_1_backpressure; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [31:0] x286_lb2_0_io_rPort_1_output_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [2:0] x286_lb2_0_io_rPort_0_banks_1; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [2:0] x286_lb2_0_io_rPort_0_banks_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [8:0] x286_lb2_0_io_rPort_0_ofs_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire  x286_lb2_0_io_rPort_0_en_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire  x286_lb2_0_io_rPort_0_backpressure; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [31:0] x286_lb2_0_io_rPort_0_output_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [2:0] x286_lb2_0_io_wPort_1_banks_1; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [2:0] x286_lb2_0_io_wPort_1_banks_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [8:0] x286_lb2_0_io_wPort_1_ofs_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [31:0] x286_lb2_0_io_wPort_1_data_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire  x286_lb2_0_io_wPort_1_en_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [2:0] x286_lb2_0_io_wPort_0_banks_1; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [2:0] x286_lb2_0_io_wPort_0_banks_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [8:0] x286_lb2_0_io_wPort_0_ofs_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire [31:0] x286_lb2_0_io_wPort_0_data_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire  x286_lb2_0_io_wPort_0_en_0; // @[m_x286_lb2_0.scala 33:17:@33510.4]
  wire  x524_sub_1_clock; // @[Math.scala 191:24:@33637.4]
  wire  x524_sub_1_reset; // @[Math.scala 191:24:@33637.4]
  wire [31:0] x524_sub_1_io_a; // @[Math.scala 191:24:@33637.4]
  wire [31:0] x524_sub_1_io_b; // @[Math.scala 191:24:@33637.4]
  wire  x524_sub_1_io_flow; // @[Math.scala 191:24:@33637.4]
  wire [31:0] x524_sub_1_io_result; // @[Math.scala 191:24:@33637.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@33664.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@33664.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@33664.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@33664.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@33664.4]
  wire  x295_sum_1_clock; // @[Math.scala 150:24:@33673.4]
  wire  x295_sum_1_reset; // @[Math.scala 150:24:@33673.4]
  wire [31:0] x295_sum_1_io_a; // @[Math.scala 150:24:@33673.4]
  wire [31:0] x295_sum_1_io_b; // @[Math.scala 150:24:@33673.4]
  wire  x295_sum_1_io_flow; // @[Math.scala 150:24:@33673.4]
  wire [31:0] x295_sum_1_io_result; // @[Math.scala 150:24:@33673.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@33683.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@33683.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@33683.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@33683.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@33683.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@33692.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@33692.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@33692.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@33692.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@33692.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@33701.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@33701.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@33701.4]
  wire [31:0] RetimeWrapper_4_io_in; // @[package.scala 93:22:@33701.4]
  wire [31:0] RetimeWrapper_4_io_out; // @[package.scala 93:22:@33701.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@33710.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@33710.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@33710.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@33710.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@33710.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@33719.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@33719.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@33719.4]
  wire [31:0] RetimeWrapper_6_io_in; // @[package.scala 93:22:@33719.4]
  wire [31:0] RetimeWrapper_6_io_out; // @[package.scala 93:22:@33719.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@33728.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@33728.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@33728.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@33728.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@33728.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@33739.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@33739.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@33739.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@33739.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@33739.4]
  wire  x297_rdcol_1_clock; // @[Math.scala 150:24:@33762.4]
  wire  x297_rdcol_1_reset; // @[Math.scala 150:24:@33762.4]
  wire [31:0] x297_rdcol_1_io_a; // @[Math.scala 150:24:@33762.4]
  wire [31:0] x297_rdcol_1_io_b; // @[Math.scala 150:24:@33762.4]
  wire  x297_rdcol_1_io_flow; // @[Math.scala 150:24:@33762.4]
  wire [31:0] x297_rdcol_1_io_result; // @[Math.scala 150:24:@33762.4]
  wire  x301_sum_1_clock; // @[Math.scala 150:24:@33802.4]
  wire  x301_sum_1_reset; // @[Math.scala 150:24:@33802.4]
  wire [31:0] x301_sum_1_io_a; // @[Math.scala 150:24:@33802.4]
  wire [31:0] x301_sum_1_io_b; // @[Math.scala 150:24:@33802.4]
  wire  x301_sum_1_io_flow; // @[Math.scala 150:24:@33802.4]
  wire [31:0] x301_sum_1_io_result; // @[Math.scala 150:24:@33802.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@33812.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@33812.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@33812.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@33812.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@33812.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@33821.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@33821.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@33821.4]
  wire [31:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@33821.4]
  wire [31:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@33821.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@33830.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@33830.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@33830.4]
  wire [31:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@33830.4]
  wire [31:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@33830.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@33841.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@33841.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@33841.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@33841.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@33841.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@33862.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@33862.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@33862.4]
  wire [31:0] RetimeWrapper_13_io_in; // @[package.scala 93:22:@33862.4]
  wire [31:0] RetimeWrapper_13_io_out; // @[package.scala 93:22:@33862.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@33878.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@33878.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@33878.4]
  wire [31:0] RetimeWrapper_14_io_in; // @[package.scala 93:22:@33878.4]
  wire [31:0] RetimeWrapper_14_io_out; // @[package.scala 93:22:@33878.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@33894.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@33894.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@33894.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@33894.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@33894.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@33909.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@33909.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@33909.4]
  wire [31:0] RetimeWrapper_16_io_in; // @[package.scala 93:22:@33909.4]
  wire [31:0] RetimeWrapper_16_io_out; // @[package.scala 93:22:@33909.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@33918.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@33918.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@33918.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@33918.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@33918.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@33927.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@33927.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@33927.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@33927.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@33927.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@33936.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@33936.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@33936.4]
  wire [31:0] RetimeWrapper_19_io_in; // @[package.scala 93:22:@33936.4]
  wire [31:0] RetimeWrapper_19_io_out; // @[package.scala 93:22:@33936.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@33945.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@33945.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@33945.4]
  wire [31:0] RetimeWrapper_20_io_in; // @[package.scala 93:22:@33945.4]
  wire [31:0] RetimeWrapper_20_io_out; // @[package.scala 93:22:@33945.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@33954.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@33954.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@33954.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@33954.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@33954.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@33966.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@33966.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@33966.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@33966.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@33966.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@33987.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@33987.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@33987.4]
  wire [31:0] RetimeWrapper_23_io_in; // @[package.scala 93:22:@33987.4]
  wire [31:0] RetimeWrapper_23_io_out; // @[package.scala 93:22:@33987.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@34011.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@34011.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@34011.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@34011.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@34011.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@34020.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@34020.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@34020.4]
  wire [31:0] RetimeWrapper_25_io_in; // @[package.scala 93:22:@34020.4]
  wire [31:0] RetimeWrapper_25_io_out; // @[package.scala 93:22:@34020.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@34029.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@34029.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@34029.4]
  wire [31:0] RetimeWrapper_26_io_in; // @[package.scala 93:22:@34029.4]
  wire [31:0] RetimeWrapper_26_io_out; // @[package.scala 93:22:@34029.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@34041.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@34041.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@34041.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@34041.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@34041.4]
  wire  x315_rdcol_1_clock; // @[Math.scala 150:24:@34064.4]
  wire  x315_rdcol_1_reset; // @[Math.scala 150:24:@34064.4]
  wire [31:0] x315_rdcol_1_io_a; // @[Math.scala 150:24:@34064.4]
  wire [31:0] x315_rdcol_1_io_b; // @[Math.scala 150:24:@34064.4]
  wire  x315_rdcol_1_io_flow; // @[Math.scala 150:24:@34064.4]
  wire [31:0] x315_rdcol_1_io_result; // @[Math.scala 150:24:@34064.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@34115.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@34115.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@34115.4]
  wire [31:0] RetimeWrapper_28_io_in; // @[package.scala 93:22:@34115.4]
  wire [31:0] RetimeWrapper_28_io_out; // @[package.scala 93:22:@34115.4]
  wire  x321_sum_1_clock; // @[Math.scala 150:24:@34124.4]
  wire  x321_sum_1_reset; // @[Math.scala 150:24:@34124.4]
  wire [31:0] x321_sum_1_io_a; // @[Math.scala 150:24:@34124.4]
  wire [31:0] x321_sum_1_io_b; // @[Math.scala 150:24:@34124.4]
  wire  x321_sum_1_io_flow; // @[Math.scala 150:24:@34124.4]
  wire [31:0] x321_sum_1_io_result; // @[Math.scala 150:24:@34124.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@34134.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@34134.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@34134.4]
  wire [31:0] RetimeWrapper_29_io_in; // @[package.scala 93:22:@34134.4]
  wire [31:0] RetimeWrapper_29_io_out; // @[package.scala 93:22:@34134.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@34143.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@34143.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@34143.4]
  wire [31:0] RetimeWrapper_30_io_in; // @[package.scala 93:22:@34143.4]
  wire [31:0] RetimeWrapper_30_io_out; // @[package.scala 93:22:@34143.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@34152.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@34152.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@34152.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@34152.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@34152.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@34164.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@34164.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@34164.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@34164.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@34164.4]
  wire  x324_rdcol_1_clock; // @[Math.scala 150:24:@34187.4]
  wire  x324_rdcol_1_reset; // @[Math.scala 150:24:@34187.4]
  wire [31:0] x324_rdcol_1_io_a; // @[Math.scala 150:24:@34187.4]
  wire [31:0] x324_rdcol_1_io_b; // @[Math.scala 150:24:@34187.4]
  wire  x324_rdcol_1_io_flow; // @[Math.scala 150:24:@34187.4]
  wire [31:0] x324_rdcol_1_io_result; // @[Math.scala 150:24:@34187.4]
  wire  x330_sum_1_clock; // @[Math.scala 150:24:@34238.4]
  wire  x330_sum_1_reset; // @[Math.scala 150:24:@34238.4]
  wire [31:0] x330_sum_1_io_a; // @[Math.scala 150:24:@34238.4]
  wire [31:0] x330_sum_1_io_b; // @[Math.scala 150:24:@34238.4]
  wire  x330_sum_1_io_flow; // @[Math.scala 150:24:@34238.4]
  wire [31:0] x330_sum_1_io_result; // @[Math.scala 150:24:@34238.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@34248.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@34248.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@34248.4]
  wire [31:0] RetimeWrapper_33_io_in; // @[package.scala 93:22:@34248.4]
  wire [31:0] RetimeWrapper_33_io_out; // @[package.scala 93:22:@34248.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@34257.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@34257.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@34257.4]
  wire [31:0] RetimeWrapper_34_io_in; // @[package.scala 93:22:@34257.4]
  wire [31:0] RetimeWrapper_34_io_out; // @[package.scala 93:22:@34257.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@34266.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@34266.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@34266.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@34266.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@34266.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@34278.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@34278.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@34278.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@34278.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@34278.4]
  wire  x333_rdrow_1_clock; // @[Math.scala 191:24:@34301.4]
  wire  x333_rdrow_1_reset; // @[Math.scala 191:24:@34301.4]
  wire [31:0] x333_rdrow_1_io_a; // @[Math.scala 191:24:@34301.4]
  wire [31:0] x333_rdrow_1_io_b; // @[Math.scala 191:24:@34301.4]
  wire  x333_rdrow_1_io_flow; // @[Math.scala 191:24:@34301.4]
  wire [31:0] x333_rdrow_1_io_result; // @[Math.scala 191:24:@34301.4]
  wire  x532_sub_1_clock; // @[Math.scala 191:24:@34373.4]
  wire  x532_sub_1_reset; // @[Math.scala 191:24:@34373.4]
  wire [31:0] x532_sub_1_io_a; // @[Math.scala 191:24:@34373.4]
  wire [31:0] x532_sub_1_io_b; // @[Math.scala 191:24:@34373.4]
  wire  x532_sub_1_io_flow; // @[Math.scala 191:24:@34373.4]
  wire [31:0] x532_sub_1_io_result; // @[Math.scala 191:24:@34373.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@34383.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@34383.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@34383.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@34383.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@34383.4]
  wire  x341_sum_1_clock; // @[Math.scala 150:24:@34392.4]
  wire  x341_sum_1_reset; // @[Math.scala 150:24:@34392.4]
  wire [31:0] x341_sum_1_io_a; // @[Math.scala 150:24:@34392.4]
  wire [31:0] x341_sum_1_io_b; // @[Math.scala 150:24:@34392.4]
  wire  x341_sum_1_io_flow; // @[Math.scala 150:24:@34392.4]
  wire [31:0] x341_sum_1_io_result; // @[Math.scala 150:24:@34392.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@34402.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@34402.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@34402.4]
  wire [31:0] RetimeWrapper_38_io_in; // @[package.scala 93:22:@34402.4]
  wire [31:0] RetimeWrapper_38_io_out; // @[package.scala 93:22:@34402.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@34411.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@34411.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@34411.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@34411.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@34411.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@34423.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@34423.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@34423.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@34423.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@34423.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@34444.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@34444.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@34444.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@34444.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@34444.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@34459.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@34459.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@34459.4]
  wire [31:0] RetimeWrapper_42_io_in; // @[package.scala 93:22:@34459.4]
  wire [31:0] RetimeWrapper_42_io_out; // @[package.scala 93:22:@34459.4]
  wire  x346_sum_1_clock; // @[Math.scala 150:24:@34470.4]
  wire  x346_sum_1_reset; // @[Math.scala 150:24:@34470.4]
  wire [31:0] x346_sum_1_io_a; // @[Math.scala 150:24:@34470.4]
  wire [31:0] x346_sum_1_io_b; // @[Math.scala 150:24:@34470.4]
  wire  x346_sum_1_io_flow; // @[Math.scala 150:24:@34470.4]
  wire [31:0] x346_sum_1_io_result; // @[Math.scala 150:24:@34470.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@34480.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@34480.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@34480.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@34480.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@34480.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@34492.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@34492.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@34492.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@34492.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@34492.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@34519.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@34519.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@34519.4]
  wire [31:0] RetimeWrapper_45_io_in; // @[package.scala 93:22:@34519.4]
  wire [31:0] RetimeWrapper_45_io_out; // @[package.scala 93:22:@34519.4]
  wire  x351_sum_1_clock; // @[Math.scala 150:24:@34528.4]
  wire  x351_sum_1_reset; // @[Math.scala 150:24:@34528.4]
  wire [31:0] x351_sum_1_io_a; // @[Math.scala 150:24:@34528.4]
  wire [31:0] x351_sum_1_io_b; // @[Math.scala 150:24:@34528.4]
  wire  x351_sum_1_io_flow; // @[Math.scala 150:24:@34528.4]
  wire [31:0] x351_sum_1_io_result; // @[Math.scala 150:24:@34528.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@34538.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@34538.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@34538.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@34538.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@34538.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@34550.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@34550.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@34550.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@34550.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@34550.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@34577.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@34577.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@34577.4]
  wire [31:0] RetimeWrapper_48_io_in; // @[package.scala 93:22:@34577.4]
  wire [31:0] RetimeWrapper_48_io_out; // @[package.scala 93:22:@34577.4]
  wire  x356_sum_1_clock; // @[Math.scala 150:24:@34586.4]
  wire  x356_sum_1_reset; // @[Math.scala 150:24:@34586.4]
  wire [31:0] x356_sum_1_io_a; // @[Math.scala 150:24:@34586.4]
  wire [31:0] x356_sum_1_io_b; // @[Math.scala 150:24:@34586.4]
  wire  x356_sum_1_io_flow; // @[Math.scala 150:24:@34586.4]
  wire [31:0] x356_sum_1_io_result; // @[Math.scala 150:24:@34586.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@34596.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@34596.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@34596.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@34596.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@34596.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@34608.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@34608.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@34608.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@34608.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@34608.4]
  wire  x359_rdrow_1_clock; // @[Math.scala 191:24:@34631.4]
  wire  x359_rdrow_1_reset; // @[Math.scala 191:24:@34631.4]
  wire [31:0] x359_rdrow_1_io_a; // @[Math.scala 191:24:@34631.4]
  wire [31:0] x359_rdrow_1_io_b; // @[Math.scala 191:24:@34631.4]
  wire  x359_rdrow_1_io_flow; // @[Math.scala 191:24:@34631.4]
  wire [31:0] x359_rdrow_1_io_result; // @[Math.scala 191:24:@34631.4]
  wire  x537_sub_1_clock; // @[Math.scala 191:24:@34703.4]
  wire  x537_sub_1_reset; // @[Math.scala 191:24:@34703.4]
  wire [31:0] x537_sub_1_io_a; // @[Math.scala 191:24:@34703.4]
  wire [31:0] x537_sub_1_io_b; // @[Math.scala 191:24:@34703.4]
  wire  x537_sub_1_io_flow; // @[Math.scala 191:24:@34703.4]
  wire [31:0] x537_sub_1_io_result; // @[Math.scala 191:24:@34703.4]
  wire  x367_sum_1_clock; // @[Math.scala 150:24:@34713.4]
  wire  x367_sum_1_reset; // @[Math.scala 150:24:@34713.4]
  wire [31:0] x367_sum_1_io_a; // @[Math.scala 150:24:@34713.4]
  wire [31:0] x367_sum_1_io_b; // @[Math.scala 150:24:@34713.4]
  wire  x367_sum_1_io_flow; // @[Math.scala 150:24:@34713.4]
  wire [31:0] x367_sum_1_io_result; // @[Math.scala 150:24:@34713.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@34723.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@34723.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@34723.4]
  wire [31:0] RetimeWrapper_51_io_in; // @[package.scala 93:22:@34723.4]
  wire [31:0] RetimeWrapper_51_io_out; // @[package.scala 93:22:@34723.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@34732.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@34732.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@34732.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@34732.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@34732.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@34744.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@34744.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@34744.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@34744.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@34744.4]
  wire  x372_sum_1_clock; // @[Math.scala 150:24:@34771.4]
  wire  x372_sum_1_reset; // @[Math.scala 150:24:@34771.4]
  wire [31:0] x372_sum_1_io_a; // @[Math.scala 150:24:@34771.4]
  wire [31:0] x372_sum_1_io_b; // @[Math.scala 150:24:@34771.4]
  wire  x372_sum_1_io_flow; // @[Math.scala 150:24:@34771.4]
  wire [31:0] x372_sum_1_io_result; // @[Math.scala 150:24:@34771.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@34781.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@34781.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@34781.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@34781.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@34781.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@34793.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@34793.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@34793.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@34793.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@34793.4]
  wire  x377_sum_1_clock; // @[Math.scala 150:24:@34820.4]
  wire  x377_sum_1_reset; // @[Math.scala 150:24:@34820.4]
  wire [31:0] x377_sum_1_io_a; // @[Math.scala 150:24:@34820.4]
  wire [31:0] x377_sum_1_io_b; // @[Math.scala 150:24:@34820.4]
  wire  x377_sum_1_io_flow; // @[Math.scala 150:24:@34820.4]
  wire [31:0] x377_sum_1_io_result; // @[Math.scala 150:24:@34820.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@34830.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@34830.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@34830.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@34830.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@34830.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@34842.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@34842.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@34842.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@34842.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@34842.4]
  wire  x382_sum_1_clock; // @[Math.scala 150:24:@34871.4]
  wire  x382_sum_1_reset; // @[Math.scala 150:24:@34871.4]
  wire [31:0] x382_sum_1_io_a; // @[Math.scala 150:24:@34871.4]
  wire [31:0] x382_sum_1_io_b; // @[Math.scala 150:24:@34871.4]
  wire  x382_sum_1_io_flow; // @[Math.scala 150:24:@34871.4]
  wire [31:0] x382_sum_1_io_result; // @[Math.scala 150:24:@34871.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@34881.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@34881.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@34881.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@34881.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@34881.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@34893.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@34893.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@34893.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@34893.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@34893.4]
  wire  x385_1_clock; // @[Math.scala 262:24:@34916.4]
  wire [31:0] x385_1_io_a; // @[Math.scala 262:24:@34916.4]
  wire [31:0] x385_1_io_b; // @[Math.scala 262:24:@34916.4]
  wire  x385_1_io_flow; // @[Math.scala 262:24:@34916.4]
  wire [31:0] x385_1_io_result; // @[Math.scala 262:24:@34916.4]
  wire  x386_1_clock; // @[Math.scala 262:24:@34928.4]
  wire [31:0] x386_1_io_a; // @[Math.scala 262:24:@34928.4]
  wire [31:0] x386_1_io_b; // @[Math.scala 262:24:@34928.4]
  wire  x386_1_io_flow; // @[Math.scala 262:24:@34928.4]
  wire [31:0] x386_1_io_result; // @[Math.scala 262:24:@34928.4]
  wire  x387_1_clock; // @[Math.scala 262:24:@34940.4]
  wire [31:0] x387_1_io_a; // @[Math.scala 262:24:@34940.4]
  wire [31:0] x387_1_io_b; // @[Math.scala 262:24:@34940.4]
  wire  x387_1_io_flow; // @[Math.scala 262:24:@34940.4]
  wire [31:0] x387_1_io_result; // @[Math.scala 262:24:@34940.4]
  wire  x388_1_clock; // @[Math.scala 262:24:@34952.4]
  wire [31:0] x388_1_io_a; // @[Math.scala 262:24:@34952.4]
  wire [31:0] x388_1_io_b; // @[Math.scala 262:24:@34952.4]
  wire  x388_1_io_flow; // @[Math.scala 262:24:@34952.4]
  wire [31:0] x388_1_io_result; // @[Math.scala 262:24:@34952.4]
  wire  x389_1_clock; // @[Math.scala 262:24:@34964.4]
  wire [31:0] x389_1_io_a; // @[Math.scala 262:24:@34964.4]
  wire [31:0] x389_1_io_b; // @[Math.scala 262:24:@34964.4]
  wire  x389_1_io_flow; // @[Math.scala 262:24:@34964.4]
  wire [31:0] x389_1_io_result; // @[Math.scala 262:24:@34964.4]
  wire  x390_1_clock; // @[Math.scala 262:24:@34976.4]
  wire [31:0] x390_1_io_a; // @[Math.scala 262:24:@34976.4]
  wire [31:0] x390_1_io_b; // @[Math.scala 262:24:@34976.4]
  wire  x390_1_io_flow; // @[Math.scala 262:24:@34976.4]
  wire [31:0] x390_1_io_result; // @[Math.scala 262:24:@34976.4]
  wire  x391_1_clock; // @[Math.scala 262:24:@34988.4]
  wire [31:0] x391_1_io_a; // @[Math.scala 262:24:@34988.4]
  wire [31:0] x391_1_io_b; // @[Math.scala 262:24:@34988.4]
  wire  x391_1_io_flow; // @[Math.scala 262:24:@34988.4]
  wire [31:0] x391_1_io_result; // @[Math.scala 262:24:@34988.4]
  wire  x392_1_clock; // @[Math.scala 262:24:@35000.4]
  wire [31:0] x392_1_io_a; // @[Math.scala 262:24:@35000.4]
  wire [31:0] x392_1_io_b; // @[Math.scala 262:24:@35000.4]
  wire  x392_1_io_flow; // @[Math.scala 262:24:@35000.4]
  wire [31:0] x392_1_io_result; // @[Math.scala 262:24:@35000.4]
  wire  x393_1_clock; // @[Math.scala 262:24:@35012.4]
  wire [31:0] x393_1_io_a; // @[Math.scala 262:24:@35012.4]
  wire [31:0] x393_1_io_b; // @[Math.scala 262:24:@35012.4]
  wire  x393_1_io_flow; // @[Math.scala 262:24:@35012.4]
  wire [31:0] x393_1_io_result; // @[Math.scala 262:24:@35012.4]
  wire  x394_x7_1_clock; // @[Math.scala 150:24:@35022.4]
  wire  x394_x7_1_reset; // @[Math.scala 150:24:@35022.4]
  wire [31:0] x394_x7_1_io_a; // @[Math.scala 150:24:@35022.4]
  wire [31:0] x394_x7_1_io_b; // @[Math.scala 150:24:@35022.4]
  wire  x394_x7_1_io_flow; // @[Math.scala 150:24:@35022.4]
  wire [31:0] x394_x7_1_io_result; // @[Math.scala 150:24:@35022.4]
  wire  x395_x8_1_clock; // @[Math.scala 150:24:@35032.4]
  wire  x395_x8_1_reset; // @[Math.scala 150:24:@35032.4]
  wire [31:0] x395_x8_1_io_a; // @[Math.scala 150:24:@35032.4]
  wire [31:0] x395_x8_1_io_b; // @[Math.scala 150:24:@35032.4]
  wire  x395_x8_1_io_flow; // @[Math.scala 150:24:@35032.4]
  wire [31:0] x395_x8_1_io_result; // @[Math.scala 150:24:@35032.4]
  wire  x396_x7_1_clock; // @[Math.scala 150:24:@35042.4]
  wire  x396_x7_1_reset; // @[Math.scala 150:24:@35042.4]
  wire [31:0] x396_x7_1_io_a; // @[Math.scala 150:24:@35042.4]
  wire [31:0] x396_x7_1_io_b; // @[Math.scala 150:24:@35042.4]
  wire  x396_x7_1_io_flow; // @[Math.scala 150:24:@35042.4]
  wire [31:0] x396_x7_1_io_result; // @[Math.scala 150:24:@35042.4]
  wire  x397_x8_1_clock; // @[Math.scala 150:24:@35052.4]
  wire  x397_x8_1_reset; // @[Math.scala 150:24:@35052.4]
  wire [31:0] x397_x8_1_io_a; // @[Math.scala 150:24:@35052.4]
  wire [31:0] x397_x8_1_io_b; // @[Math.scala 150:24:@35052.4]
  wire  x397_x8_1_io_flow; // @[Math.scala 150:24:@35052.4]
  wire [31:0] x397_x8_1_io_result; // @[Math.scala 150:24:@35052.4]
  wire  x398_x7_1_clock; // @[Math.scala 150:24:@35062.4]
  wire  x398_x7_1_reset; // @[Math.scala 150:24:@35062.4]
  wire [31:0] x398_x7_1_io_a; // @[Math.scala 150:24:@35062.4]
  wire [31:0] x398_x7_1_io_b; // @[Math.scala 150:24:@35062.4]
  wire  x398_x7_1_io_flow; // @[Math.scala 150:24:@35062.4]
  wire [31:0] x398_x7_1_io_result; // @[Math.scala 150:24:@35062.4]
  wire  x399_x8_1_clock; // @[Math.scala 150:24:@35072.4]
  wire  x399_x8_1_reset; // @[Math.scala 150:24:@35072.4]
  wire [31:0] x399_x8_1_io_a; // @[Math.scala 150:24:@35072.4]
  wire [31:0] x399_x8_1_io_b; // @[Math.scala 150:24:@35072.4]
  wire  x399_x8_1_io_flow; // @[Math.scala 150:24:@35072.4]
  wire [31:0] x399_x8_1_io_result; // @[Math.scala 150:24:@35072.4]
  wire  x400_x7_1_clock; // @[Math.scala 150:24:@35082.4]
  wire  x400_x7_1_reset; // @[Math.scala 150:24:@35082.4]
  wire [31:0] x400_x7_1_io_a; // @[Math.scala 150:24:@35082.4]
  wire [31:0] x400_x7_1_io_b; // @[Math.scala 150:24:@35082.4]
  wire  x400_x7_1_io_flow; // @[Math.scala 150:24:@35082.4]
  wire [31:0] x400_x7_1_io_result; // @[Math.scala 150:24:@35082.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@35092.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@35092.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@35092.4]
  wire [31:0] RetimeWrapper_60_io_in; // @[package.scala 93:22:@35092.4]
  wire [31:0] RetimeWrapper_60_io_out; // @[package.scala 93:22:@35092.4]
  wire  x401_sum_1_clock; // @[Math.scala 150:24:@35101.4]
  wire  x401_sum_1_reset; // @[Math.scala 150:24:@35101.4]
  wire [31:0] x401_sum_1_io_a; // @[Math.scala 150:24:@35101.4]
  wire [31:0] x401_sum_1_io_b; // @[Math.scala 150:24:@35101.4]
  wire  x401_sum_1_io_flow; // @[Math.scala 150:24:@35101.4]
  wire [31:0] x401_sum_1_io_result; // @[Math.scala 150:24:@35101.4]
  wire [31:0] x402_1_io_b; // @[Math.scala 720:24:@35111.4]
  wire [31:0] x402_1_io_result; // @[Math.scala 720:24:@35111.4]
  wire  x403_mul_1_clock; // @[Math.scala 262:24:@35122.4]
  wire [31:0] x403_mul_1_io_a; // @[Math.scala 262:24:@35122.4]
  wire [31:0] x403_mul_1_io_b; // @[Math.scala 262:24:@35122.4]
  wire  x403_mul_1_io_flow; // @[Math.scala 262:24:@35122.4]
  wire [31:0] x403_mul_1_io_result; // @[Math.scala 262:24:@35122.4]
  wire [31:0] x404_1_io_b; // @[Math.scala 720:24:@35132.4]
  wire [31:0] x404_1_io_result; // @[Math.scala 720:24:@35132.4]
  wire  x405_1_clock; // @[Math.scala 262:24:@35143.4]
  wire [31:0] x405_1_io_a; // @[Math.scala 262:24:@35143.4]
  wire [31:0] x405_1_io_b; // @[Math.scala 262:24:@35143.4]
  wire  x405_1_io_flow; // @[Math.scala 262:24:@35143.4]
  wire [31:0] x405_1_io_result; // @[Math.scala 262:24:@35143.4]
  wire  x406_1_clock; // @[Math.scala 262:24:@35155.4]
  wire [31:0] x406_1_io_a; // @[Math.scala 262:24:@35155.4]
  wire [31:0] x406_1_io_b; // @[Math.scala 262:24:@35155.4]
  wire  x406_1_io_flow; // @[Math.scala 262:24:@35155.4]
  wire [31:0] x406_1_io_result; // @[Math.scala 262:24:@35155.4]
  wire  x407_1_clock; // @[Math.scala 262:24:@35167.4]
  wire [31:0] x407_1_io_a; // @[Math.scala 262:24:@35167.4]
  wire [31:0] x407_1_io_b; // @[Math.scala 262:24:@35167.4]
  wire  x407_1_io_flow; // @[Math.scala 262:24:@35167.4]
  wire [31:0] x407_1_io_result; // @[Math.scala 262:24:@35167.4]
  wire  x408_1_clock; // @[Math.scala 262:24:@35179.4]
  wire [31:0] x408_1_io_a; // @[Math.scala 262:24:@35179.4]
  wire [31:0] x408_1_io_b; // @[Math.scala 262:24:@35179.4]
  wire  x408_1_io_flow; // @[Math.scala 262:24:@35179.4]
  wire [31:0] x408_1_io_result; // @[Math.scala 262:24:@35179.4]
  wire  x409_1_clock; // @[Math.scala 262:24:@35191.4]
  wire [31:0] x409_1_io_a; // @[Math.scala 262:24:@35191.4]
  wire [31:0] x409_1_io_b; // @[Math.scala 262:24:@35191.4]
  wire  x409_1_io_flow; // @[Math.scala 262:24:@35191.4]
  wire [31:0] x409_1_io_result; // @[Math.scala 262:24:@35191.4]
  wire  x410_1_clock; // @[Math.scala 262:24:@35203.4]
  wire [31:0] x410_1_io_a; // @[Math.scala 262:24:@35203.4]
  wire [31:0] x410_1_io_b; // @[Math.scala 262:24:@35203.4]
  wire  x410_1_io_flow; // @[Math.scala 262:24:@35203.4]
  wire [31:0] x410_1_io_result; // @[Math.scala 262:24:@35203.4]
  wire  x411_1_clock; // @[Math.scala 262:24:@35215.4]
  wire [31:0] x411_1_io_a; // @[Math.scala 262:24:@35215.4]
  wire [31:0] x411_1_io_b; // @[Math.scala 262:24:@35215.4]
  wire  x411_1_io_flow; // @[Math.scala 262:24:@35215.4]
  wire [31:0] x411_1_io_result; // @[Math.scala 262:24:@35215.4]
  wire  x412_1_clock; // @[Math.scala 262:24:@35227.4]
  wire [31:0] x412_1_io_a; // @[Math.scala 262:24:@35227.4]
  wire [31:0] x412_1_io_b; // @[Math.scala 262:24:@35227.4]
  wire  x412_1_io_flow; // @[Math.scala 262:24:@35227.4]
  wire [31:0] x412_1_io_result; // @[Math.scala 262:24:@35227.4]
  wire  x413_1_clock; // @[Math.scala 262:24:@35239.4]
  wire [31:0] x413_1_io_a; // @[Math.scala 262:24:@35239.4]
  wire [31:0] x413_1_io_b; // @[Math.scala 262:24:@35239.4]
  wire  x413_1_io_flow; // @[Math.scala 262:24:@35239.4]
  wire [31:0] x413_1_io_result; // @[Math.scala 262:24:@35239.4]
  wire  x414_x7_1_clock; // @[Math.scala 150:24:@35249.4]
  wire  x414_x7_1_reset; // @[Math.scala 150:24:@35249.4]
  wire [31:0] x414_x7_1_io_a; // @[Math.scala 150:24:@35249.4]
  wire [31:0] x414_x7_1_io_b; // @[Math.scala 150:24:@35249.4]
  wire  x414_x7_1_io_flow; // @[Math.scala 150:24:@35249.4]
  wire [31:0] x414_x7_1_io_result; // @[Math.scala 150:24:@35249.4]
  wire  x415_x8_1_clock; // @[Math.scala 150:24:@35259.4]
  wire  x415_x8_1_reset; // @[Math.scala 150:24:@35259.4]
  wire [31:0] x415_x8_1_io_a; // @[Math.scala 150:24:@35259.4]
  wire [31:0] x415_x8_1_io_b; // @[Math.scala 150:24:@35259.4]
  wire  x415_x8_1_io_flow; // @[Math.scala 150:24:@35259.4]
  wire [31:0] x415_x8_1_io_result; // @[Math.scala 150:24:@35259.4]
  wire  x416_x7_1_clock; // @[Math.scala 150:24:@35269.4]
  wire  x416_x7_1_reset; // @[Math.scala 150:24:@35269.4]
  wire [31:0] x416_x7_1_io_a; // @[Math.scala 150:24:@35269.4]
  wire [31:0] x416_x7_1_io_b; // @[Math.scala 150:24:@35269.4]
  wire  x416_x7_1_io_flow; // @[Math.scala 150:24:@35269.4]
  wire [31:0] x416_x7_1_io_result; // @[Math.scala 150:24:@35269.4]
  wire  x417_x8_1_clock; // @[Math.scala 150:24:@35279.4]
  wire  x417_x8_1_reset; // @[Math.scala 150:24:@35279.4]
  wire [31:0] x417_x8_1_io_a; // @[Math.scala 150:24:@35279.4]
  wire [31:0] x417_x8_1_io_b; // @[Math.scala 150:24:@35279.4]
  wire  x417_x8_1_io_flow; // @[Math.scala 150:24:@35279.4]
  wire [31:0] x417_x8_1_io_result; // @[Math.scala 150:24:@35279.4]
  wire  x418_x7_1_clock; // @[Math.scala 150:24:@35289.4]
  wire  x418_x7_1_reset; // @[Math.scala 150:24:@35289.4]
  wire [31:0] x418_x7_1_io_a; // @[Math.scala 150:24:@35289.4]
  wire [31:0] x418_x7_1_io_b; // @[Math.scala 150:24:@35289.4]
  wire  x418_x7_1_io_flow; // @[Math.scala 150:24:@35289.4]
  wire [31:0] x418_x7_1_io_result; // @[Math.scala 150:24:@35289.4]
  wire  x419_x8_1_clock; // @[Math.scala 150:24:@35299.4]
  wire  x419_x8_1_reset; // @[Math.scala 150:24:@35299.4]
  wire [31:0] x419_x8_1_io_a; // @[Math.scala 150:24:@35299.4]
  wire [31:0] x419_x8_1_io_b; // @[Math.scala 150:24:@35299.4]
  wire  x419_x8_1_io_flow; // @[Math.scala 150:24:@35299.4]
  wire [31:0] x419_x8_1_io_result; // @[Math.scala 150:24:@35299.4]
  wire  x420_x7_1_clock; // @[Math.scala 150:24:@35309.4]
  wire  x420_x7_1_reset; // @[Math.scala 150:24:@35309.4]
  wire [31:0] x420_x7_1_io_a; // @[Math.scala 150:24:@35309.4]
  wire [31:0] x420_x7_1_io_b; // @[Math.scala 150:24:@35309.4]
  wire  x420_x7_1_io_flow; // @[Math.scala 150:24:@35309.4]
  wire [31:0] x420_x7_1_io_result; // @[Math.scala 150:24:@35309.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@35319.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@35319.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@35319.4]
  wire [31:0] RetimeWrapper_61_io_in; // @[package.scala 93:22:@35319.4]
  wire [31:0] RetimeWrapper_61_io_out; // @[package.scala 93:22:@35319.4]
  wire  x421_sum_1_clock; // @[Math.scala 150:24:@35328.4]
  wire  x421_sum_1_reset; // @[Math.scala 150:24:@35328.4]
  wire [31:0] x421_sum_1_io_a; // @[Math.scala 150:24:@35328.4]
  wire [31:0] x421_sum_1_io_b; // @[Math.scala 150:24:@35328.4]
  wire  x421_sum_1_io_flow; // @[Math.scala 150:24:@35328.4]
  wire [31:0] x421_sum_1_io_result; // @[Math.scala 150:24:@35328.4]
  wire [31:0] x422_1_io_b; // @[Math.scala 720:24:@35338.4]
  wire [31:0] x422_1_io_result; // @[Math.scala 720:24:@35338.4]
  wire  x423_mul_1_clock; // @[Math.scala 262:24:@35349.4]
  wire [31:0] x423_mul_1_io_a; // @[Math.scala 262:24:@35349.4]
  wire [31:0] x423_mul_1_io_b; // @[Math.scala 262:24:@35349.4]
  wire  x423_mul_1_io_flow; // @[Math.scala 262:24:@35349.4]
  wire [31:0] x423_mul_1_io_result; // @[Math.scala 262:24:@35349.4]
  wire [31:0] x424_1_io_b; // @[Math.scala 720:24:@35359.4]
  wire [31:0] x424_1_io_result; // @[Math.scala 720:24:@35359.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@35368.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@35368.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@35368.4]
  wire [31:0] RetimeWrapper_62_io_in; // @[package.scala 93:22:@35368.4]
  wire [31:0] RetimeWrapper_62_io_out; // @[package.scala 93:22:@35368.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@35377.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@35377.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@35377.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@35377.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@35377.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@35386.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@35386.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@35386.4]
  wire [31:0] RetimeWrapper_64_io_in; // @[package.scala 93:22:@35386.4]
  wire [31:0] RetimeWrapper_64_io_out; // @[package.scala 93:22:@35386.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@35395.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@35395.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@35395.4]
  wire [31:0] RetimeWrapper_65_io_in; // @[package.scala 93:22:@35395.4]
  wire [31:0] RetimeWrapper_65_io_out; // @[package.scala 93:22:@35395.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@35404.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@35404.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@35404.4]
  wire [31:0] RetimeWrapper_66_io_in; // @[package.scala 93:22:@35404.4]
  wire [31:0] RetimeWrapper_66_io_out; // @[package.scala 93:22:@35404.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@35413.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@35413.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@35413.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@35413.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@35413.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@35424.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@35424.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@35424.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@35424.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@35424.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@35445.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@35445.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@35445.4]
  wire [31:0] RetimeWrapper_69_io_in; // @[package.scala 93:22:@35445.4]
  wire [31:0] RetimeWrapper_69_io_out; // @[package.scala 93:22:@35445.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@35454.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@35454.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@35454.4]
  wire [31:0] RetimeWrapper_70_io_in; // @[package.scala 93:22:@35454.4]
  wire [31:0] RetimeWrapper_70_io_out; // @[package.scala 93:22:@35454.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@35463.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@35463.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@35463.4]
  wire [31:0] RetimeWrapper_71_io_in; // @[package.scala 93:22:@35463.4]
  wire [31:0] RetimeWrapper_71_io_out; // @[package.scala 93:22:@35463.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@35474.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@35474.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@35474.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@35474.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@35474.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@35495.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@35495.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@35495.4]
  wire [31:0] RetimeWrapper_73_io_in; // @[package.scala 93:22:@35495.4]
  wire [31:0] RetimeWrapper_73_io_out; // @[package.scala 93:22:@35495.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@35504.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@35504.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@35504.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@35504.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@35504.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@35513.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@35513.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@35513.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@35513.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@35513.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@35522.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@35522.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@35522.4]
  wire [31:0] RetimeWrapper_76_io_in; // @[package.scala 93:22:@35522.4]
  wire [31:0] RetimeWrapper_76_io_out; // @[package.scala 93:22:@35522.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@35531.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@35531.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@35531.4]
  wire [31:0] RetimeWrapper_77_io_in; // @[package.scala 93:22:@35531.4]
  wire [31:0] RetimeWrapper_77_io_out; // @[package.scala 93:22:@35531.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@35540.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@35540.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@35540.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@35540.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@35540.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@35552.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@35552.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@35552.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@35552.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@35552.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@35573.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@35573.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@35573.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@35573.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@35573.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@35582.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@35582.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@35582.4]
  wire [31:0] RetimeWrapper_81_io_in; // @[package.scala 93:22:@35582.4]
  wire [31:0] RetimeWrapper_81_io_out; // @[package.scala 93:22:@35582.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@35591.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@35591.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@35591.4]
  wire [31:0] RetimeWrapper_82_io_in; // @[package.scala 93:22:@35591.4]
  wire [31:0] RetimeWrapper_82_io_out; // @[package.scala 93:22:@35591.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@35603.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@35603.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@35603.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@35603.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@35603.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@35624.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@35624.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@35624.4]
  wire [31:0] RetimeWrapper_84_io_in; // @[package.scala 93:22:@35624.4]
  wire [31:0] RetimeWrapper_84_io_out; // @[package.scala 93:22:@35624.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@35633.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@35633.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@35633.4]
  wire [31:0] RetimeWrapper_85_io_in; // @[package.scala 93:22:@35633.4]
  wire [31:0] RetimeWrapper_85_io_out; // @[package.scala 93:22:@35633.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@35642.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@35642.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@35642.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@35642.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@35642.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@35654.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@35654.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@35654.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@35654.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@35654.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@35675.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@35675.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@35675.4]
  wire [31:0] RetimeWrapper_88_io_in; // @[package.scala 93:22:@35675.4]
  wire [31:0] RetimeWrapper_88_io_out; // @[package.scala 93:22:@35675.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@35684.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@35684.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@35684.4]
  wire [31:0] RetimeWrapper_89_io_in; // @[package.scala 93:22:@35684.4]
  wire [31:0] RetimeWrapper_89_io_out; // @[package.scala 93:22:@35684.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@35693.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@35693.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@35693.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@35693.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@35693.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@35705.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@35705.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@35705.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@35705.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@35705.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@35726.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@35726.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@35726.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@35726.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@35726.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@35735.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@35735.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@35735.4]
  wire [31:0] RetimeWrapper_93_io_in; // @[package.scala 93:22:@35735.4]
  wire [31:0] RetimeWrapper_93_io_out; // @[package.scala 93:22:@35735.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@35747.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@35747.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@35747.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@35747.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@35747.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@35768.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@35768.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@35768.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@35768.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@35768.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@35777.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@35777.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@35777.4]
  wire [31:0] RetimeWrapper_96_io_in; // @[package.scala 93:22:@35777.4]
  wire [31:0] RetimeWrapper_96_io_out; // @[package.scala 93:22:@35777.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@35789.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@35789.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@35789.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@35789.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@35789.4]
  wire  x441_1_clock; // @[Math.scala 262:24:@35814.4]
  wire [31:0] x441_1_io_a; // @[Math.scala 262:24:@35814.4]
  wire [31:0] x441_1_io_b; // @[Math.scala 262:24:@35814.4]
  wire  x441_1_io_flow; // @[Math.scala 262:24:@35814.4]
  wire [31:0] x441_1_io_result; // @[Math.scala 262:24:@35814.4]
  wire  x442_1_clock; // @[Math.scala 262:24:@35826.4]
  wire [31:0] x442_1_io_a; // @[Math.scala 262:24:@35826.4]
  wire [31:0] x442_1_io_b; // @[Math.scala 262:24:@35826.4]
  wire  x442_1_io_flow; // @[Math.scala 262:24:@35826.4]
  wire [31:0] x442_1_io_result; // @[Math.scala 262:24:@35826.4]
  wire  x443_1_clock; // @[Math.scala 262:24:@35838.4]
  wire [31:0] x443_1_io_a; // @[Math.scala 262:24:@35838.4]
  wire [31:0] x443_1_io_b; // @[Math.scala 262:24:@35838.4]
  wire  x443_1_io_flow; // @[Math.scala 262:24:@35838.4]
  wire [31:0] x443_1_io_result; // @[Math.scala 262:24:@35838.4]
  wire  x444_1_clock; // @[Math.scala 262:24:@35850.4]
  wire [31:0] x444_1_io_a; // @[Math.scala 262:24:@35850.4]
  wire [31:0] x444_1_io_b; // @[Math.scala 262:24:@35850.4]
  wire  x444_1_io_flow; // @[Math.scala 262:24:@35850.4]
  wire [31:0] x444_1_io_result; // @[Math.scala 262:24:@35850.4]
  wire  x445_x9_1_clock; // @[Math.scala 150:24:@35860.4]
  wire  x445_x9_1_reset; // @[Math.scala 150:24:@35860.4]
  wire [31:0] x445_x9_1_io_a; // @[Math.scala 150:24:@35860.4]
  wire [31:0] x445_x9_1_io_b; // @[Math.scala 150:24:@35860.4]
  wire  x445_x9_1_io_flow; // @[Math.scala 150:24:@35860.4]
  wire [31:0] x445_x9_1_io_result; // @[Math.scala 150:24:@35860.4]
  wire  x446_x10_1_clock; // @[Math.scala 150:24:@35872.4]
  wire  x446_x10_1_reset; // @[Math.scala 150:24:@35872.4]
  wire [31:0] x446_x10_1_io_a; // @[Math.scala 150:24:@35872.4]
  wire [31:0] x446_x10_1_io_b; // @[Math.scala 150:24:@35872.4]
  wire  x446_x10_1_io_flow; // @[Math.scala 150:24:@35872.4]
  wire [31:0] x446_x10_1_io_result; // @[Math.scala 150:24:@35872.4]
  wire  x447_sum_1_clock; // @[Math.scala 150:24:@35882.4]
  wire  x447_sum_1_reset; // @[Math.scala 150:24:@35882.4]
  wire [31:0] x447_sum_1_io_a; // @[Math.scala 150:24:@35882.4]
  wire [31:0] x447_sum_1_io_b; // @[Math.scala 150:24:@35882.4]
  wire  x447_sum_1_io_flow; // @[Math.scala 150:24:@35882.4]
  wire [31:0] x447_sum_1_io_result; // @[Math.scala 150:24:@35882.4]
  wire [31:0] x448_1_io_b; // @[Math.scala 720:24:@35892.4]
  wire [31:0] x448_1_io_result; // @[Math.scala 720:24:@35892.4]
  wire  x449_mul_1_clock; // @[Math.scala 262:24:@35903.4]
  wire [31:0] x449_mul_1_io_a; // @[Math.scala 262:24:@35903.4]
  wire [31:0] x449_mul_1_io_b; // @[Math.scala 262:24:@35903.4]
  wire  x449_mul_1_io_flow; // @[Math.scala 262:24:@35903.4]
  wire [31:0] x449_mul_1_io_result; // @[Math.scala 262:24:@35903.4]
  wire [31:0] x450_1_io_b; // @[Math.scala 720:24:@35913.4]
  wire [31:0] x450_1_io_result; // @[Math.scala 720:24:@35913.4]
  wire  x451_1_clock; // @[Math.scala 262:24:@35924.4]
  wire [31:0] x451_1_io_a; // @[Math.scala 262:24:@35924.4]
  wire [31:0] x451_1_io_b; // @[Math.scala 262:24:@35924.4]
  wire  x451_1_io_flow; // @[Math.scala 262:24:@35924.4]
  wire [31:0] x451_1_io_result; // @[Math.scala 262:24:@35924.4]
  wire  x452_1_clock; // @[Math.scala 262:24:@35936.4]
  wire [31:0] x452_1_io_a; // @[Math.scala 262:24:@35936.4]
  wire [31:0] x452_1_io_b; // @[Math.scala 262:24:@35936.4]
  wire  x452_1_io_flow; // @[Math.scala 262:24:@35936.4]
  wire [31:0] x452_1_io_result; // @[Math.scala 262:24:@35936.4]
  wire  x453_1_clock; // @[Math.scala 262:24:@35948.4]
  wire [31:0] x453_1_io_a; // @[Math.scala 262:24:@35948.4]
  wire [31:0] x453_1_io_b; // @[Math.scala 262:24:@35948.4]
  wire  x453_1_io_flow; // @[Math.scala 262:24:@35948.4]
  wire [31:0] x453_1_io_result; // @[Math.scala 262:24:@35948.4]
  wire  x454_1_clock; // @[Math.scala 262:24:@35960.4]
  wire [31:0] x454_1_io_a; // @[Math.scala 262:24:@35960.4]
  wire [31:0] x454_1_io_b; // @[Math.scala 262:24:@35960.4]
  wire  x454_1_io_flow; // @[Math.scala 262:24:@35960.4]
  wire [31:0] x454_1_io_result; // @[Math.scala 262:24:@35960.4]
  wire  x455_x9_1_clock; // @[Math.scala 150:24:@35970.4]
  wire  x455_x9_1_reset; // @[Math.scala 150:24:@35970.4]
  wire [31:0] x455_x9_1_io_a; // @[Math.scala 150:24:@35970.4]
  wire [31:0] x455_x9_1_io_b; // @[Math.scala 150:24:@35970.4]
  wire  x455_x9_1_io_flow; // @[Math.scala 150:24:@35970.4]
  wire [31:0] x455_x9_1_io_result; // @[Math.scala 150:24:@35970.4]
  wire  x456_x10_1_clock; // @[Math.scala 150:24:@35980.4]
  wire  x456_x10_1_reset; // @[Math.scala 150:24:@35980.4]
  wire [31:0] x456_x10_1_io_a; // @[Math.scala 150:24:@35980.4]
  wire [31:0] x456_x10_1_io_b; // @[Math.scala 150:24:@35980.4]
  wire  x456_x10_1_io_flow; // @[Math.scala 150:24:@35980.4]
  wire [31:0] x456_x10_1_io_result; // @[Math.scala 150:24:@35980.4]
  wire  x457_sum_1_clock; // @[Math.scala 150:24:@35990.4]
  wire  x457_sum_1_reset; // @[Math.scala 150:24:@35990.4]
  wire [31:0] x457_sum_1_io_a; // @[Math.scala 150:24:@35990.4]
  wire [31:0] x457_sum_1_io_b; // @[Math.scala 150:24:@35990.4]
  wire  x457_sum_1_io_flow; // @[Math.scala 150:24:@35990.4]
  wire [31:0] x457_sum_1_io_result; // @[Math.scala 150:24:@35990.4]
  wire [31:0] x458_1_io_b; // @[Math.scala 720:24:@36000.4]
  wire [31:0] x458_1_io_result; // @[Math.scala 720:24:@36000.4]
  wire  x459_mul_1_clock; // @[Math.scala 262:24:@36011.4]
  wire [31:0] x459_mul_1_io_a; // @[Math.scala 262:24:@36011.4]
  wire [31:0] x459_mul_1_io_b; // @[Math.scala 262:24:@36011.4]
  wire  x459_mul_1_io_flow; // @[Math.scala 262:24:@36011.4]
  wire [31:0] x459_mul_1_io_result; // @[Math.scala 262:24:@36011.4]
  wire [31:0] x460_1_io_b; // @[Math.scala 720:24:@36021.4]
  wire [31:0] x460_1_io_result; // @[Math.scala 720:24:@36021.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@36036.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@36036.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@36036.4]
  wire [63:0] RetimeWrapper_98_io_in; // @[package.scala 93:22:@36036.4]
  wire [63:0] RetimeWrapper_98_io_out; // @[package.scala 93:22:@36036.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@36045.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@36045.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@36045.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@36045.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@36045.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@36054.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@36054.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@36054.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@36054.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@36054.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@36063.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@36063.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@36063.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@36063.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@36063.4]
  wire  b281; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 62:18:@33392.4]
  wire  b282; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 63:18:@33393.4]
  wire  _T_205; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 67:30:@33395.4]
  wire  _T_206; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 67:37:@33396.4]
  wire  _T_210; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 69:76:@33401.4]
  wire  _T_211; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 69:62:@33402.4]
  wire  _T_213; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 69:101:@33403.4]
  wire [63:0] x543_x283_D1_0_number; // @[package.scala 96:25:@33412.4 package.scala 96:25:@33413.4]
  wire [31:0] b279_number; // @[Math.scala 723:22:@33377.4 Math.scala 724:14:@33378.4]
  wire [31:0] _T_244; // @[Math.scala 406:49:@33578.4]
  wire [31:0] _T_246; // @[Math.scala 406:56:@33580.4]
  wire [31:0] _T_247; // @[Math.scala 406:56:@33581.4]
  wire [31:0] x519_number; // @[implicits.scala 133:21:@33582.4]
  wire [31:0] _T_257; // @[Math.scala 406:49:@33591.4]
  wire [31:0] _T_259; // @[Math.scala 406:56:@33593.4]
  wire [31:0] _T_260; // @[Math.scala 406:56:@33594.4]
  wire [31:0] b280_number; // @[Math.scala 723:22:@33389.4 Math.scala 724:14:@33390.4]
  wire [31:0] _T_269; // @[Math.scala 406:49:@33602.4]
  wire [31:0] _T_271; // @[Math.scala 406:56:@33604.4]
  wire [31:0] _T_272; // @[Math.scala 406:56:@33605.4]
  wire  _T_276; // @[FixedPoint.scala 50:25:@33611.4]
  wire [1:0] _T_280; // @[Bitwise.scala 72:12:@33613.4]
  wire [29:0] _T_281; // @[FixedPoint.scala 18:52:@33614.4]
  wire  _T_287; // @[Math.scala 451:55:@33616.4]
  wire [1:0] _T_288; // @[FixedPoint.scala 18:52:@33617.4]
  wire  _T_294; // @[Math.scala 451:110:@33619.4]
  wire  _T_295; // @[Math.scala 451:94:@33620.4]
  wire [31:0] _T_297; // @[Cat.scala 30:58:@33622.4]
  wire [31:0] x292_1_number; // @[Math.scala 454:20:@33623.4]
  wire [40:0] _GEN_0; // @[Math.scala 461:32:@33628.4]
  wire [40:0] _T_302; // @[Math.scala 461:32:@33628.4]
  wire [36:0] _GEN_1; // @[Math.scala 461:32:@33633.4]
  wire [36:0] _T_305; // @[Math.scala 461:32:@33633.4]
  wire  _T_311; // @[FixedPoint.scala 50:25:@33648.4]
  wire [1:0] _T_315; // @[Bitwise.scala 72:12:@33650.4]
  wire [29:0] _T_316; // @[FixedPoint.scala 18:52:@33651.4]
  wire  _T_322; // @[Math.scala 451:55:@33653.4]
  wire [1:0] _T_323; // @[FixedPoint.scala 18:52:@33654.4]
  wire  _T_329; // @[Math.scala 451:110:@33656.4]
  wire  _T_330; // @[Math.scala 451:94:@33657.4]
  wire [31:0] _T_332; // @[Cat.scala 30:58:@33659.4]
  wire  _T_360; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 118:101:@33736.4]
  wire  _T_364; // @[package.scala 96:25:@33744.4 package.scala 96:25:@33745.4]
  wire  _T_366; // @[implicits.scala 55:10:@33746.4]
  wire  _T_367; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 118:118:@33747.4]
  wire  _T_369; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 118:206:@33749.4]
  wire  _T_370; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 118:225:@33750.4]
  wire  x546_b281_D3; // @[package.scala 96:25:@33697.4 package.scala 96:25:@33698.4]
  wire  _T_371; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 118:251:@33751.4]
  wire  x550_b282_D3; // @[package.scala 96:25:@33733.4 package.scala 96:25:@33734.4]
  wire [31:0] x297_rdcol_number; // @[Math.scala 154:22:@33768.4 Math.scala 155:14:@33769.4]
  wire [31:0] _T_388; // @[Math.scala 406:49:@33777.4]
  wire [31:0] _T_390; // @[Math.scala 406:56:@33779.4]
  wire [31:0] _T_391; // @[Math.scala 406:56:@33780.4]
  wire  _T_395; // @[FixedPoint.scala 50:25:@33786.4]
  wire [1:0] _T_399; // @[Bitwise.scala 72:12:@33788.4]
  wire [29:0] _T_400; // @[FixedPoint.scala 18:52:@33789.4]
  wire  _T_406; // @[Math.scala 451:55:@33791.4]
  wire [1:0] _T_407; // @[FixedPoint.scala 18:52:@33792.4]
  wire  _T_413; // @[Math.scala 451:110:@33794.4]
  wire  _T_414; // @[Math.scala 451:94:@33795.4]
  wire [31:0] _T_416; // @[Cat.scala 30:58:@33797.4]
  wire  _T_436; // @[package.scala 96:25:@33846.4 package.scala 96:25:@33847.4]
  wire  _T_438; // @[implicits.scala 55:10:@33848.4]
  wire  _T_439; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 139:118:@33849.4]
  wire  _T_441; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 139:206:@33851.4]
  wire  _T_442; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 139:225:@33852.4]
  wire  _T_443; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 139:251:@33853.4]
  wire [31:0] x554_b279_D6_number; // @[package.scala 96:25:@33867.4 package.scala 96:25:@33868.4]
  wire [31:0] _T_453; // @[Math.scala 476:37:@33873.4]
  wire  x304; // @[Math.scala 476:44:@33875.4]
  wire [31:0] x555_x297_rdcol_D6_number; // @[package.scala 96:25:@33883.4 package.scala 96:25:@33884.4]
  wire [31:0] _T_464; // @[Math.scala 476:37:@33889.4]
  wire  x305; // @[Math.scala 476:44:@33891.4]
  wire  x556_x304_D1; // @[package.scala 96:25:@33899.4 package.scala 96:25:@33900.4]
  wire  x306; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 152:24:@33903.4]
  wire  _T_503; // @[package.scala 96:25:@33971.4 package.scala 96:25:@33972.4]
  wire  _T_505; // @[implicits.scala 55:10:@33973.4]
  wire  _T_506; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 171:146:@33974.4]
  wire  x558_x307_D2; // @[package.scala 96:25:@33923.4 package.scala 96:25:@33924.4]
  wire  _T_507; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 171:234:@33975.4]
  wire  x559_b281_D9; // @[package.scala 96:25:@33932.4 package.scala 96:25:@33933.4]
  wire  _T_508; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 171:242:@33976.4]
  wire  x562_b282_D9; // @[package.scala 96:25:@33959.4 package.scala 96:25:@33960.4]
  wire [31:0] x563_b280_D6_number; // @[package.scala 96:25:@33992.4 package.scala 96:25:@33993.4]
  wire [31:0] _T_521; // @[Math.scala 476:37:@34000.4]
  wire  x310; // @[Math.scala 476:44:@34002.4]
  wire  x311; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 187:59:@34005.4]
  wire  _T_548; // @[package.scala 96:25:@34046.4 package.scala 96:25:@34047.4]
  wire  _T_550; // @[implicits.scala 55:10:@34048.4]
  wire  _T_551; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 200:194:@34049.4]
  wire  x564_x312_D3; // @[package.scala 96:25:@34016.4 package.scala 96:25:@34017.4]
  wire  _T_552; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 200:282:@34050.4]
  wire  _T_553; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 200:290:@34051.4]
  wire [31:0] x315_rdcol_number; // @[Math.scala 154:22:@34070.4 Math.scala 155:14:@34071.4]
  wire [31:0] _T_568; // @[Math.scala 476:37:@34076.4]
  wire  x316; // @[Math.scala 476:44:@34078.4]
  wire  x317; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 208:59:@34081.4]
  wire [31:0] _T_584; // @[Math.scala 406:56:@34092.4]
  wire [31:0] _T_585; // @[Math.scala 406:56:@34093.4]
  wire  _T_589; // @[FixedPoint.scala 50:25:@34099.4]
  wire [1:0] _T_593; // @[Bitwise.scala 72:12:@34101.4]
  wire [29:0] _T_594; // @[FixedPoint.scala 18:52:@34102.4]
  wire  _T_600; // @[Math.scala 451:55:@34104.4]
  wire [1:0] _T_601; // @[FixedPoint.scala 18:52:@34105.4]
  wire  _T_607; // @[Math.scala 451:110:@34107.4]
  wire  _T_608; // @[Math.scala 451:94:@34108.4]
  wire [31:0] _T_610; // @[Cat.scala 30:58:@34110.4]
  wire  _T_639; // @[package.scala 96:25:@34169.4 package.scala 96:25:@34170.4]
  wire  _T_641; // @[implicits.scala 55:10:@34171.4]
  wire  _T_642; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 229:194:@34172.4]
  wire  x570_x318_D2; // @[package.scala 96:25:@34157.4 package.scala 96:25:@34158.4]
  wire  _T_643; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 229:282:@34173.4]
  wire  _T_644; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 229:290:@34174.4]
  wire [31:0] x324_rdcol_number; // @[Math.scala 154:22:@34193.4 Math.scala 155:14:@34194.4]
  wire [31:0] _T_659; // @[Math.scala 476:37:@34199.4]
  wire  x325; // @[Math.scala 476:44:@34201.4]
  wire  x326; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 237:59:@34204.4]
  wire [31:0] _T_675; // @[Math.scala 406:56:@34215.4]
  wire [31:0] _T_676; // @[Math.scala 406:56:@34216.4]
  wire  _T_680; // @[FixedPoint.scala 50:25:@34222.4]
  wire [1:0] _T_684; // @[Bitwise.scala 72:12:@34224.4]
  wire [29:0] _T_685; // @[FixedPoint.scala 18:52:@34225.4]
  wire  _T_691; // @[Math.scala 451:55:@34227.4]
  wire [1:0] _T_692; // @[FixedPoint.scala 18:52:@34228.4]
  wire  _T_698; // @[Math.scala 451:110:@34230.4]
  wire  _T_699; // @[Math.scala 451:94:@34231.4]
  wire [31:0] _T_701; // @[Cat.scala 30:58:@34233.4]
  wire  _T_727; // @[package.scala 96:25:@34283.4 package.scala 96:25:@34284.4]
  wire  _T_729; // @[implicits.scala 55:10:@34285.4]
  wire  _T_730; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 256:194:@34286.4]
  wire  x573_x327_D2; // @[package.scala 96:25:@34271.4 package.scala 96:25:@34272.4]
  wire  _T_731; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 256:282:@34287.4]
  wire  _T_732; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 256:290:@34288.4]
  wire [31:0] x333_rdrow_number; // @[Math.scala 195:22:@34307.4 Math.scala 196:14:@34308.4]
  wire [31:0] _T_749; // @[Math.scala 406:49:@34314.4]
  wire [31:0] _T_751; // @[Math.scala 406:56:@34316.4]
  wire [31:0] _T_752; // @[Math.scala 406:56:@34317.4]
  wire [31:0] x528_number; // @[implicits.scala 133:21:@34318.4]
  wire  x335; // @[Math.scala 476:44:@34326.4]
  wire  x336; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 266:24:@34329.4]
  wire [31:0] _T_773; // @[Math.scala 406:49:@34338.4]
  wire [31:0] _T_775; // @[Math.scala 406:56:@34340.4]
  wire [31:0] _T_776; // @[Math.scala 406:56:@34341.4]
  wire  _T_780; // @[FixedPoint.scala 50:25:@34347.4]
  wire [1:0] _T_784; // @[Bitwise.scala 72:12:@34349.4]
  wire [29:0] _T_785; // @[FixedPoint.scala 18:52:@34350.4]
  wire  _T_791; // @[Math.scala 451:55:@34352.4]
  wire [1:0] _T_792; // @[FixedPoint.scala 18:52:@34353.4]
  wire  _T_798; // @[Math.scala 451:110:@34355.4]
  wire  _T_799; // @[Math.scala 451:94:@34356.4]
  wire [31:0] _T_801; // @[Cat.scala 30:58:@34358.4]
  wire [31:0] x339_1_number; // @[Math.scala 454:20:@34359.4]
  wire [40:0] _GEN_2; // @[Math.scala 461:32:@34364.4]
  wire [40:0] _T_806; // @[Math.scala 461:32:@34364.4]
  wire [36:0] _GEN_3; // @[Math.scala 461:32:@34369.4]
  wire [36:0] _T_809; // @[Math.scala 461:32:@34369.4]
  wire  _T_836; // @[package.scala 96:25:@34428.4 package.scala 96:25:@34429.4]
  wire  _T_838; // @[implicits.scala 55:10:@34430.4]
  wire  _T_839; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 291:194:@34431.4]
  wire  x576_x337_D2; // @[package.scala 96:25:@34416.4 package.scala 96:25:@34417.4]
  wire  _T_840; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 291:282:@34432.4]
  wire  _T_841; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 291:290:@34433.4]
  wire  x577_x310_D1; // @[package.scala 96:25:@34449.4 package.scala 96:25:@34450.4]
  wire  x344; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 303:59:@34453.4]
  wire  _T_873; // @[package.scala 96:25:@34497.4 package.scala 96:25:@34498.4]
  wire  _T_875; // @[implicits.scala 55:10:@34499.4]
  wire  _T_876; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 318:194:@34500.4]
  wire  x579_x345_D2; // @[package.scala 96:25:@34485.4 package.scala 96:25:@34486.4]
  wire  _T_877; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 318:282:@34501.4]
  wire  _T_878; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 318:290:@34502.4]
  wire  x349; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 322:59:@34513.4]
  wire  _T_905; // @[package.scala 96:25:@34555.4 package.scala 96:25:@34556.4]
  wire  _T_907; // @[implicits.scala 55:10:@34557.4]
  wire  _T_908; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 335:194:@34558.4]
  wire  x581_x350_D2; // @[package.scala 96:25:@34543.4 package.scala 96:25:@34544.4]
  wire  _T_909; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 335:282:@34559.4]
  wire  _T_910; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 335:290:@34560.4]
  wire  x354; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 339:59:@34571.4]
  wire  _T_937; // @[package.scala 96:25:@34613.4 package.scala 96:25:@34614.4]
  wire  _T_939; // @[implicits.scala 55:10:@34615.4]
  wire  _T_940; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 352:194:@34616.4]
  wire  x583_x355_D2; // @[package.scala 96:25:@34601.4 package.scala 96:25:@34602.4]
  wire  _T_941; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 352:282:@34617.4]
  wire  _T_942; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 352:290:@34618.4]
  wire [31:0] x359_rdrow_number; // @[Math.scala 195:22:@34637.4 Math.scala 196:14:@34638.4]
  wire [31:0] _T_959; // @[Math.scala 406:49:@34644.4]
  wire [31:0] _T_961; // @[Math.scala 406:56:@34646.4]
  wire [31:0] _T_962; // @[Math.scala 406:56:@34647.4]
  wire [31:0] x533_number; // @[implicits.scala 133:21:@34648.4]
  wire  x361; // @[Math.scala 476:44:@34656.4]
  wire  x362; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 362:24:@34659.4]
  wire [31:0] _T_983; // @[Math.scala 406:49:@34668.4]
  wire [31:0] _T_985; // @[Math.scala 406:56:@34670.4]
  wire [31:0] _T_986; // @[Math.scala 406:56:@34671.4]
  wire  _T_990; // @[FixedPoint.scala 50:25:@34677.4]
  wire [1:0] _T_994; // @[Bitwise.scala 72:12:@34679.4]
  wire [29:0] _T_995; // @[FixedPoint.scala 18:52:@34680.4]
  wire  _T_1001; // @[Math.scala 451:55:@34682.4]
  wire [1:0] _T_1002; // @[FixedPoint.scala 18:52:@34683.4]
  wire  _T_1008; // @[Math.scala 451:110:@34685.4]
  wire  _T_1009; // @[Math.scala 451:94:@34686.4]
  wire [31:0] _T_1011; // @[Cat.scala 30:58:@34688.4]
  wire [31:0] x365_1_number; // @[Math.scala 454:20:@34689.4]
  wire [40:0] _GEN_4; // @[Math.scala 461:32:@34694.4]
  wire [40:0] _T_1016; // @[Math.scala 461:32:@34694.4]
  wire [36:0] _GEN_5; // @[Math.scala 461:32:@34699.4]
  wire [36:0] _T_1019; // @[Math.scala 461:32:@34699.4]
  wire  _T_1043; // @[package.scala 96:25:@34749.4 package.scala 96:25:@34750.4]
  wire  _T_1045; // @[implicits.scala 55:10:@34751.4]
  wire  _T_1046; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 385:194:@34752.4]
  wire  x585_x363_D2; // @[package.scala 96:25:@34737.4 package.scala 96:25:@34738.4]
  wire  _T_1047; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 385:282:@34753.4]
  wire  _T_1048; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 385:290:@34754.4]
  wire  x370; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 389:24:@34765.4]
  wire  _T_1072; // @[package.scala 96:25:@34798.4 package.scala 96:25:@34799.4]
  wire  _T_1074; // @[implicits.scala 55:10:@34800.4]
  wire  _T_1075; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 400:194:@34801.4]
  wire  x586_x371_D2; // @[package.scala 96:25:@34786.4 package.scala 96:25:@34787.4]
  wire  _T_1076; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 400:282:@34802.4]
  wire  _T_1077; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 400:290:@34803.4]
  wire  x375; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 404:24:@34814.4]
  wire  _T_1101; // @[package.scala 96:25:@34847.4 package.scala 96:25:@34848.4]
  wire  _T_1103; // @[implicits.scala 55:10:@34849.4]
  wire  _T_1104; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 415:194:@34850.4]
  wire  x587_x376_D2; // @[package.scala 96:25:@34835.4 package.scala 96:25:@34836.4]
  wire  _T_1105; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 415:282:@34851.4]
  wire  _T_1106; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 415:290:@34852.4]
  wire  x380; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 425:59:@34863.4]
  wire  _T_1132; // @[package.scala 96:25:@34898.4 package.scala 96:25:@34899.4]
  wire  _T_1134; // @[implicits.scala 55:10:@34900.4]
  wire  _T_1135; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 438:194:@34901.4]
  wire  x588_x381_D2; // @[package.scala 96:25:@34886.4 package.scala 96:25:@34887.4]
  wire  _T_1136; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 438:282:@34902.4]
  wire  _T_1137; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 438:290:@34903.4]
  wire  _T_1369; // @[package.scala 96:25:@35429.4 package.scala 96:25:@35430.4]
  wire  _T_1371; // @[implicits.scala 55:10:@35431.4]
  wire  _T_1372; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 548:167:@35432.4]
  wire  _T_1374; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 548:256:@35434.4]
  wire  _T_1375; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 548:275:@35435.4]
  wire  x592_b281_D28; // @[package.scala 96:25:@35382.4 package.scala 96:25:@35383.4]
  wire  _T_1376; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 548:301:@35436.4]
  wire  x596_b282_D28; // @[package.scala 96:25:@35418.4 package.scala 96:25:@35419.4]
  wire  _T_1392; // @[package.scala 96:25:@35479.4 package.scala 96:25:@35480.4]
  wire  _T_1394; // @[implicits.scala 55:10:@35481.4]
  wire  _T_1395; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 559:167:@35482.4]
  wire  _T_1397; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 559:256:@35484.4]
  wire  _T_1398; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 559:275:@35485.4]
  wire  _T_1399; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 559:301:@35486.4]
  wire  _T_1430; // @[package.scala 96:25:@35557.4 package.scala 96:25:@35558.4]
  wire  _T_1432; // @[implicits.scala 55:10:@35559.4]
  wire  _T_1433; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 577:195:@35560.4]
  wire  x601_x307_D22; // @[package.scala 96:25:@35509.4 package.scala 96:25:@35510.4]
  wire  _T_1434; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 577:284:@35561.4]
  wire  x602_b281_D29; // @[package.scala 96:25:@35518.4 package.scala 96:25:@35519.4]
  wire  _T_1435; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 577:292:@35562.4]
  wire  x605_b282_D29; // @[package.scala 96:25:@35545.4 package.scala 96:25:@35546.4]
  wire  _T_1458; // @[package.scala 96:25:@35608.4 package.scala 96:25:@35609.4]
  wire  _T_1460; // @[implicits.scala 55:10:@35610.4]
  wire  _T_1461; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 590:195:@35611.4]
  wire  x606_x312_D23; // @[package.scala 96:25:@35578.4 package.scala 96:25:@35579.4]
  wire  _T_1462; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 590:284:@35612.4]
  wire  _T_1463; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 590:292:@35613.4]
  wire  _T_1486; // @[package.scala 96:25:@35659.4 package.scala 96:25:@35660.4]
  wire  _T_1488; // @[implicits.scala 55:10:@35661.4]
  wire  _T_1489; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 603:195:@35662.4]
  wire  x611_x318_D22; // @[package.scala 96:25:@35647.4 package.scala 96:25:@35648.4]
  wire  _T_1490; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 603:284:@35663.4]
  wire  _T_1491; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 603:292:@35664.4]
  wire  _T_1514; // @[package.scala 96:25:@35710.4 package.scala 96:25:@35711.4]
  wire  _T_1516; // @[implicits.scala 55:10:@35712.4]
  wire  _T_1517; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 616:195:@35713.4]
  wire  x614_x337_D22; // @[package.scala 96:25:@35698.4 package.scala 96:25:@35699.4]
  wire  _T_1518; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 616:284:@35714.4]
  wire  _T_1519; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 616:292:@35715.4]
  wire  _T_1539; // @[package.scala 96:25:@35752.4 package.scala 96:25:@35753.4]
  wire  _T_1541; // @[implicits.scala 55:10:@35754.4]
  wire  _T_1542; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 627:195:@35755.4]
  wire  x615_x345_D22; // @[package.scala 96:25:@35731.4 package.scala 96:25:@35732.4]
  wire  _T_1543; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 627:284:@35756.4]
  wire  _T_1544; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 627:292:@35757.4]
  wire  _T_1564; // @[package.scala 96:25:@35794.4 package.scala 96:25:@35795.4]
  wire  _T_1566; // @[implicits.scala 55:10:@35796.4]
  wire  _T_1567; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 638:195:@35797.4]
  wire  x617_x350_D22; // @[package.scala 96:25:@35773.4 package.scala 96:25:@35774.4]
  wire  _T_1568; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 638:284:@35798.4]
  wire  _T_1569; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 638:292:@35799.4]
  wire [31:0] x450_number; // @[Math.scala 723:22:@35918.4 Math.scala 724:14:@35919.4]
  wire [31:0] x460_number; // @[Math.scala 723:22:@36026.4 Math.scala 724:14:@36027.4]
  wire  _T_1697; // @[package.scala 96:25:@36068.4 package.scala 96:25:@36069.4]
  wire  _T_1699; // @[implicits.scala 55:10:@36070.4]
  wire  x620_b281_D48; // @[package.scala 96:25:@36059.4 package.scala 96:25:@36060.4]
  wire  _T_1700; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 700:117:@36071.4]
  wire  x619_b282_D48; // @[package.scala 96:25:@36050.4 package.scala 96:25:@36051.4]
  wire  _T_1701; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 700:123:@36072.4]
  wire [31:0] x547_x520_D3_number; // @[package.scala 96:25:@33706.4 package.scala 96:25:@33707.4]
  wire [31:0] x548_x521_D3_number; // @[package.scala 96:25:@33715.4 package.scala 96:25:@33716.4]
  wire [31:0] x549_x295_sum_D1_number; // @[package.scala 96:25:@33724.4 package.scala 96:25:@33725.4]
  wire [31:0] x551_x301_sum_D1_number; // @[package.scala 96:25:@33817.4 package.scala 96:25:@33818.4]
  wire [31:0] x553_x525_D2_number; // @[package.scala 96:25:@33835.4 package.scala 96:25:@33836.4]
  wire [31:0] x557_x301_sum_D7_number; // @[package.scala 96:25:@33914.4 package.scala 96:25:@33915.4]
  wire [31:0] x560_x520_D9_number; // @[package.scala 96:25:@33941.4 package.scala 96:25:@33942.4]
  wire [31:0] x561_x525_D8_number; // @[package.scala 96:25:@33950.4 package.scala 96:25:@33951.4]
  wire [31:0] x565_x521_D9_number; // @[package.scala 96:25:@34025.4 package.scala 96:25:@34026.4]
  wire [31:0] x566_x295_sum_D7_number; // @[package.scala 96:25:@34034.4 package.scala 96:25:@34035.4]
  wire [31:0] x568_x321_sum_D1_number; // @[package.scala 96:25:@34139.4 package.scala 96:25:@34140.4]
  wire [31:0] x569_x526_D2_number; // @[package.scala 96:25:@34148.4 package.scala 96:25:@34149.4]
  wire [31:0] x571_x527_D2_number; // @[package.scala 96:25:@34253.4 package.scala 96:25:@34254.4]
  wire [31:0] x572_x330_sum_D1_number; // @[package.scala 96:25:@34262.4 package.scala 96:25:@34263.4]
  wire [31:0] x341_sum_number; // @[Math.scala 154:22:@34398.4 Math.scala 155:14:@34399.4]
  wire [31:0] x575_x529_D2_number; // @[package.scala 96:25:@34407.4 package.scala 96:25:@34408.4]
  wire [31:0] x346_sum_number; // @[Math.scala 154:22:@34476.4 Math.scala 155:14:@34477.4]
  wire [31:0] x351_sum_number; // @[Math.scala 154:22:@34534.4 Math.scala 155:14:@34535.4]
  wire [31:0] x356_sum_number; // @[Math.scala 154:22:@34592.4 Math.scala 155:14:@34593.4]
  wire [31:0] x367_sum_number; // @[Math.scala 154:22:@34719.4 Math.scala 155:14:@34720.4]
  wire [31:0] x584_x534_D2_number; // @[package.scala 96:25:@34728.4 package.scala 96:25:@34729.4]
  wire [31:0] x372_sum_number; // @[Math.scala 154:22:@34777.4 Math.scala 155:14:@34778.4]
  wire [31:0] x377_sum_number; // @[Math.scala 154:22:@34826.4 Math.scala 155:14:@34827.4]
  wire [31:0] x382_sum_number; // @[Math.scala 154:22:@34877.4 Math.scala 155:14:@34878.4]
  wire [31:0] x593_x520_D28_number; // @[package.scala 96:25:@35391.4 package.scala 96:25:@35392.4]
  wire [31:0] x594_x521_D28_number; // @[package.scala 96:25:@35400.4 package.scala 96:25:@35401.4]
  wire [31:0] x595_x295_sum_D26_number; // @[package.scala 96:25:@35409.4 package.scala 96:25:@35410.4]
  wire [31:0] x598_x301_sum_D26_number; // @[package.scala 96:25:@35459.4 package.scala 96:25:@35460.4]
  wire [31:0] x599_x525_D27_number; // @[package.scala 96:25:@35468.4 package.scala 96:25:@35469.4]
  wire [31:0] x600_x301_sum_D27_number; // @[package.scala 96:25:@35500.4 package.scala 96:25:@35501.4]
  wire [31:0] x603_x520_D29_number; // @[package.scala 96:25:@35527.4 package.scala 96:25:@35528.4]
  wire [31:0] x604_x525_D28_number; // @[package.scala 96:25:@35536.4 package.scala 96:25:@35537.4]
  wire [31:0] x607_x521_D29_number; // @[package.scala 96:25:@35587.4 package.scala 96:25:@35588.4]
  wire [31:0] x608_x295_sum_D27_number; // @[package.scala 96:25:@35596.4 package.scala 96:25:@35597.4]
  wire [31:0] x609_x321_sum_D21_number; // @[package.scala 96:25:@35629.4 package.scala 96:25:@35630.4]
  wire [31:0] x610_x526_D22_number; // @[package.scala 96:25:@35638.4 package.scala 96:25:@35639.4]
  wire [31:0] x612_x529_D22_number; // @[package.scala 96:25:@35680.4 package.scala 96:25:@35681.4]
  wire [31:0] x613_x341_sum_D20_number; // @[package.scala 96:25:@35689.4 package.scala 96:25:@35690.4]
  wire [31:0] x616_x346_sum_D20_number; // @[package.scala 96:25:@35740.4 package.scala 96:25:@35741.4]
  wire [31:0] x618_x351_sum_D20_number; // @[package.scala 96:25:@35782.4 package.scala 96:25:@35783.4]
  _ _ ( // @[Math.scala 720:24:@33372.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@33384.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  RetimeWrapper_50 RetimeWrapper ( // @[package.scala 93:22:@33407.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x285_lb_0 x285_lb_0 ( // @[m_x285_lb_0.scala 39:17:@33417.4]
    .clock(x285_lb_0_clock),
    .reset(x285_lb_0_reset),
    .io_rPort_11_banks_1(x285_lb_0_io_rPort_11_banks_1),
    .io_rPort_11_banks_0(x285_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x285_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x285_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x285_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x285_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_1(x285_lb_0_io_rPort_10_banks_1),
    .io_rPort_10_banks_0(x285_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x285_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x285_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x285_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x285_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_1(x285_lb_0_io_rPort_9_banks_1),
    .io_rPort_9_banks_0(x285_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x285_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x285_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x285_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x285_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_1(x285_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x285_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x285_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x285_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x285_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x285_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x285_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x285_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x285_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x285_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x285_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x285_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x285_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x285_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x285_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x285_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x285_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x285_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x285_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x285_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x285_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x285_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x285_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x285_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x285_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x285_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x285_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x285_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x285_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x285_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x285_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x285_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x285_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x285_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x285_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x285_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x285_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x285_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x285_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x285_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x285_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x285_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x285_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x285_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x285_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x285_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x285_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x285_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x285_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x285_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x285_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x285_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x285_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x285_lb_0_io_rPort_0_output_0),
    .io_wPort_1_banks_1(x285_lb_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x285_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x285_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x285_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x285_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x285_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x285_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x285_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x285_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x285_lb_0_io_wPort_0_en_0)
  );
  x286_lb2_0 x286_lb2_0 ( // @[m_x286_lb2_0.scala 33:17:@33510.4]
    .clock(x286_lb2_0_clock),
    .reset(x286_lb2_0_reset),
    .io_rPort_5_banks_1(x286_lb2_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x286_lb2_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x286_lb2_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x286_lb2_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x286_lb2_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x286_lb2_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x286_lb2_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x286_lb2_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x286_lb2_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x286_lb2_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x286_lb2_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x286_lb2_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x286_lb2_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x286_lb2_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x286_lb2_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x286_lb2_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x286_lb2_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x286_lb2_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x286_lb2_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x286_lb2_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x286_lb2_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x286_lb2_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x286_lb2_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x286_lb2_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x286_lb2_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x286_lb2_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x286_lb2_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x286_lb2_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x286_lb2_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x286_lb2_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x286_lb2_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x286_lb2_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x286_lb2_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x286_lb2_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x286_lb2_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x286_lb2_0_io_rPort_0_output_0),
    .io_wPort_1_banks_1(x286_lb2_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x286_lb2_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x286_lb2_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x286_lb2_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x286_lb2_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x286_lb2_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x286_lb2_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x286_lb2_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x286_lb2_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x286_lb2_0_io_wPort_0_en_0)
  );
  x516_sub x524_sub_1 ( // @[Math.scala 191:24:@33637.4]
    .clock(x524_sub_1_clock),
    .reset(x524_sub_1_reset),
    .io_a(x524_sub_1_io_a),
    .io_b(x524_sub_1_io_b),
    .io_flow(x524_sub_1_io_flow),
    .io_result(x524_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_1 ( // @[package.scala 93:22:@33664.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x264_sum x295_sum_1 ( // @[Math.scala 150:24:@33673.4]
    .clock(x295_sum_1_clock),
    .reset(x295_sum_1_reset),
    .io_a(x295_sum_1_io_a),
    .io_b(x295_sum_1_io_b),
    .io_flow(x295_sum_1_io_flow),
    .io_result(x295_sum_1_io_result)
  );
  RetimeWrapper_230 RetimeWrapper_2 ( // @[package.scala 93:22:@33683.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_3 ( // @[package.scala 93:22:@33692.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_232 RetimeWrapper_4 ( // @[package.scala 93:22:@33701.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_232 RetimeWrapper_5 ( // @[package.scala 93:22:@33710.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_6 ( // @[package.scala 93:22:@33719.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_7 ( // @[package.scala 93:22:@33728.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_8 ( // @[package.scala 93:22:@33739.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  x264_sum x297_rdcol_1 ( // @[Math.scala 150:24:@33762.4]
    .clock(x297_rdcol_1_clock),
    .reset(x297_rdcol_1_reset),
    .io_a(x297_rdcol_1_io_a),
    .io_b(x297_rdcol_1_io_b),
    .io_flow(x297_rdcol_1_io_flow),
    .io_result(x297_rdcol_1_io_result)
  );
  x264_sum x301_sum_1 ( // @[Math.scala 150:24:@33802.4]
    .clock(x301_sum_1_clock),
    .reset(x301_sum_1_reset),
    .io_a(x301_sum_1_io_a),
    .io_b(x301_sum_1_io_b),
    .io_flow(x301_sum_1_io_flow),
    .io_result(x301_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_9 ( // @[package.scala 93:22:@33812.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_230 RetimeWrapper_10 ( // @[package.scala 93:22:@33821.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_230 RetimeWrapper_11 ( // @[package.scala 93:22:@33830.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_12 ( // @[package.scala 93:22:@33841.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_243 RetimeWrapper_13 ( // @[package.scala 93:22:@33862.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_243 RetimeWrapper_14 ( // @[package.scala 93:22:@33878.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 ( // @[package.scala 93:22:@33894.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_246 RetimeWrapper_16 ( // @[package.scala 93:22:@33909.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@33918.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_248 RetimeWrapper_18 ( // @[package.scala 93:22:@33927.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_249 RetimeWrapper_19 ( // @[package.scala 93:22:@33936.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_250 RetimeWrapper_20 ( // @[package.scala 93:22:@33945.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_248 RetimeWrapper_21 ( // @[package.scala 93:22:@33954.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_248 RetimeWrapper_22 ( // @[package.scala 93:22:@33966.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_243 RetimeWrapper_23 ( // @[package.scala 93:22:@33987.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_24 ( // @[package.scala 93:22:@34011.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_249 RetimeWrapper_25 ( // @[package.scala 93:22:@34020.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_246 RetimeWrapper_26 ( // @[package.scala 93:22:@34029.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_248 RetimeWrapper_27 ( // @[package.scala 93:22:@34041.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  x264_sum x315_rdcol_1 ( // @[Math.scala 150:24:@34064.4]
    .clock(x315_rdcol_1_clock),
    .reset(x315_rdcol_1_reset),
    .io_a(x315_rdcol_1_io_a),
    .io_b(x315_rdcol_1_io_b),
    .io_flow(x315_rdcol_1_io_flow),
    .io_result(x315_rdcol_1_io_result)
  );
  RetimeWrapper_243 RetimeWrapper_28 ( // @[package.scala 93:22:@34115.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  x264_sum x321_sum_1 ( // @[Math.scala 150:24:@34124.4]
    .clock(x321_sum_1_clock),
    .reset(x321_sum_1_reset),
    .io_a(x321_sum_1_io_a),
    .io_b(x321_sum_1_io_b),
    .io_flow(x321_sum_1_io_flow),
    .io_result(x321_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_29 ( // @[package.scala 93:22:@34134.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_230 RetimeWrapper_30 ( // @[package.scala 93:22:@34143.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@34152.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_248 RetimeWrapper_32 ( // @[package.scala 93:22:@34164.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  x264_sum x324_rdcol_1 ( // @[Math.scala 150:24:@34187.4]
    .clock(x324_rdcol_1_clock),
    .reset(x324_rdcol_1_reset),
    .io_a(x324_rdcol_1_io_a),
    .io_b(x324_rdcol_1_io_b),
    .io_flow(x324_rdcol_1_io_flow),
    .io_result(x324_rdcol_1_io_result)
  );
  x264_sum x330_sum_1 ( // @[Math.scala 150:24:@34238.4]
    .clock(x330_sum_1_clock),
    .reset(x330_sum_1_reset),
    .io_a(x330_sum_1_io_a),
    .io_b(x330_sum_1_io_b),
    .io_flow(x330_sum_1_io_flow),
    .io_result(x330_sum_1_io_result)
  );
  RetimeWrapper_230 RetimeWrapper_33 ( // @[package.scala 93:22:@34248.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_34 ( // @[package.scala 93:22:@34257.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@34266.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_248 RetimeWrapper_36 ( // @[package.scala 93:22:@34278.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  x516_sub x333_rdrow_1 ( // @[Math.scala 191:24:@34301.4]
    .clock(x333_rdrow_1_clock),
    .reset(x333_rdrow_1_reset),
    .io_a(x333_rdrow_1_io_a),
    .io_b(x333_rdrow_1_io_b),
    .io_flow(x333_rdrow_1_io_flow),
    .io_result(x333_rdrow_1_io_result)
  );
  x516_sub x532_sub_1 ( // @[Math.scala 191:24:@34373.4]
    .clock(x532_sub_1_clock),
    .reset(x532_sub_1_reset),
    .io_a(x532_sub_1_io_a),
    .io_b(x532_sub_1_io_b),
    .io_flow(x532_sub_1_io_flow),
    .io_result(x532_sub_1_io_result)
  );
  RetimeWrapper_246 RetimeWrapper_37 ( // @[package.scala 93:22:@34383.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  x264_sum x341_sum_1 ( // @[Math.scala 150:24:@34392.4]
    .clock(x341_sum_1_clock),
    .reset(x341_sum_1_reset),
    .io_a(x341_sum_1_io_a),
    .io_b(x341_sum_1_io_b),
    .io_flow(x341_sum_1_io_flow),
    .io_result(x341_sum_1_io_result)
  );
  RetimeWrapper_230 RetimeWrapper_38 ( // @[package.scala 93:22:@34402.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@34411.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_248 RetimeWrapper_40 ( // @[package.scala 93:22:@34423.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper RetimeWrapper_41 ( // @[package.scala 93:22:@34444.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_250 RetimeWrapper_42 ( // @[package.scala 93:22:@34459.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  x264_sum x346_sum_1 ( // @[Math.scala 150:24:@34470.4]
    .clock(x346_sum_1_clock),
    .reset(x346_sum_1_reset),
    .io_a(x346_sum_1_io_a),
    .io_b(x346_sum_1_io_b),
    .io_flow(x346_sum_1_io_flow),
    .io_result(x346_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@34480.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_248 RetimeWrapper_44 ( // @[package.scala 93:22:@34492.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_45 ( // @[package.scala 93:22:@34519.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  x264_sum x351_sum_1 ( // @[Math.scala 150:24:@34528.4]
    .clock(x351_sum_1_clock),
    .reset(x351_sum_1_reset),
    .io_a(x351_sum_1_io_a),
    .io_b(x351_sum_1_io_b),
    .io_flow(x351_sum_1_io_flow),
    .io_result(x351_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@34538.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_248 RetimeWrapper_47 ( // @[package.scala 93:22:@34550.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_48 ( // @[package.scala 93:22:@34577.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  x264_sum x356_sum_1 ( // @[Math.scala 150:24:@34586.4]
    .clock(x356_sum_1_clock),
    .reset(x356_sum_1_reset),
    .io_a(x356_sum_1_io_a),
    .io_b(x356_sum_1_io_b),
    .io_flow(x356_sum_1_io_flow),
    .io_result(x356_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@34596.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_248 RetimeWrapper_50 ( // @[package.scala 93:22:@34608.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  x516_sub x359_rdrow_1 ( // @[Math.scala 191:24:@34631.4]
    .clock(x359_rdrow_1_clock),
    .reset(x359_rdrow_1_reset),
    .io_a(x359_rdrow_1_io_a),
    .io_b(x359_rdrow_1_io_b),
    .io_flow(x359_rdrow_1_io_flow),
    .io_result(x359_rdrow_1_io_result)
  );
  x516_sub x537_sub_1 ( // @[Math.scala 191:24:@34703.4]
    .clock(x537_sub_1_clock),
    .reset(x537_sub_1_reset),
    .io_a(x537_sub_1_io_a),
    .io_b(x537_sub_1_io_b),
    .io_flow(x537_sub_1_io_flow),
    .io_result(x537_sub_1_io_result)
  );
  x264_sum x367_sum_1 ( // @[Math.scala 150:24:@34713.4]
    .clock(x367_sum_1_clock),
    .reset(x367_sum_1_reset),
    .io_a(x367_sum_1_io_a),
    .io_b(x367_sum_1_io_b),
    .io_flow(x367_sum_1_io_flow),
    .io_result(x367_sum_1_io_result)
  );
  RetimeWrapper_230 RetimeWrapper_51 ( // @[package.scala 93:22:@34723.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@34732.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_248 RetimeWrapper_53 ( // @[package.scala 93:22:@34744.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  x264_sum x372_sum_1 ( // @[Math.scala 150:24:@34771.4]
    .clock(x372_sum_1_clock),
    .reset(x372_sum_1_reset),
    .io_a(x372_sum_1_io_a),
    .io_b(x372_sum_1_io_b),
    .io_flow(x372_sum_1_io_flow),
    .io_result(x372_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@34781.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_248 RetimeWrapper_55 ( // @[package.scala 93:22:@34793.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  x264_sum x377_sum_1 ( // @[Math.scala 150:24:@34820.4]
    .clock(x377_sum_1_clock),
    .reset(x377_sum_1_reset),
    .io_a(x377_sum_1_io_a),
    .io_b(x377_sum_1_io_b),
    .io_flow(x377_sum_1_io_flow),
    .io_result(x377_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@34830.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_248 RetimeWrapper_57 ( // @[package.scala 93:22:@34842.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  x264_sum x382_sum_1 ( // @[Math.scala 150:24:@34871.4]
    .clock(x382_sum_1_clock),
    .reset(x382_sum_1_reset),
    .io_a(x382_sum_1_io_a),
    .io_b(x382_sum_1_io_b),
    .io_flow(x382_sum_1_io_flow),
    .io_result(x382_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@34881.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_248 RetimeWrapper_59 ( // @[package.scala 93:22:@34893.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  x385 x385_1 ( // @[Math.scala 262:24:@34916.4]
    .clock(x385_1_clock),
    .io_a(x385_1_io_a),
    .io_b(x385_1_io_b),
    .io_flow(x385_1_io_flow),
    .io_result(x385_1_io_result)
  );
  x385 x386_1 ( // @[Math.scala 262:24:@34928.4]
    .clock(x386_1_clock),
    .io_a(x386_1_io_a),
    .io_b(x386_1_io_b),
    .io_flow(x386_1_io_flow),
    .io_result(x386_1_io_result)
  );
  x385 x387_1 ( // @[Math.scala 262:24:@34940.4]
    .clock(x387_1_clock),
    .io_a(x387_1_io_a),
    .io_b(x387_1_io_b),
    .io_flow(x387_1_io_flow),
    .io_result(x387_1_io_result)
  );
  x385 x388_1 ( // @[Math.scala 262:24:@34952.4]
    .clock(x388_1_clock),
    .io_a(x388_1_io_a),
    .io_b(x388_1_io_b),
    .io_flow(x388_1_io_flow),
    .io_result(x388_1_io_result)
  );
  x385 x389_1 ( // @[Math.scala 262:24:@34964.4]
    .clock(x389_1_clock),
    .io_a(x389_1_io_a),
    .io_b(x389_1_io_b),
    .io_flow(x389_1_io_flow),
    .io_result(x389_1_io_result)
  );
  x385 x390_1 ( // @[Math.scala 262:24:@34976.4]
    .clock(x390_1_clock),
    .io_a(x390_1_io_a),
    .io_b(x390_1_io_b),
    .io_flow(x390_1_io_flow),
    .io_result(x390_1_io_result)
  );
  x385 x391_1 ( // @[Math.scala 262:24:@34988.4]
    .clock(x391_1_clock),
    .io_a(x391_1_io_a),
    .io_b(x391_1_io_b),
    .io_flow(x391_1_io_flow),
    .io_result(x391_1_io_result)
  );
  x385 x392_1 ( // @[Math.scala 262:24:@35000.4]
    .clock(x392_1_clock),
    .io_a(x392_1_io_a),
    .io_b(x392_1_io_b),
    .io_flow(x392_1_io_flow),
    .io_result(x392_1_io_result)
  );
  x385 x393_1 ( // @[Math.scala 262:24:@35012.4]
    .clock(x393_1_clock),
    .io_a(x393_1_io_a),
    .io_b(x393_1_io_b),
    .io_flow(x393_1_io_flow),
    .io_result(x393_1_io_result)
  );
  x394_x7 x394_x7_1 ( // @[Math.scala 150:24:@35022.4]
    .clock(x394_x7_1_clock),
    .reset(x394_x7_1_reset),
    .io_a(x394_x7_1_io_a),
    .io_b(x394_x7_1_io_b),
    .io_flow(x394_x7_1_io_flow),
    .io_result(x394_x7_1_io_result)
  );
  x394_x7 x395_x8_1 ( // @[Math.scala 150:24:@35032.4]
    .clock(x395_x8_1_clock),
    .reset(x395_x8_1_reset),
    .io_a(x395_x8_1_io_a),
    .io_b(x395_x8_1_io_b),
    .io_flow(x395_x8_1_io_flow),
    .io_result(x395_x8_1_io_result)
  );
  x394_x7 x396_x7_1 ( // @[Math.scala 150:24:@35042.4]
    .clock(x396_x7_1_clock),
    .reset(x396_x7_1_reset),
    .io_a(x396_x7_1_io_a),
    .io_b(x396_x7_1_io_b),
    .io_flow(x396_x7_1_io_flow),
    .io_result(x396_x7_1_io_result)
  );
  x394_x7 x397_x8_1 ( // @[Math.scala 150:24:@35052.4]
    .clock(x397_x8_1_clock),
    .reset(x397_x8_1_reset),
    .io_a(x397_x8_1_io_a),
    .io_b(x397_x8_1_io_b),
    .io_flow(x397_x8_1_io_flow),
    .io_result(x397_x8_1_io_result)
  );
  x394_x7 x398_x7_1 ( // @[Math.scala 150:24:@35062.4]
    .clock(x398_x7_1_clock),
    .reset(x398_x7_1_reset),
    .io_a(x398_x7_1_io_a),
    .io_b(x398_x7_1_io_b),
    .io_flow(x398_x7_1_io_flow),
    .io_result(x398_x7_1_io_result)
  );
  x394_x7 x399_x8_1 ( // @[Math.scala 150:24:@35072.4]
    .clock(x399_x8_1_clock),
    .reset(x399_x8_1_reset),
    .io_a(x399_x8_1_io_a),
    .io_b(x399_x8_1_io_b),
    .io_flow(x399_x8_1_io_flow),
    .io_result(x399_x8_1_io_result)
  );
  x394_x7 x400_x7_1 ( // @[Math.scala 150:24:@35082.4]
    .clock(x400_x7_1_clock),
    .reset(x400_x7_1_reset),
    .io_a(x400_x7_1_io_a),
    .io_b(x400_x7_1_io_b),
    .io_flow(x400_x7_1_io_flow),
    .io_result(x400_x7_1_io_result)
  );
  RetimeWrapper_232 RetimeWrapper_60 ( // @[package.scala 93:22:@35092.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  x394_x7 x401_sum_1 ( // @[Math.scala 150:24:@35101.4]
    .clock(x401_sum_1_clock),
    .reset(x401_sum_1_reset),
    .io_a(x401_sum_1_io_a),
    .io_b(x401_sum_1_io_b),
    .io_flow(x401_sum_1_io_flow),
    .io_result(x401_sum_1_io_result)
  );
  x402 x402_1 ( // @[Math.scala 720:24:@35111.4]
    .io_b(x402_1_io_b),
    .io_result(x402_1_io_result)
  );
  x403_mul x403_mul_1 ( // @[Math.scala 262:24:@35122.4]
    .clock(x403_mul_1_clock),
    .io_a(x403_mul_1_io_a),
    .io_b(x403_mul_1_io_b),
    .io_flow(x403_mul_1_io_flow),
    .io_result(x403_mul_1_io_result)
  );
  x404 x404_1 ( // @[Math.scala 720:24:@35132.4]
    .io_b(x404_1_io_b),
    .io_result(x404_1_io_result)
  );
  x385 x405_1 ( // @[Math.scala 262:24:@35143.4]
    .clock(x405_1_clock),
    .io_a(x405_1_io_a),
    .io_b(x405_1_io_b),
    .io_flow(x405_1_io_flow),
    .io_result(x405_1_io_result)
  );
  x385 x406_1 ( // @[Math.scala 262:24:@35155.4]
    .clock(x406_1_clock),
    .io_a(x406_1_io_a),
    .io_b(x406_1_io_b),
    .io_flow(x406_1_io_flow),
    .io_result(x406_1_io_result)
  );
  x385 x407_1 ( // @[Math.scala 262:24:@35167.4]
    .clock(x407_1_clock),
    .io_a(x407_1_io_a),
    .io_b(x407_1_io_b),
    .io_flow(x407_1_io_flow),
    .io_result(x407_1_io_result)
  );
  x385 x408_1 ( // @[Math.scala 262:24:@35179.4]
    .clock(x408_1_clock),
    .io_a(x408_1_io_a),
    .io_b(x408_1_io_b),
    .io_flow(x408_1_io_flow),
    .io_result(x408_1_io_result)
  );
  x385 x409_1 ( // @[Math.scala 262:24:@35191.4]
    .clock(x409_1_clock),
    .io_a(x409_1_io_a),
    .io_b(x409_1_io_b),
    .io_flow(x409_1_io_flow),
    .io_result(x409_1_io_result)
  );
  x385 x410_1 ( // @[Math.scala 262:24:@35203.4]
    .clock(x410_1_clock),
    .io_a(x410_1_io_a),
    .io_b(x410_1_io_b),
    .io_flow(x410_1_io_flow),
    .io_result(x410_1_io_result)
  );
  x385 x411_1 ( // @[Math.scala 262:24:@35215.4]
    .clock(x411_1_clock),
    .io_a(x411_1_io_a),
    .io_b(x411_1_io_b),
    .io_flow(x411_1_io_flow),
    .io_result(x411_1_io_result)
  );
  x385 x412_1 ( // @[Math.scala 262:24:@35227.4]
    .clock(x412_1_clock),
    .io_a(x412_1_io_a),
    .io_b(x412_1_io_b),
    .io_flow(x412_1_io_flow),
    .io_result(x412_1_io_result)
  );
  x385 x413_1 ( // @[Math.scala 262:24:@35239.4]
    .clock(x413_1_clock),
    .io_a(x413_1_io_a),
    .io_b(x413_1_io_b),
    .io_flow(x413_1_io_flow),
    .io_result(x413_1_io_result)
  );
  x394_x7 x414_x7_1 ( // @[Math.scala 150:24:@35249.4]
    .clock(x414_x7_1_clock),
    .reset(x414_x7_1_reset),
    .io_a(x414_x7_1_io_a),
    .io_b(x414_x7_1_io_b),
    .io_flow(x414_x7_1_io_flow),
    .io_result(x414_x7_1_io_result)
  );
  x394_x7 x415_x8_1 ( // @[Math.scala 150:24:@35259.4]
    .clock(x415_x8_1_clock),
    .reset(x415_x8_1_reset),
    .io_a(x415_x8_1_io_a),
    .io_b(x415_x8_1_io_b),
    .io_flow(x415_x8_1_io_flow),
    .io_result(x415_x8_1_io_result)
  );
  x394_x7 x416_x7_1 ( // @[Math.scala 150:24:@35269.4]
    .clock(x416_x7_1_clock),
    .reset(x416_x7_1_reset),
    .io_a(x416_x7_1_io_a),
    .io_b(x416_x7_1_io_b),
    .io_flow(x416_x7_1_io_flow),
    .io_result(x416_x7_1_io_result)
  );
  x394_x7 x417_x8_1 ( // @[Math.scala 150:24:@35279.4]
    .clock(x417_x8_1_clock),
    .reset(x417_x8_1_reset),
    .io_a(x417_x8_1_io_a),
    .io_b(x417_x8_1_io_b),
    .io_flow(x417_x8_1_io_flow),
    .io_result(x417_x8_1_io_result)
  );
  x394_x7 x418_x7_1 ( // @[Math.scala 150:24:@35289.4]
    .clock(x418_x7_1_clock),
    .reset(x418_x7_1_reset),
    .io_a(x418_x7_1_io_a),
    .io_b(x418_x7_1_io_b),
    .io_flow(x418_x7_1_io_flow),
    .io_result(x418_x7_1_io_result)
  );
  x394_x7 x419_x8_1 ( // @[Math.scala 150:24:@35299.4]
    .clock(x419_x8_1_clock),
    .reset(x419_x8_1_reset),
    .io_a(x419_x8_1_io_a),
    .io_b(x419_x8_1_io_b),
    .io_flow(x419_x8_1_io_flow),
    .io_result(x419_x8_1_io_result)
  );
  x394_x7 x420_x7_1 ( // @[Math.scala 150:24:@35309.4]
    .clock(x420_x7_1_clock),
    .reset(x420_x7_1_reset),
    .io_a(x420_x7_1_io_a),
    .io_b(x420_x7_1_io_b),
    .io_flow(x420_x7_1_io_flow),
    .io_result(x420_x7_1_io_result)
  );
  RetimeWrapper_232 RetimeWrapper_61 ( // @[package.scala 93:22:@35319.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  x394_x7 x421_sum_1 ( // @[Math.scala 150:24:@35328.4]
    .clock(x421_sum_1_clock),
    .reset(x421_sum_1_reset),
    .io_a(x421_sum_1_io_a),
    .io_b(x421_sum_1_io_b),
    .io_flow(x421_sum_1_io_flow),
    .io_result(x421_sum_1_io_result)
  );
  x402 x422_1 ( // @[Math.scala 720:24:@35338.4]
    .io_b(x422_1_io_b),
    .io_result(x422_1_io_result)
  );
  x403_mul x423_mul_1 ( // @[Math.scala 262:24:@35349.4]
    .clock(x423_mul_1_clock),
    .io_a(x423_mul_1_io_a),
    .io_b(x423_mul_1_io_b),
    .io_flow(x423_mul_1_io_flow),
    .io_result(x423_mul_1_io_result)
  );
  x404 x424_1 ( // @[Math.scala 720:24:@35359.4]
    .io_b(x424_1_io_b),
    .io_result(x424_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_62 ( // @[package.scala 93:22:@35368.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_325 RetimeWrapper_63 ( // @[package.scala 93:22:@35377.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_64 ( // @[package.scala 93:22:@35386.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_65 ( // @[package.scala 93:22:@35395.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_328 RetimeWrapper_66 ( // @[package.scala 93:22:@35404.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_325 RetimeWrapper_67 ( // @[package.scala 93:22:@35413.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_325 RetimeWrapper_68 ( // @[package.scala 93:22:@35424.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_69 ( // @[package.scala 93:22:@35445.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_328 RetimeWrapper_70 ( // @[package.scala 93:22:@35454.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_71 ( // @[package.scala 93:22:@35463.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_325 RetimeWrapper_72 ( // @[package.scala 93:22:@35474.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_73 ( // @[package.scala 93:22:@35495.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_336 RetimeWrapper_74 ( // @[package.scala 93:22:@35504.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_337 RetimeWrapper_75 ( // @[package.scala 93:22:@35513.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_338 RetimeWrapper_76 ( // @[package.scala 93:22:@35522.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_326 RetimeWrapper_77 ( // @[package.scala 93:22:@35531.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_337 RetimeWrapper_78 ( // @[package.scala 93:22:@35540.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_337 RetimeWrapper_79 ( // @[package.scala 93:22:@35552.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_342 RetimeWrapper_80 ( // @[package.scala 93:22:@35573.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_338 RetimeWrapper_81 ( // @[package.scala 93:22:@35582.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_333 RetimeWrapper_82 ( // @[package.scala 93:22:@35591.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_337 RetimeWrapper_83 ( // @[package.scala 93:22:@35603.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_346 RetimeWrapper_84 ( // @[package.scala 93:22:@35624.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_347 RetimeWrapper_85 ( // @[package.scala 93:22:@35633.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_336 RetimeWrapper_86 ( // @[package.scala 93:22:@35642.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_337 RetimeWrapper_87 ( // @[package.scala 93:22:@35654.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_347 RetimeWrapper_88 ( // @[package.scala 93:22:@35675.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_351 RetimeWrapper_89 ( // @[package.scala 93:22:@35684.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_336 RetimeWrapper_90 ( // @[package.scala 93:22:@35693.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_337 RetimeWrapper_91 ( // @[package.scala 93:22:@35705.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_336 RetimeWrapper_92 ( // @[package.scala 93:22:@35726.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_351 RetimeWrapper_93 ( // @[package.scala 93:22:@35735.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_337 RetimeWrapper_94 ( // @[package.scala 93:22:@35747.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_336 RetimeWrapper_95 ( // @[package.scala 93:22:@35768.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_351 RetimeWrapper_96 ( // @[package.scala 93:22:@35777.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_337 RetimeWrapper_97 ( // @[package.scala 93:22:@35789.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  x385 x441_1 ( // @[Math.scala 262:24:@35814.4]
    .clock(x441_1_clock),
    .io_a(x441_1_io_a),
    .io_b(x441_1_io_b),
    .io_flow(x441_1_io_flow),
    .io_result(x441_1_io_result)
  );
  x385 x442_1 ( // @[Math.scala 262:24:@35826.4]
    .clock(x442_1_clock),
    .io_a(x442_1_io_a),
    .io_b(x442_1_io_b),
    .io_flow(x442_1_io_flow),
    .io_result(x442_1_io_result)
  );
  x385 x443_1 ( // @[Math.scala 262:24:@35838.4]
    .clock(x443_1_clock),
    .io_a(x443_1_io_a),
    .io_b(x443_1_io_b),
    .io_flow(x443_1_io_flow),
    .io_result(x443_1_io_result)
  );
  x385 x444_1 ( // @[Math.scala 262:24:@35850.4]
    .clock(x444_1_clock),
    .io_a(x444_1_io_a),
    .io_b(x444_1_io_b),
    .io_flow(x444_1_io_flow),
    .io_result(x444_1_io_result)
  );
  x394_x7 x445_x9_1 ( // @[Math.scala 150:24:@35860.4]
    .clock(x445_x9_1_clock),
    .reset(x445_x9_1_reset),
    .io_a(x445_x9_1_io_a),
    .io_b(x445_x9_1_io_b),
    .io_flow(x445_x9_1_io_flow),
    .io_result(x445_x9_1_io_result)
  );
  x394_x7 x446_x10_1 ( // @[Math.scala 150:24:@35872.4]
    .clock(x446_x10_1_clock),
    .reset(x446_x10_1_reset),
    .io_a(x446_x10_1_io_a),
    .io_b(x446_x10_1_io_b),
    .io_flow(x446_x10_1_io_flow),
    .io_result(x446_x10_1_io_result)
  );
  x394_x7 x447_sum_1 ( // @[Math.scala 150:24:@35882.4]
    .clock(x447_sum_1_clock),
    .reset(x447_sum_1_reset),
    .io_a(x447_sum_1_io_a),
    .io_b(x447_sum_1_io_b),
    .io_flow(x447_sum_1_io_flow),
    .io_result(x447_sum_1_io_result)
  );
  x402 x448_1 ( // @[Math.scala 720:24:@35892.4]
    .io_b(x448_1_io_b),
    .io_result(x448_1_io_result)
  );
  x403_mul x449_mul_1 ( // @[Math.scala 262:24:@35903.4]
    .clock(x449_mul_1_clock),
    .io_a(x449_mul_1_io_a),
    .io_b(x449_mul_1_io_b),
    .io_flow(x449_mul_1_io_flow),
    .io_result(x449_mul_1_io_result)
  );
  x404 x450_1 ( // @[Math.scala 720:24:@35913.4]
    .io_b(x450_1_io_b),
    .io_result(x450_1_io_result)
  );
  x385 x451_1 ( // @[Math.scala 262:24:@35924.4]
    .clock(x451_1_clock),
    .io_a(x451_1_io_a),
    .io_b(x451_1_io_b),
    .io_flow(x451_1_io_flow),
    .io_result(x451_1_io_result)
  );
  x385 x452_1 ( // @[Math.scala 262:24:@35936.4]
    .clock(x452_1_clock),
    .io_a(x452_1_io_a),
    .io_b(x452_1_io_b),
    .io_flow(x452_1_io_flow),
    .io_result(x452_1_io_result)
  );
  x385 x453_1 ( // @[Math.scala 262:24:@35948.4]
    .clock(x453_1_clock),
    .io_a(x453_1_io_a),
    .io_b(x453_1_io_b),
    .io_flow(x453_1_io_flow),
    .io_result(x453_1_io_result)
  );
  x385 x454_1 ( // @[Math.scala 262:24:@35960.4]
    .clock(x454_1_clock),
    .io_a(x454_1_io_a),
    .io_b(x454_1_io_b),
    .io_flow(x454_1_io_flow),
    .io_result(x454_1_io_result)
  );
  x394_x7 x455_x9_1 ( // @[Math.scala 150:24:@35970.4]
    .clock(x455_x9_1_clock),
    .reset(x455_x9_1_reset),
    .io_a(x455_x9_1_io_a),
    .io_b(x455_x9_1_io_b),
    .io_flow(x455_x9_1_io_flow),
    .io_result(x455_x9_1_io_result)
  );
  x394_x7 x456_x10_1 ( // @[Math.scala 150:24:@35980.4]
    .clock(x456_x10_1_clock),
    .reset(x456_x10_1_reset),
    .io_a(x456_x10_1_io_a),
    .io_b(x456_x10_1_io_b),
    .io_flow(x456_x10_1_io_flow),
    .io_result(x456_x10_1_io_result)
  );
  x394_x7 x457_sum_1 ( // @[Math.scala 150:24:@35990.4]
    .clock(x457_sum_1_clock),
    .reset(x457_sum_1_reset),
    .io_a(x457_sum_1_io_a),
    .io_b(x457_sum_1_io_b),
    .io_flow(x457_sum_1_io_flow),
    .io_result(x457_sum_1_io_result)
  );
  x402 x458_1 ( // @[Math.scala 720:24:@36000.4]
    .io_b(x458_1_io_b),
    .io_result(x458_1_io_result)
  );
  x403_mul x459_mul_1 ( // @[Math.scala 262:24:@36011.4]
    .clock(x459_mul_1_clock),
    .io_a(x459_mul_1_io_a),
    .io_b(x459_mul_1_io_b),
    .io_flow(x459_mul_1_io_flow),
    .io_result(x459_mul_1_io_result)
  );
  x404 x460_1 ( // @[Math.scala 720:24:@36021.4]
    .io_b(x460_1_io_b),
    .io_result(x460_1_io_result)
  );
  RetimeWrapper_366 RetimeWrapper_98 ( // @[package.scala 93:22:@36036.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_367 RetimeWrapper_99 ( // @[package.scala 93:22:@36045.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_367 RetimeWrapper_100 ( // @[package.scala 93:22:@36054.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_367 RetimeWrapper_101 ( // @[package.scala 93:22:@36063.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  assign b281 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 62:18:@33392.4]
  assign b282 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 63:18:@33393.4]
  assign _T_205 = b281 & b282; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 67:30:@33395.4]
  assign _T_206 = _T_205 & io_sigsIn_datapathEn; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 67:37:@33396.4]
  assign _T_210 = io_in_x250_TID == 8'h0; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 69:76:@33401.4]
  assign _T_211 = _T_206 & _T_210; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 69:62:@33402.4]
  assign _T_213 = io_in_x250_TDEST == 8'h0; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 69:101:@33403.4]
  assign x543_x283_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@33412.4 package.scala 96:25:@33413.4]
  assign b279_number = __io_result; // @[Math.scala 723:22:@33377.4 Math.scala 724:14:@33378.4]
  assign _T_244 = $signed(b279_number); // @[Math.scala 406:49:@33578.4]
  assign _T_246 = $signed(_T_244) & $signed(32'sh3); // @[Math.scala 406:56:@33580.4]
  assign _T_247 = $signed(_T_246); // @[Math.scala 406:56:@33581.4]
  assign x519_number = $unsigned(_T_247); // @[implicits.scala 133:21:@33582.4]
  assign _T_257 = $signed(x519_number); // @[Math.scala 406:49:@33591.4]
  assign _T_259 = $signed(_T_257) & $signed(32'sh3); // @[Math.scala 406:56:@33593.4]
  assign _T_260 = $signed(_T_259); // @[Math.scala 406:56:@33594.4]
  assign b280_number = __1_io_result; // @[Math.scala 723:22:@33389.4 Math.scala 724:14:@33390.4]
  assign _T_269 = $signed(b280_number); // @[Math.scala 406:49:@33602.4]
  assign _T_271 = $signed(_T_269) & $signed(32'sh3); // @[Math.scala 406:56:@33604.4]
  assign _T_272 = $signed(_T_271); // @[Math.scala 406:56:@33605.4]
  assign _T_276 = x519_number[31]; // @[FixedPoint.scala 50:25:@33611.4]
  assign _T_280 = _T_276 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33613.4]
  assign _T_281 = x519_number[31:2]; // @[FixedPoint.scala 18:52:@33614.4]
  assign _T_287 = _T_281 == 30'h3fffffff; // @[Math.scala 451:55:@33616.4]
  assign _T_288 = x519_number[1:0]; // @[FixedPoint.scala 18:52:@33617.4]
  assign _T_294 = _T_288 != 2'h0; // @[Math.scala 451:110:@33619.4]
  assign _T_295 = _T_287 & _T_294; // @[Math.scala 451:94:@33620.4]
  assign _T_297 = {_T_280,_T_281}; // @[Cat.scala 30:58:@33622.4]
  assign x292_1_number = _T_295 ? 32'h0 : _T_297; // @[Math.scala 454:20:@33623.4]
  assign _GEN_0 = {{9'd0}, x292_1_number}; // @[Math.scala 461:32:@33628.4]
  assign _T_302 = _GEN_0 << 9; // @[Math.scala 461:32:@33628.4]
  assign _GEN_1 = {{5'd0}, x292_1_number}; // @[Math.scala 461:32:@33633.4]
  assign _T_305 = _GEN_1 << 5; // @[Math.scala 461:32:@33633.4]
  assign _T_311 = b280_number[31]; // @[FixedPoint.scala 50:25:@33648.4]
  assign _T_315 = _T_311 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33650.4]
  assign _T_316 = b280_number[31:2]; // @[FixedPoint.scala 18:52:@33651.4]
  assign _T_322 = _T_316 == 30'h3fffffff; // @[Math.scala 451:55:@33653.4]
  assign _T_323 = b280_number[1:0]; // @[FixedPoint.scala 18:52:@33654.4]
  assign _T_329 = _T_323 != 2'h0; // @[Math.scala 451:110:@33656.4]
  assign _T_330 = _T_322 & _T_329; // @[Math.scala 451:94:@33657.4]
  assign _T_332 = {_T_315,_T_316}; // @[Cat.scala 30:58:@33659.4]
  assign _T_360 = ~ io_sigsIn_break; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 118:101:@33736.4]
  assign _T_364 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@33744.4 package.scala 96:25:@33745.4]
  assign _T_366 = io_rr ? _T_364 : 1'h0; // @[implicits.scala 55:10:@33746.4]
  assign _T_367 = _T_360 & _T_366; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 118:118:@33747.4]
  assign _T_369 = _T_367 & _T_360; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 118:206:@33749.4]
  assign _T_370 = _T_369 & io_sigsIn_backpressure; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 118:225:@33750.4]
  assign x546_b281_D3 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@33697.4 package.scala 96:25:@33698.4]
  assign _T_371 = _T_370 & x546_b281_D3; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 118:251:@33751.4]
  assign x550_b282_D3 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@33733.4 package.scala 96:25:@33734.4]
  assign x297_rdcol_number = x297_rdcol_1_io_result; // @[Math.scala 154:22:@33768.4 Math.scala 155:14:@33769.4]
  assign _T_388 = $signed(x297_rdcol_number); // @[Math.scala 406:49:@33777.4]
  assign _T_390 = $signed(_T_388) & $signed(32'sh3); // @[Math.scala 406:56:@33779.4]
  assign _T_391 = $signed(_T_390); // @[Math.scala 406:56:@33780.4]
  assign _T_395 = x297_rdcol_number[31]; // @[FixedPoint.scala 50:25:@33786.4]
  assign _T_399 = _T_395 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@33788.4]
  assign _T_400 = x297_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@33789.4]
  assign _T_406 = _T_400 == 30'h3fffffff; // @[Math.scala 451:55:@33791.4]
  assign _T_407 = x297_rdcol_number[1:0]; // @[FixedPoint.scala 18:52:@33792.4]
  assign _T_413 = _T_407 != 2'h0; // @[Math.scala 451:110:@33794.4]
  assign _T_414 = _T_406 & _T_413; // @[Math.scala 451:94:@33795.4]
  assign _T_416 = {_T_399,_T_400}; // @[Cat.scala 30:58:@33797.4]
  assign _T_436 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@33846.4 package.scala 96:25:@33847.4]
  assign _T_438 = io_rr ? _T_436 : 1'h0; // @[implicits.scala 55:10:@33848.4]
  assign _T_439 = _T_360 & _T_438; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 139:118:@33849.4]
  assign _T_441 = _T_439 & _T_360; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 139:206:@33851.4]
  assign _T_442 = _T_441 & io_sigsIn_backpressure; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 139:225:@33852.4]
  assign _T_443 = _T_442 & x546_b281_D3; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 139:251:@33853.4]
  assign x554_b279_D6_number = RetimeWrapper_13_io_out; // @[package.scala 96:25:@33867.4 package.scala 96:25:@33868.4]
  assign _T_453 = $signed(x554_b279_D6_number); // @[Math.scala 476:37:@33873.4]
  assign x304 = $signed(_T_453) < $signed(32'sh0); // @[Math.scala 476:44:@33875.4]
  assign x555_x297_rdcol_D6_number = RetimeWrapper_14_io_out; // @[package.scala 96:25:@33883.4 package.scala 96:25:@33884.4]
  assign _T_464 = $signed(x555_x297_rdcol_D6_number); // @[Math.scala 476:37:@33889.4]
  assign x305 = $signed(_T_464) < $signed(32'sh0); // @[Math.scala 476:44:@33891.4]
  assign x556_x304_D1 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@33899.4 package.scala 96:25:@33900.4]
  assign x306 = x556_x304_D1 | x305; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 152:24:@33903.4]
  assign _T_503 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@33971.4 package.scala 96:25:@33972.4]
  assign _T_505 = io_rr ? _T_503 : 1'h0; // @[implicits.scala 55:10:@33973.4]
  assign _T_506 = _T_360 & _T_505; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 171:146:@33974.4]
  assign x558_x307_D2 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@33923.4 package.scala 96:25:@33924.4]
  assign _T_507 = _T_506 & x558_x307_D2; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 171:234:@33975.4]
  assign x559_b281_D9 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@33932.4 package.scala 96:25:@33933.4]
  assign _T_508 = _T_507 & x559_b281_D9; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 171:242:@33976.4]
  assign x562_b282_D9 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@33959.4 package.scala 96:25:@33960.4]
  assign x563_b280_D6_number = RetimeWrapper_23_io_out; // @[package.scala 96:25:@33992.4 package.scala 96:25:@33993.4]
  assign _T_521 = $signed(x563_b280_D6_number); // @[Math.scala 476:37:@34000.4]
  assign x310 = $signed(_T_521) < $signed(32'sh0); // @[Math.scala 476:44:@34002.4]
  assign x311 = x304 | x310; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 187:59:@34005.4]
  assign _T_548 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@34046.4 package.scala 96:25:@34047.4]
  assign _T_550 = io_rr ? _T_548 : 1'h0; // @[implicits.scala 55:10:@34048.4]
  assign _T_551 = _T_360 & _T_550; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 200:194:@34049.4]
  assign x564_x312_D3 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@34016.4 package.scala 96:25:@34017.4]
  assign _T_552 = _T_551 & x564_x312_D3; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 200:282:@34050.4]
  assign _T_553 = _T_552 & x559_b281_D9; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 200:290:@34051.4]
  assign x315_rdcol_number = x315_rdcol_1_io_result; // @[Math.scala 154:22:@34070.4 Math.scala 155:14:@34071.4]
  assign _T_568 = $signed(x315_rdcol_number); // @[Math.scala 476:37:@34076.4]
  assign x316 = $signed(_T_568) < $signed(32'sh0); // @[Math.scala 476:44:@34078.4]
  assign x317 = x556_x304_D1 | x316; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 208:59:@34081.4]
  assign _T_584 = $signed(_T_568) & $signed(32'sh3); // @[Math.scala 406:56:@34092.4]
  assign _T_585 = $signed(_T_584); // @[Math.scala 406:56:@34093.4]
  assign _T_589 = x315_rdcol_number[31]; // @[FixedPoint.scala 50:25:@34099.4]
  assign _T_593 = _T_589 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@34101.4]
  assign _T_594 = x315_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@34102.4]
  assign _T_600 = _T_594 == 30'h3fffffff; // @[Math.scala 451:55:@34104.4]
  assign _T_601 = x315_rdcol_number[1:0]; // @[FixedPoint.scala 18:52:@34105.4]
  assign _T_607 = _T_601 != 2'h0; // @[Math.scala 451:110:@34107.4]
  assign _T_608 = _T_600 & _T_607; // @[Math.scala 451:94:@34108.4]
  assign _T_610 = {_T_593,_T_594}; // @[Cat.scala 30:58:@34110.4]
  assign _T_639 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@34169.4 package.scala 96:25:@34170.4]
  assign _T_641 = io_rr ? _T_639 : 1'h0; // @[implicits.scala 55:10:@34171.4]
  assign _T_642 = _T_360 & _T_641; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 229:194:@34172.4]
  assign x570_x318_D2 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@34157.4 package.scala 96:25:@34158.4]
  assign _T_643 = _T_642 & x570_x318_D2; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 229:282:@34173.4]
  assign _T_644 = _T_643 & x559_b281_D9; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 229:290:@34174.4]
  assign x324_rdcol_number = x324_rdcol_1_io_result; // @[Math.scala 154:22:@34193.4 Math.scala 155:14:@34194.4]
  assign _T_659 = $signed(x324_rdcol_number); // @[Math.scala 476:37:@34199.4]
  assign x325 = $signed(_T_659) < $signed(32'sh0); // @[Math.scala 476:44:@34201.4]
  assign x326 = x556_x304_D1 | x325; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 237:59:@34204.4]
  assign _T_675 = $signed(_T_659) & $signed(32'sh3); // @[Math.scala 406:56:@34215.4]
  assign _T_676 = $signed(_T_675); // @[Math.scala 406:56:@34216.4]
  assign _T_680 = x324_rdcol_number[31]; // @[FixedPoint.scala 50:25:@34222.4]
  assign _T_684 = _T_680 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@34224.4]
  assign _T_685 = x324_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@34225.4]
  assign _T_691 = _T_685 == 30'h3fffffff; // @[Math.scala 451:55:@34227.4]
  assign _T_692 = x324_rdcol_number[1:0]; // @[FixedPoint.scala 18:52:@34228.4]
  assign _T_698 = _T_692 != 2'h0; // @[Math.scala 451:110:@34230.4]
  assign _T_699 = _T_691 & _T_698; // @[Math.scala 451:94:@34231.4]
  assign _T_701 = {_T_684,_T_685}; // @[Cat.scala 30:58:@34233.4]
  assign _T_727 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@34283.4 package.scala 96:25:@34284.4]
  assign _T_729 = io_rr ? _T_727 : 1'h0; // @[implicits.scala 55:10:@34285.4]
  assign _T_730 = _T_360 & _T_729; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 256:194:@34286.4]
  assign x573_x327_D2 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@34271.4 package.scala 96:25:@34272.4]
  assign _T_731 = _T_730 & x573_x327_D2; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 256:282:@34287.4]
  assign _T_732 = _T_731 & x559_b281_D9; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 256:290:@34288.4]
  assign x333_rdrow_number = x333_rdrow_1_io_result; // @[Math.scala 195:22:@34307.4 Math.scala 196:14:@34308.4]
  assign _T_749 = $signed(x333_rdrow_number); // @[Math.scala 406:49:@34314.4]
  assign _T_751 = $signed(_T_749) & $signed(32'sh3); // @[Math.scala 406:56:@34316.4]
  assign _T_752 = $signed(_T_751); // @[Math.scala 406:56:@34317.4]
  assign x528_number = $unsigned(_T_752); // @[implicits.scala 133:21:@34318.4]
  assign x335 = $signed(_T_749) < $signed(32'sh0); // @[Math.scala 476:44:@34326.4]
  assign x336 = x335 | x305; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 266:24:@34329.4]
  assign _T_773 = $signed(x528_number); // @[Math.scala 406:49:@34338.4]
  assign _T_775 = $signed(_T_773) & $signed(32'sh3); // @[Math.scala 406:56:@34340.4]
  assign _T_776 = $signed(_T_775); // @[Math.scala 406:56:@34341.4]
  assign _T_780 = x528_number[31]; // @[FixedPoint.scala 50:25:@34347.4]
  assign _T_784 = _T_780 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@34349.4]
  assign _T_785 = x528_number[31:2]; // @[FixedPoint.scala 18:52:@34350.4]
  assign _T_791 = _T_785 == 30'h3fffffff; // @[Math.scala 451:55:@34352.4]
  assign _T_792 = x528_number[1:0]; // @[FixedPoint.scala 18:52:@34353.4]
  assign _T_798 = _T_792 != 2'h0; // @[Math.scala 451:110:@34355.4]
  assign _T_799 = _T_791 & _T_798; // @[Math.scala 451:94:@34356.4]
  assign _T_801 = {_T_784,_T_785}; // @[Cat.scala 30:58:@34358.4]
  assign x339_1_number = _T_799 ? 32'h0 : _T_801; // @[Math.scala 454:20:@34359.4]
  assign _GEN_2 = {{9'd0}, x339_1_number}; // @[Math.scala 461:32:@34364.4]
  assign _T_806 = _GEN_2 << 9; // @[Math.scala 461:32:@34364.4]
  assign _GEN_3 = {{5'd0}, x339_1_number}; // @[Math.scala 461:32:@34369.4]
  assign _T_809 = _GEN_3 << 5; // @[Math.scala 461:32:@34369.4]
  assign _T_836 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@34428.4 package.scala 96:25:@34429.4]
  assign _T_838 = io_rr ? _T_836 : 1'h0; // @[implicits.scala 55:10:@34430.4]
  assign _T_839 = _T_360 & _T_838; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 291:194:@34431.4]
  assign x576_x337_D2 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@34416.4 package.scala 96:25:@34417.4]
  assign _T_840 = _T_839 & x576_x337_D2; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 291:282:@34432.4]
  assign _T_841 = _T_840 & x559_b281_D9; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 291:290:@34433.4]
  assign x577_x310_D1 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@34449.4 package.scala 96:25:@34450.4]
  assign x344 = x335 | x577_x310_D1; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 303:59:@34453.4]
  assign _T_873 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@34497.4 package.scala 96:25:@34498.4]
  assign _T_875 = io_rr ? _T_873 : 1'h0; // @[implicits.scala 55:10:@34499.4]
  assign _T_876 = _T_360 & _T_875; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 318:194:@34500.4]
  assign x579_x345_D2 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@34485.4 package.scala 96:25:@34486.4]
  assign _T_877 = _T_876 & x579_x345_D2; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 318:282:@34501.4]
  assign _T_878 = _T_877 & x559_b281_D9; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 318:290:@34502.4]
  assign x349 = x335 | x316; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 322:59:@34513.4]
  assign _T_905 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@34555.4 package.scala 96:25:@34556.4]
  assign _T_907 = io_rr ? _T_905 : 1'h0; // @[implicits.scala 55:10:@34557.4]
  assign _T_908 = _T_360 & _T_907; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 335:194:@34558.4]
  assign x581_x350_D2 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@34543.4 package.scala 96:25:@34544.4]
  assign _T_909 = _T_908 & x581_x350_D2; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 335:282:@34559.4]
  assign _T_910 = _T_909 & x559_b281_D9; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 335:290:@34560.4]
  assign x354 = x335 | x325; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 339:59:@34571.4]
  assign _T_937 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@34613.4 package.scala 96:25:@34614.4]
  assign _T_939 = io_rr ? _T_937 : 1'h0; // @[implicits.scala 55:10:@34615.4]
  assign _T_940 = _T_360 & _T_939; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 352:194:@34616.4]
  assign x583_x355_D2 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@34601.4 package.scala 96:25:@34602.4]
  assign _T_941 = _T_940 & x583_x355_D2; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 352:282:@34617.4]
  assign _T_942 = _T_941 & x559_b281_D9; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 352:290:@34618.4]
  assign x359_rdrow_number = x359_rdrow_1_io_result; // @[Math.scala 195:22:@34637.4 Math.scala 196:14:@34638.4]
  assign _T_959 = $signed(x359_rdrow_number); // @[Math.scala 406:49:@34644.4]
  assign _T_961 = $signed(_T_959) & $signed(32'sh3); // @[Math.scala 406:56:@34646.4]
  assign _T_962 = $signed(_T_961); // @[Math.scala 406:56:@34647.4]
  assign x533_number = $unsigned(_T_962); // @[implicits.scala 133:21:@34648.4]
  assign x361 = $signed(_T_959) < $signed(32'sh0); // @[Math.scala 476:44:@34656.4]
  assign x362 = x361 | x305; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 362:24:@34659.4]
  assign _T_983 = $signed(x533_number); // @[Math.scala 406:49:@34668.4]
  assign _T_985 = $signed(_T_983) & $signed(32'sh3); // @[Math.scala 406:56:@34670.4]
  assign _T_986 = $signed(_T_985); // @[Math.scala 406:56:@34671.4]
  assign _T_990 = x533_number[31]; // @[FixedPoint.scala 50:25:@34677.4]
  assign _T_994 = _T_990 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@34679.4]
  assign _T_995 = x533_number[31:2]; // @[FixedPoint.scala 18:52:@34680.4]
  assign _T_1001 = _T_995 == 30'h3fffffff; // @[Math.scala 451:55:@34682.4]
  assign _T_1002 = x533_number[1:0]; // @[FixedPoint.scala 18:52:@34683.4]
  assign _T_1008 = _T_1002 != 2'h0; // @[Math.scala 451:110:@34685.4]
  assign _T_1009 = _T_1001 & _T_1008; // @[Math.scala 451:94:@34686.4]
  assign _T_1011 = {_T_994,_T_995}; // @[Cat.scala 30:58:@34688.4]
  assign x365_1_number = _T_1009 ? 32'h0 : _T_1011; // @[Math.scala 454:20:@34689.4]
  assign _GEN_4 = {{9'd0}, x365_1_number}; // @[Math.scala 461:32:@34694.4]
  assign _T_1016 = _GEN_4 << 9; // @[Math.scala 461:32:@34694.4]
  assign _GEN_5 = {{5'd0}, x365_1_number}; // @[Math.scala 461:32:@34699.4]
  assign _T_1019 = _GEN_5 << 5; // @[Math.scala 461:32:@34699.4]
  assign _T_1043 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@34749.4 package.scala 96:25:@34750.4]
  assign _T_1045 = io_rr ? _T_1043 : 1'h0; // @[implicits.scala 55:10:@34751.4]
  assign _T_1046 = _T_360 & _T_1045; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 385:194:@34752.4]
  assign x585_x363_D2 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@34737.4 package.scala 96:25:@34738.4]
  assign _T_1047 = _T_1046 & x585_x363_D2; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 385:282:@34753.4]
  assign _T_1048 = _T_1047 & x559_b281_D9; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 385:290:@34754.4]
  assign x370 = x361 | x577_x310_D1; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 389:24:@34765.4]
  assign _T_1072 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@34798.4 package.scala 96:25:@34799.4]
  assign _T_1074 = io_rr ? _T_1072 : 1'h0; // @[implicits.scala 55:10:@34800.4]
  assign _T_1075 = _T_360 & _T_1074; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 400:194:@34801.4]
  assign x586_x371_D2 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@34786.4 package.scala 96:25:@34787.4]
  assign _T_1076 = _T_1075 & x586_x371_D2; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 400:282:@34802.4]
  assign _T_1077 = _T_1076 & x559_b281_D9; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 400:290:@34803.4]
  assign x375 = x361 | x316; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 404:24:@34814.4]
  assign _T_1101 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@34847.4 package.scala 96:25:@34848.4]
  assign _T_1103 = io_rr ? _T_1101 : 1'h0; // @[implicits.scala 55:10:@34849.4]
  assign _T_1104 = _T_360 & _T_1103; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 415:194:@34850.4]
  assign x587_x376_D2 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@34835.4 package.scala 96:25:@34836.4]
  assign _T_1105 = _T_1104 & x587_x376_D2; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 415:282:@34851.4]
  assign _T_1106 = _T_1105 & x559_b281_D9; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 415:290:@34852.4]
  assign x380 = x361 | x325; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 425:59:@34863.4]
  assign _T_1132 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@34898.4 package.scala 96:25:@34899.4]
  assign _T_1134 = io_rr ? _T_1132 : 1'h0; // @[implicits.scala 55:10:@34900.4]
  assign _T_1135 = _T_360 & _T_1134; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 438:194:@34901.4]
  assign x588_x381_D2 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@34886.4 package.scala 96:25:@34887.4]
  assign _T_1136 = _T_1135 & x588_x381_D2; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 438:282:@34902.4]
  assign _T_1137 = _T_1136 & x559_b281_D9; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 438:290:@34903.4]
  assign _T_1369 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@35429.4 package.scala 96:25:@35430.4]
  assign _T_1371 = io_rr ? _T_1369 : 1'h0; // @[implicits.scala 55:10:@35431.4]
  assign _T_1372 = _T_360 & _T_1371; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 548:167:@35432.4]
  assign _T_1374 = _T_1372 & _T_360; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 548:256:@35434.4]
  assign _T_1375 = _T_1374 & io_sigsIn_backpressure; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 548:275:@35435.4]
  assign x592_b281_D28 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@35382.4 package.scala 96:25:@35383.4]
  assign _T_1376 = _T_1375 & x592_b281_D28; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 548:301:@35436.4]
  assign x596_b282_D28 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@35418.4 package.scala 96:25:@35419.4]
  assign _T_1392 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@35479.4 package.scala 96:25:@35480.4]
  assign _T_1394 = io_rr ? _T_1392 : 1'h0; // @[implicits.scala 55:10:@35481.4]
  assign _T_1395 = _T_360 & _T_1394; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 559:167:@35482.4]
  assign _T_1397 = _T_1395 & _T_360; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 559:256:@35484.4]
  assign _T_1398 = _T_1397 & io_sigsIn_backpressure; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 559:275:@35485.4]
  assign _T_1399 = _T_1398 & x592_b281_D28; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 559:301:@35486.4]
  assign _T_1430 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@35557.4 package.scala 96:25:@35558.4]
  assign _T_1432 = io_rr ? _T_1430 : 1'h0; // @[implicits.scala 55:10:@35559.4]
  assign _T_1433 = _T_360 & _T_1432; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 577:195:@35560.4]
  assign x601_x307_D22 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@35509.4 package.scala 96:25:@35510.4]
  assign _T_1434 = _T_1433 & x601_x307_D22; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 577:284:@35561.4]
  assign x602_b281_D29 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@35518.4 package.scala 96:25:@35519.4]
  assign _T_1435 = _T_1434 & x602_b281_D29; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 577:292:@35562.4]
  assign x605_b282_D29 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@35545.4 package.scala 96:25:@35546.4]
  assign _T_1458 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@35608.4 package.scala 96:25:@35609.4]
  assign _T_1460 = io_rr ? _T_1458 : 1'h0; // @[implicits.scala 55:10:@35610.4]
  assign _T_1461 = _T_360 & _T_1460; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 590:195:@35611.4]
  assign x606_x312_D23 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@35578.4 package.scala 96:25:@35579.4]
  assign _T_1462 = _T_1461 & x606_x312_D23; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 590:284:@35612.4]
  assign _T_1463 = _T_1462 & x602_b281_D29; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 590:292:@35613.4]
  assign _T_1486 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@35659.4 package.scala 96:25:@35660.4]
  assign _T_1488 = io_rr ? _T_1486 : 1'h0; // @[implicits.scala 55:10:@35661.4]
  assign _T_1489 = _T_360 & _T_1488; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 603:195:@35662.4]
  assign x611_x318_D22 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@35647.4 package.scala 96:25:@35648.4]
  assign _T_1490 = _T_1489 & x611_x318_D22; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 603:284:@35663.4]
  assign _T_1491 = _T_1490 & x602_b281_D29; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 603:292:@35664.4]
  assign _T_1514 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@35710.4 package.scala 96:25:@35711.4]
  assign _T_1516 = io_rr ? _T_1514 : 1'h0; // @[implicits.scala 55:10:@35712.4]
  assign _T_1517 = _T_360 & _T_1516; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 616:195:@35713.4]
  assign x614_x337_D22 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@35698.4 package.scala 96:25:@35699.4]
  assign _T_1518 = _T_1517 & x614_x337_D22; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 616:284:@35714.4]
  assign _T_1519 = _T_1518 & x602_b281_D29; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 616:292:@35715.4]
  assign _T_1539 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@35752.4 package.scala 96:25:@35753.4]
  assign _T_1541 = io_rr ? _T_1539 : 1'h0; // @[implicits.scala 55:10:@35754.4]
  assign _T_1542 = _T_360 & _T_1541; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 627:195:@35755.4]
  assign x615_x345_D22 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@35731.4 package.scala 96:25:@35732.4]
  assign _T_1543 = _T_1542 & x615_x345_D22; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 627:284:@35756.4]
  assign _T_1544 = _T_1543 & x602_b281_D29; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 627:292:@35757.4]
  assign _T_1564 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@35794.4 package.scala 96:25:@35795.4]
  assign _T_1566 = io_rr ? _T_1564 : 1'h0; // @[implicits.scala 55:10:@35796.4]
  assign _T_1567 = _T_360 & _T_1566; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 638:195:@35797.4]
  assign x617_x350_D22 = RetimeWrapper_95_io_out; // @[package.scala 96:25:@35773.4 package.scala 96:25:@35774.4]
  assign _T_1568 = _T_1567 & x617_x350_D22; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 638:284:@35798.4]
  assign _T_1569 = _T_1568 & x602_b281_D29; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 638:292:@35799.4]
  assign x450_number = x450_1_io_result; // @[Math.scala 723:22:@35918.4 Math.scala 724:14:@35919.4]
  assign x460_number = x460_1_io_result; // @[Math.scala 723:22:@36026.4 Math.scala 724:14:@36027.4]
  assign _T_1697 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@36068.4 package.scala 96:25:@36069.4]
  assign _T_1699 = io_rr ? _T_1697 : 1'h0; // @[implicits.scala 55:10:@36070.4]
  assign x620_b281_D48 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@36059.4 package.scala 96:25:@36060.4]
  assign _T_1700 = _T_1699 & x620_b281_D48; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 700:117:@36071.4]
  assign x619_b282_D48 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@36050.4 package.scala 96:25:@36051.4]
  assign _T_1701 = _T_1700 & x619_b282_D48; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 700:123:@36072.4]
  assign x547_x520_D3_number = RetimeWrapper_4_io_out; // @[package.scala 96:25:@33706.4 package.scala 96:25:@33707.4]
  assign x548_x521_D3_number = RetimeWrapper_5_io_out; // @[package.scala 96:25:@33715.4 package.scala 96:25:@33716.4]
  assign x549_x295_sum_D1_number = RetimeWrapper_6_io_out; // @[package.scala 96:25:@33724.4 package.scala 96:25:@33725.4]
  assign x551_x301_sum_D1_number = RetimeWrapper_9_io_out; // @[package.scala 96:25:@33817.4 package.scala 96:25:@33818.4]
  assign x553_x525_D2_number = RetimeWrapper_11_io_out; // @[package.scala 96:25:@33835.4 package.scala 96:25:@33836.4]
  assign x557_x301_sum_D7_number = RetimeWrapper_16_io_out; // @[package.scala 96:25:@33914.4 package.scala 96:25:@33915.4]
  assign x560_x520_D9_number = RetimeWrapper_19_io_out; // @[package.scala 96:25:@33941.4 package.scala 96:25:@33942.4]
  assign x561_x525_D8_number = RetimeWrapper_20_io_out; // @[package.scala 96:25:@33950.4 package.scala 96:25:@33951.4]
  assign x565_x521_D9_number = RetimeWrapper_25_io_out; // @[package.scala 96:25:@34025.4 package.scala 96:25:@34026.4]
  assign x566_x295_sum_D7_number = RetimeWrapper_26_io_out; // @[package.scala 96:25:@34034.4 package.scala 96:25:@34035.4]
  assign x568_x321_sum_D1_number = RetimeWrapper_29_io_out; // @[package.scala 96:25:@34139.4 package.scala 96:25:@34140.4]
  assign x569_x526_D2_number = RetimeWrapper_30_io_out; // @[package.scala 96:25:@34148.4 package.scala 96:25:@34149.4]
  assign x571_x527_D2_number = RetimeWrapper_33_io_out; // @[package.scala 96:25:@34253.4 package.scala 96:25:@34254.4]
  assign x572_x330_sum_D1_number = RetimeWrapper_34_io_out; // @[package.scala 96:25:@34262.4 package.scala 96:25:@34263.4]
  assign x341_sum_number = x341_sum_1_io_result; // @[Math.scala 154:22:@34398.4 Math.scala 155:14:@34399.4]
  assign x575_x529_D2_number = RetimeWrapper_38_io_out; // @[package.scala 96:25:@34407.4 package.scala 96:25:@34408.4]
  assign x346_sum_number = x346_sum_1_io_result; // @[Math.scala 154:22:@34476.4 Math.scala 155:14:@34477.4]
  assign x351_sum_number = x351_sum_1_io_result; // @[Math.scala 154:22:@34534.4 Math.scala 155:14:@34535.4]
  assign x356_sum_number = x356_sum_1_io_result; // @[Math.scala 154:22:@34592.4 Math.scala 155:14:@34593.4]
  assign x367_sum_number = x367_sum_1_io_result; // @[Math.scala 154:22:@34719.4 Math.scala 155:14:@34720.4]
  assign x584_x534_D2_number = RetimeWrapper_51_io_out; // @[package.scala 96:25:@34728.4 package.scala 96:25:@34729.4]
  assign x372_sum_number = x372_sum_1_io_result; // @[Math.scala 154:22:@34777.4 Math.scala 155:14:@34778.4]
  assign x377_sum_number = x377_sum_1_io_result; // @[Math.scala 154:22:@34826.4 Math.scala 155:14:@34827.4]
  assign x382_sum_number = x382_sum_1_io_result; // @[Math.scala 154:22:@34877.4 Math.scala 155:14:@34878.4]
  assign x593_x520_D28_number = RetimeWrapper_64_io_out; // @[package.scala 96:25:@35391.4 package.scala 96:25:@35392.4]
  assign x594_x521_D28_number = RetimeWrapper_65_io_out; // @[package.scala 96:25:@35400.4 package.scala 96:25:@35401.4]
  assign x595_x295_sum_D26_number = RetimeWrapper_66_io_out; // @[package.scala 96:25:@35409.4 package.scala 96:25:@35410.4]
  assign x598_x301_sum_D26_number = RetimeWrapper_70_io_out; // @[package.scala 96:25:@35459.4 package.scala 96:25:@35460.4]
  assign x599_x525_D27_number = RetimeWrapper_71_io_out; // @[package.scala 96:25:@35468.4 package.scala 96:25:@35469.4]
  assign x600_x301_sum_D27_number = RetimeWrapper_73_io_out; // @[package.scala 96:25:@35500.4 package.scala 96:25:@35501.4]
  assign x603_x520_D29_number = RetimeWrapper_76_io_out; // @[package.scala 96:25:@35527.4 package.scala 96:25:@35528.4]
  assign x604_x525_D28_number = RetimeWrapper_77_io_out; // @[package.scala 96:25:@35536.4 package.scala 96:25:@35537.4]
  assign x607_x521_D29_number = RetimeWrapper_81_io_out; // @[package.scala 96:25:@35587.4 package.scala 96:25:@35588.4]
  assign x608_x295_sum_D27_number = RetimeWrapper_82_io_out; // @[package.scala 96:25:@35596.4 package.scala 96:25:@35597.4]
  assign x609_x321_sum_D21_number = RetimeWrapper_84_io_out; // @[package.scala 96:25:@35629.4 package.scala 96:25:@35630.4]
  assign x610_x526_D22_number = RetimeWrapper_85_io_out; // @[package.scala 96:25:@35638.4 package.scala 96:25:@35639.4]
  assign x612_x529_D22_number = RetimeWrapper_88_io_out; // @[package.scala 96:25:@35680.4 package.scala 96:25:@35681.4]
  assign x613_x341_sum_D20_number = RetimeWrapper_89_io_out; // @[package.scala 96:25:@35689.4 package.scala 96:25:@35690.4]
  assign x616_x346_sum_D20_number = RetimeWrapper_93_io_out; // @[package.scala 96:25:@35740.4 package.scala 96:25:@35741.4]
  assign x618_x351_sum_D20_number = RetimeWrapper_96_io_out; // @[package.scala 96:25:@35782.4 package.scala 96:25:@35783.4]
  assign io_in_x251_TVALID = _T_1701 & io_sigsIn_backpressure; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 700:22:@36074.4]
  assign io_in_x251_TDATA = {{192'd0}, RetimeWrapper_98_io_out}; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 701:24:@36075.4]
  assign io_in_x250_TREADY = _T_211 & _T_213; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 67:22:@33397.4 sm_x465_inr_Foreach_SAMPLER_BOX.scala 69:22:@33405.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@33375.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@33387.4]
  assign RetimeWrapper_clock = clock; // @[:@33408.4]
  assign RetimeWrapper_reset = reset; // @[:@33409.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33411.4]
  assign RetimeWrapper_io_in = io_in_x250_TDATA[63:0]; // @[package.scala 94:16:@33410.4]
  assign x285_lb_0_clock = clock; // @[:@33418.4]
  assign x285_lb_0_reset = reset; // @[:@33419.4]
  assign x285_lb_0_io_rPort_11_banks_1 = x569_x526_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34177.4]
  assign x285_lb_0_io_rPort_11_banks_0 = x560_x520_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@34176.4]
  assign x285_lb_0_io_rPort_11_ofs_0 = x568_x321_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@34178.4]
  assign x285_lb_0_io_rPort_11_en_0 = _T_644 & x562_b282_D9; // @[MemInterfaceType.scala 110:79:@34180.4]
  assign x285_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34179.4]
  assign x285_lb_0_io_rPort_10_banks_1 = x565_x521_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@34806.4]
  assign x285_lb_0_io_rPort_10_banks_0 = x584_x534_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34805.4]
  assign x285_lb_0_io_rPort_10_ofs_0 = x372_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@34807.4]
  assign x285_lb_0_io_rPort_10_en_0 = _T_1077 & x562_b282_D9; // @[MemInterfaceType.scala 110:79:@34809.4]
  assign x285_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34808.4]
  assign x285_lb_0_io_rPort_9_banks_1 = x571_x527_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34906.4]
  assign x285_lb_0_io_rPort_9_banks_0 = x584_x534_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34905.4]
  assign x285_lb_0_io_rPort_9_ofs_0 = x382_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@34907.4]
  assign x285_lb_0_io_rPort_9_en_0 = _T_1137 & x562_b282_D9; // @[MemInterfaceType.scala 110:79:@34909.4]
  assign x285_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34908.4]
  assign x285_lb_0_io_rPort_8_banks_1 = x569_x526_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34855.4]
  assign x285_lb_0_io_rPort_8_banks_0 = x584_x534_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34854.4]
  assign x285_lb_0_io_rPort_8_ofs_0 = x377_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@34856.4]
  assign x285_lb_0_io_rPort_8_en_0 = _T_1106 & x562_b282_D9; // @[MemInterfaceType.scala 110:79:@34858.4]
  assign x285_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34857.4]
  assign x285_lb_0_io_rPort_7_banks_1 = x561_x525_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@34757.4]
  assign x285_lb_0_io_rPort_7_banks_0 = x584_x534_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34756.4]
  assign x285_lb_0_io_rPort_7_ofs_0 = x367_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@34758.4]
  assign x285_lb_0_io_rPort_7_en_0 = _T_1048 & x562_b282_D9; // @[MemInterfaceType.scala 110:79:@34760.4]
  assign x285_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34759.4]
  assign x285_lb_0_io_rPort_6_banks_1 = x571_x527_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34291.4]
  assign x285_lb_0_io_rPort_6_banks_0 = x560_x520_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@34290.4]
  assign x285_lb_0_io_rPort_6_ofs_0 = x572_x330_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@34292.4]
  assign x285_lb_0_io_rPort_6_en_0 = _T_732 & x562_b282_D9; // @[MemInterfaceType.scala 110:79:@34294.4]
  assign x285_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34293.4]
  assign x285_lb_0_io_rPort_5_banks_1 = x561_x525_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@34436.4]
  assign x285_lb_0_io_rPort_5_banks_0 = x575_x529_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34435.4]
  assign x285_lb_0_io_rPort_5_ofs_0 = x341_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@34437.4]
  assign x285_lb_0_io_rPort_5_en_0 = _T_841 & x562_b282_D9; // @[MemInterfaceType.scala 110:79:@34439.4]
  assign x285_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34438.4]
  assign x285_lb_0_io_rPort_4_banks_1 = x565_x521_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@34054.4]
  assign x285_lb_0_io_rPort_4_banks_0 = x560_x520_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@34053.4]
  assign x285_lb_0_io_rPort_4_ofs_0 = x566_x295_sum_D7_number[8:0]; // @[MemInterfaceType.scala 107:54:@34055.4]
  assign x285_lb_0_io_rPort_4_en_0 = _T_553 & x562_b282_D9; // @[MemInterfaceType.scala 110:79:@34057.4]
  assign x285_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34056.4]
  assign x285_lb_0_io_rPort_3_banks_1 = x571_x527_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34621.4]
  assign x285_lb_0_io_rPort_3_banks_0 = x575_x529_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34620.4]
  assign x285_lb_0_io_rPort_3_ofs_0 = x356_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@34622.4]
  assign x285_lb_0_io_rPort_3_en_0 = _T_942 & x562_b282_D9; // @[MemInterfaceType.scala 110:79:@34624.4]
  assign x285_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34623.4]
  assign x285_lb_0_io_rPort_2_banks_1 = x561_x525_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@33979.4]
  assign x285_lb_0_io_rPort_2_banks_0 = x560_x520_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@33978.4]
  assign x285_lb_0_io_rPort_2_ofs_0 = x557_x301_sum_D7_number[8:0]; // @[MemInterfaceType.scala 107:54:@33980.4]
  assign x285_lb_0_io_rPort_2_en_0 = _T_508 & x562_b282_D9; // @[MemInterfaceType.scala 110:79:@33982.4]
  assign x285_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@33981.4]
  assign x285_lb_0_io_rPort_1_banks_1 = x569_x526_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34563.4]
  assign x285_lb_0_io_rPort_1_banks_0 = x575_x529_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34562.4]
  assign x285_lb_0_io_rPort_1_ofs_0 = x351_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@34564.4]
  assign x285_lb_0_io_rPort_1_en_0 = _T_910 & x562_b282_D9; // @[MemInterfaceType.scala 110:79:@34566.4]
  assign x285_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34565.4]
  assign x285_lb_0_io_rPort_0_banks_1 = x565_x521_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@34505.4]
  assign x285_lb_0_io_rPort_0_banks_0 = x575_x529_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@34504.4]
  assign x285_lb_0_io_rPort_0_ofs_0 = x346_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@34506.4]
  assign x285_lb_0_io_rPort_0_en_0 = _T_878 & x562_b282_D9; // @[MemInterfaceType.scala 110:79:@34508.4]
  assign x285_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@34507.4]
  assign x285_lb_0_io_wPort_1_banks_1 = x553_x525_D2_number[2:0]; // @[MemInterfaceType.scala 88:58:@33856.4]
  assign x285_lb_0_io_wPort_1_banks_0 = x547_x520_D3_number[2:0]; // @[MemInterfaceType.scala 88:58:@33855.4]
  assign x285_lb_0_io_wPort_1_ofs_0 = x551_x301_sum_D1_number[8:0]; // @[MemInterfaceType.scala 89:54:@33857.4]
  assign x285_lb_0_io_wPort_1_data_0 = RetimeWrapper_10_io_out; // @[MemInterfaceType.scala 90:56:@33858.4]
  assign x285_lb_0_io_wPort_1_en_0 = _T_443 & x550_b282_D3; // @[MemInterfaceType.scala 93:57:@33860.4]
  assign x285_lb_0_io_wPort_0_banks_1 = x548_x521_D3_number[2:0]; // @[MemInterfaceType.scala 88:58:@33754.4]
  assign x285_lb_0_io_wPort_0_banks_0 = x547_x520_D3_number[2:0]; // @[MemInterfaceType.scala 88:58:@33753.4]
  assign x285_lb_0_io_wPort_0_ofs_0 = x549_x295_sum_D1_number[8:0]; // @[MemInterfaceType.scala 89:54:@33755.4]
  assign x285_lb_0_io_wPort_0_data_0 = RetimeWrapper_2_io_out; // @[MemInterfaceType.scala 90:56:@33756.4]
  assign x285_lb_0_io_wPort_0_en_0 = _T_371 & x550_b282_D3; // @[MemInterfaceType.scala 93:57:@33758.4]
  assign x286_lb2_0_clock = clock; // @[:@33511.4]
  assign x286_lb2_0_reset = reset; // @[:@33512.4]
  assign x286_lb2_0_io_rPort_5_banks_1 = x607_x521_D29_number[2:0]; // @[MemInterfaceType.scala 106:58:@35760.4]
  assign x286_lb2_0_io_rPort_5_banks_0 = x612_x529_D22_number[2:0]; // @[MemInterfaceType.scala 106:58:@35759.4]
  assign x286_lb2_0_io_rPort_5_ofs_0 = x616_x346_sum_D20_number[8:0]; // @[MemInterfaceType.scala 107:54:@35761.4]
  assign x286_lb2_0_io_rPort_5_en_0 = _T_1544 & x605_b282_D29; // @[MemInterfaceType.scala 110:79:@35763.4]
  assign x286_lb2_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35762.4]
  assign x286_lb2_0_io_rPort_4_banks_1 = x610_x526_D22_number[2:0]; // @[MemInterfaceType.scala 106:58:@35667.4]
  assign x286_lb2_0_io_rPort_4_banks_0 = x603_x520_D29_number[2:0]; // @[MemInterfaceType.scala 106:58:@35666.4]
  assign x286_lb2_0_io_rPort_4_ofs_0 = x609_x321_sum_D21_number[8:0]; // @[MemInterfaceType.scala 107:54:@35668.4]
  assign x286_lb2_0_io_rPort_4_en_0 = _T_1491 & x605_b282_D29; // @[MemInterfaceType.scala 110:79:@35670.4]
  assign x286_lb2_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35669.4]
  assign x286_lb2_0_io_rPort_3_banks_1 = x607_x521_D29_number[2:0]; // @[MemInterfaceType.scala 106:58:@35616.4]
  assign x286_lb2_0_io_rPort_3_banks_0 = x603_x520_D29_number[2:0]; // @[MemInterfaceType.scala 106:58:@35615.4]
  assign x286_lb2_0_io_rPort_3_ofs_0 = x608_x295_sum_D27_number[8:0]; // @[MemInterfaceType.scala 107:54:@35617.4]
  assign x286_lb2_0_io_rPort_3_en_0 = _T_1463 & x605_b282_D29; // @[MemInterfaceType.scala 110:79:@35619.4]
  assign x286_lb2_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35618.4]
  assign x286_lb2_0_io_rPort_2_banks_1 = x604_x525_D28_number[2:0]; // @[MemInterfaceType.scala 106:58:@35718.4]
  assign x286_lb2_0_io_rPort_2_banks_0 = x612_x529_D22_number[2:0]; // @[MemInterfaceType.scala 106:58:@35717.4]
  assign x286_lb2_0_io_rPort_2_ofs_0 = x613_x341_sum_D20_number[8:0]; // @[MemInterfaceType.scala 107:54:@35719.4]
  assign x286_lb2_0_io_rPort_2_en_0 = _T_1519 & x605_b282_D29; // @[MemInterfaceType.scala 110:79:@35721.4]
  assign x286_lb2_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35720.4]
  assign x286_lb2_0_io_rPort_1_banks_1 = x604_x525_D28_number[2:0]; // @[MemInterfaceType.scala 106:58:@35565.4]
  assign x286_lb2_0_io_rPort_1_banks_0 = x603_x520_D29_number[2:0]; // @[MemInterfaceType.scala 106:58:@35564.4]
  assign x286_lb2_0_io_rPort_1_ofs_0 = x600_x301_sum_D27_number[8:0]; // @[MemInterfaceType.scala 107:54:@35566.4]
  assign x286_lb2_0_io_rPort_1_en_0 = _T_1435 & x605_b282_D29; // @[MemInterfaceType.scala 110:79:@35568.4]
  assign x286_lb2_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35567.4]
  assign x286_lb2_0_io_rPort_0_banks_1 = x610_x526_D22_number[2:0]; // @[MemInterfaceType.scala 106:58:@35802.4]
  assign x286_lb2_0_io_rPort_0_banks_0 = x612_x529_D22_number[2:0]; // @[MemInterfaceType.scala 106:58:@35801.4]
  assign x286_lb2_0_io_rPort_0_ofs_0 = x618_x351_sum_D20_number[8:0]; // @[MemInterfaceType.scala 107:54:@35803.4]
  assign x286_lb2_0_io_rPort_0_en_0 = _T_1569 & x605_b282_D29; // @[MemInterfaceType.scala 110:79:@35805.4]
  assign x286_lb2_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@35804.4]
  assign x286_lb2_0_io_wPort_1_banks_1 = x599_x525_D27_number[2:0]; // @[MemInterfaceType.scala 88:58:@35489.4]
  assign x286_lb2_0_io_wPort_1_banks_0 = x593_x520_D28_number[2:0]; // @[MemInterfaceType.scala 88:58:@35488.4]
  assign x286_lb2_0_io_wPort_1_ofs_0 = x598_x301_sum_D26_number[8:0]; // @[MemInterfaceType.scala 89:54:@35490.4]
  assign x286_lb2_0_io_wPort_1_data_0 = RetimeWrapper_69_io_out; // @[MemInterfaceType.scala 90:56:@35491.4]
  assign x286_lb2_0_io_wPort_1_en_0 = _T_1399 & x596_b282_D28; // @[MemInterfaceType.scala 93:57:@35493.4]
  assign x286_lb2_0_io_wPort_0_banks_1 = x594_x521_D28_number[2:0]; // @[MemInterfaceType.scala 88:58:@35439.4]
  assign x286_lb2_0_io_wPort_0_banks_0 = x593_x520_D28_number[2:0]; // @[MemInterfaceType.scala 88:58:@35438.4]
  assign x286_lb2_0_io_wPort_0_ofs_0 = x595_x295_sum_D26_number[8:0]; // @[MemInterfaceType.scala 89:54:@35440.4]
  assign x286_lb2_0_io_wPort_0_data_0 = RetimeWrapper_62_io_out; // @[MemInterfaceType.scala 90:56:@35441.4]
  assign x286_lb2_0_io_wPort_0_en_0 = _T_1376 & x596_b282_D28; // @[MemInterfaceType.scala 93:57:@35443.4]
  assign x524_sub_1_clock = clock; // @[:@33638.4]
  assign x524_sub_1_reset = reset; // @[:@33639.4]
  assign x524_sub_1_io_a = _T_302[31:0]; // @[Math.scala 192:17:@33640.4]
  assign x524_sub_1_io_b = _T_305[31:0]; // @[Math.scala 193:17:@33641.4]
  assign x524_sub_1_io_flow = io_in_x251_TREADY; // @[Math.scala 194:20:@33642.4]
  assign RetimeWrapper_1_clock = clock; // @[:@33665.4]
  assign RetimeWrapper_1_reset = reset; // @[:@33666.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33668.4]
  assign RetimeWrapper_1_io_in = _T_330 ? 32'h0 : _T_332; // @[package.scala 94:16:@33667.4]
  assign x295_sum_1_clock = clock; // @[:@33674.4]
  assign x295_sum_1_reset = reset; // @[:@33675.4]
  assign x295_sum_1_io_a = x524_sub_1_io_result; // @[Math.scala 151:17:@33676.4]
  assign x295_sum_1_io_b = RetimeWrapper_1_io_out; // @[Math.scala 152:17:@33677.4]
  assign x295_sum_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@33678.4]
  assign RetimeWrapper_2_clock = clock; // @[:@33684.4]
  assign RetimeWrapper_2_reset = reset; // @[:@33685.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33687.4]
  assign RetimeWrapper_2_io_in = x543_x283_D1_0_number[31:0]; // @[package.scala 94:16:@33686.4]
  assign RetimeWrapper_3_clock = clock; // @[:@33693.4]
  assign RetimeWrapper_3_reset = reset; // @[:@33694.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33696.4]
  assign RetimeWrapper_3_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@33695.4]
  assign RetimeWrapper_4_clock = clock; // @[:@33702.4]
  assign RetimeWrapper_4_reset = reset; // @[:@33703.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33705.4]
  assign RetimeWrapper_4_io_in = $unsigned(_T_260); // @[package.scala 94:16:@33704.4]
  assign RetimeWrapper_5_clock = clock; // @[:@33711.4]
  assign RetimeWrapper_5_reset = reset; // @[:@33712.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33714.4]
  assign RetimeWrapper_5_io_in = $unsigned(_T_272); // @[package.scala 94:16:@33713.4]
  assign RetimeWrapper_6_clock = clock; // @[:@33720.4]
  assign RetimeWrapper_6_reset = reset; // @[:@33721.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33723.4]
  assign RetimeWrapper_6_io_in = x295_sum_1_io_result; // @[package.scala 94:16:@33722.4]
  assign RetimeWrapper_7_clock = clock; // @[:@33729.4]
  assign RetimeWrapper_7_reset = reset; // @[:@33730.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33732.4]
  assign RetimeWrapper_7_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@33731.4]
  assign RetimeWrapper_8_clock = clock; // @[:@33740.4]
  assign RetimeWrapper_8_reset = reset; // @[:@33741.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33743.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33742.4]
  assign x297_rdcol_1_clock = clock; // @[:@33763.4]
  assign x297_rdcol_1_reset = reset; // @[:@33764.4]
  assign x297_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@33765.4]
  assign x297_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@33766.4]
  assign x297_rdcol_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@33767.4]
  assign x301_sum_1_clock = clock; // @[:@33803.4]
  assign x301_sum_1_reset = reset; // @[:@33804.4]
  assign x301_sum_1_io_a = x524_sub_1_io_result; // @[Math.scala 151:17:@33805.4]
  assign x301_sum_1_io_b = _T_414 ? 32'h0 : _T_416; // @[Math.scala 152:17:@33806.4]
  assign x301_sum_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@33807.4]
  assign RetimeWrapper_9_clock = clock; // @[:@33813.4]
  assign RetimeWrapper_9_reset = reset; // @[:@33814.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33816.4]
  assign RetimeWrapper_9_io_in = x301_sum_1_io_result; // @[package.scala 94:16:@33815.4]
  assign RetimeWrapper_10_clock = clock; // @[:@33822.4]
  assign RetimeWrapper_10_reset = reset; // @[:@33823.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33825.4]
  assign RetimeWrapper_10_io_in = x543_x283_D1_0_number[63:32]; // @[package.scala 94:16:@33824.4]
  assign RetimeWrapper_11_clock = clock; // @[:@33831.4]
  assign RetimeWrapper_11_reset = reset; // @[:@33832.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33834.4]
  assign RetimeWrapper_11_io_in = $unsigned(_T_391); // @[package.scala 94:16:@33833.4]
  assign RetimeWrapper_12_clock = clock; // @[:@33842.4]
  assign RetimeWrapper_12_reset = reset; // @[:@33843.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33845.4]
  assign RetimeWrapper_12_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33844.4]
  assign RetimeWrapper_13_clock = clock; // @[:@33863.4]
  assign RetimeWrapper_13_reset = reset; // @[:@33864.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33866.4]
  assign RetimeWrapper_13_io_in = __io_result; // @[package.scala 94:16:@33865.4]
  assign RetimeWrapper_14_clock = clock; // @[:@33879.4]
  assign RetimeWrapper_14_reset = reset; // @[:@33880.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33882.4]
  assign RetimeWrapper_14_io_in = x297_rdcol_1_io_result; // @[package.scala 94:16:@33881.4]
  assign RetimeWrapper_15_clock = clock; // @[:@33895.4]
  assign RetimeWrapper_15_reset = reset; // @[:@33896.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33898.4]
  assign RetimeWrapper_15_io_in = $signed(_T_453) < $signed(32'sh0); // @[package.scala 94:16:@33897.4]
  assign RetimeWrapper_16_clock = clock; // @[:@33910.4]
  assign RetimeWrapper_16_reset = reset; // @[:@33911.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33913.4]
  assign RetimeWrapper_16_io_in = x301_sum_1_io_result; // @[package.scala 94:16:@33912.4]
  assign RetimeWrapper_17_clock = clock; // @[:@33919.4]
  assign RetimeWrapper_17_reset = reset; // @[:@33920.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33922.4]
  assign RetimeWrapper_17_io_in = ~ x306; // @[package.scala 94:16:@33921.4]
  assign RetimeWrapper_18_clock = clock; // @[:@33928.4]
  assign RetimeWrapper_18_reset = reset; // @[:@33929.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33931.4]
  assign RetimeWrapper_18_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@33930.4]
  assign RetimeWrapper_19_clock = clock; // @[:@33937.4]
  assign RetimeWrapper_19_reset = reset; // @[:@33938.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33940.4]
  assign RetimeWrapper_19_io_in = $unsigned(_T_260); // @[package.scala 94:16:@33939.4]
  assign RetimeWrapper_20_clock = clock; // @[:@33946.4]
  assign RetimeWrapper_20_reset = reset; // @[:@33947.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33949.4]
  assign RetimeWrapper_20_io_in = $unsigned(_T_391); // @[package.scala 94:16:@33948.4]
  assign RetimeWrapper_21_clock = clock; // @[:@33955.4]
  assign RetimeWrapper_21_reset = reset; // @[:@33956.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33958.4]
  assign RetimeWrapper_21_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@33957.4]
  assign RetimeWrapper_22_clock = clock; // @[:@33967.4]
  assign RetimeWrapper_22_reset = reset; // @[:@33968.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33970.4]
  assign RetimeWrapper_22_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@33969.4]
  assign RetimeWrapper_23_clock = clock; // @[:@33988.4]
  assign RetimeWrapper_23_reset = reset; // @[:@33989.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@33991.4]
  assign RetimeWrapper_23_io_in = __1_io_result; // @[package.scala 94:16:@33990.4]
  assign RetimeWrapper_24_clock = clock; // @[:@34012.4]
  assign RetimeWrapper_24_reset = reset; // @[:@34013.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34015.4]
  assign RetimeWrapper_24_io_in = ~ x311; // @[package.scala 94:16:@34014.4]
  assign RetimeWrapper_25_clock = clock; // @[:@34021.4]
  assign RetimeWrapper_25_reset = reset; // @[:@34022.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34024.4]
  assign RetimeWrapper_25_io_in = $unsigned(_T_272); // @[package.scala 94:16:@34023.4]
  assign RetimeWrapper_26_clock = clock; // @[:@34030.4]
  assign RetimeWrapper_26_reset = reset; // @[:@34031.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34033.4]
  assign RetimeWrapper_26_io_in = x295_sum_1_io_result; // @[package.scala 94:16:@34032.4]
  assign RetimeWrapper_27_clock = clock; // @[:@34042.4]
  assign RetimeWrapper_27_reset = reset; // @[:@34043.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34045.4]
  assign RetimeWrapper_27_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34044.4]
  assign x315_rdcol_1_clock = clock; // @[:@34065.4]
  assign x315_rdcol_1_reset = reset; // @[:@34066.4]
  assign x315_rdcol_1_io_a = RetimeWrapper_23_io_out; // @[Math.scala 151:17:@34067.4]
  assign x315_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@34068.4]
  assign x315_rdcol_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@34069.4]
  assign RetimeWrapper_28_clock = clock; // @[:@34116.4]
  assign RetimeWrapper_28_reset = reset; // @[:@34117.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34119.4]
  assign RetimeWrapper_28_io_in = x524_sub_1_io_result; // @[package.scala 94:16:@34118.4]
  assign x321_sum_1_clock = clock; // @[:@34125.4]
  assign x321_sum_1_reset = reset; // @[:@34126.4]
  assign x321_sum_1_io_a = RetimeWrapper_28_io_out; // @[Math.scala 151:17:@34127.4]
  assign x321_sum_1_io_b = _T_608 ? 32'h0 : _T_610; // @[Math.scala 152:17:@34128.4]
  assign x321_sum_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@34129.4]
  assign RetimeWrapper_29_clock = clock; // @[:@34135.4]
  assign RetimeWrapper_29_reset = reset; // @[:@34136.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34138.4]
  assign RetimeWrapper_29_io_in = x321_sum_1_io_result; // @[package.scala 94:16:@34137.4]
  assign RetimeWrapper_30_clock = clock; // @[:@34144.4]
  assign RetimeWrapper_30_reset = reset; // @[:@34145.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34147.4]
  assign RetimeWrapper_30_io_in = $unsigned(_T_585); // @[package.scala 94:16:@34146.4]
  assign RetimeWrapper_31_clock = clock; // @[:@34153.4]
  assign RetimeWrapper_31_reset = reset; // @[:@34154.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34156.4]
  assign RetimeWrapper_31_io_in = ~ x317; // @[package.scala 94:16:@34155.4]
  assign RetimeWrapper_32_clock = clock; // @[:@34165.4]
  assign RetimeWrapper_32_reset = reset; // @[:@34166.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34168.4]
  assign RetimeWrapper_32_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34167.4]
  assign x324_rdcol_1_clock = clock; // @[:@34188.4]
  assign x324_rdcol_1_reset = reset; // @[:@34189.4]
  assign x324_rdcol_1_io_a = RetimeWrapper_23_io_out; // @[Math.scala 151:17:@34190.4]
  assign x324_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@34191.4]
  assign x324_rdcol_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@34192.4]
  assign x330_sum_1_clock = clock; // @[:@34239.4]
  assign x330_sum_1_reset = reset; // @[:@34240.4]
  assign x330_sum_1_io_a = RetimeWrapper_28_io_out; // @[Math.scala 151:17:@34241.4]
  assign x330_sum_1_io_b = _T_699 ? 32'h0 : _T_701; // @[Math.scala 152:17:@34242.4]
  assign x330_sum_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@34243.4]
  assign RetimeWrapper_33_clock = clock; // @[:@34249.4]
  assign RetimeWrapper_33_reset = reset; // @[:@34250.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34252.4]
  assign RetimeWrapper_33_io_in = $unsigned(_T_676); // @[package.scala 94:16:@34251.4]
  assign RetimeWrapper_34_clock = clock; // @[:@34258.4]
  assign RetimeWrapper_34_reset = reset; // @[:@34259.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34261.4]
  assign RetimeWrapper_34_io_in = x330_sum_1_io_result; // @[package.scala 94:16:@34260.4]
  assign RetimeWrapper_35_clock = clock; // @[:@34267.4]
  assign RetimeWrapper_35_reset = reset; // @[:@34268.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34270.4]
  assign RetimeWrapper_35_io_in = ~ x326; // @[package.scala 94:16:@34269.4]
  assign RetimeWrapper_36_clock = clock; // @[:@34279.4]
  assign RetimeWrapper_36_reset = reset; // @[:@34280.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34282.4]
  assign RetimeWrapper_36_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34281.4]
  assign x333_rdrow_1_clock = clock; // @[:@34302.4]
  assign x333_rdrow_1_reset = reset; // @[:@34303.4]
  assign x333_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@34304.4]
  assign x333_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@34305.4]
  assign x333_rdrow_1_io_flow = io_in_x251_TREADY; // @[Math.scala 194:20:@34306.4]
  assign x532_sub_1_clock = clock; // @[:@34374.4]
  assign x532_sub_1_reset = reset; // @[:@34375.4]
  assign x532_sub_1_io_a = _T_806[31:0]; // @[Math.scala 192:17:@34376.4]
  assign x532_sub_1_io_b = _T_809[31:0]; // @[Math.scala 193:17:@34377.4]
  assign x532_sub_1_io_flow = io_in_x251_TREADY; // @[Math.scala 194:20:@34378.4]
  assign RetimeWrapper_37_clock = clock; // @[:@34384.4]
  assign RetimeWrapper_37_reset = reset; // @[:@34385.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34387.4]
  assign RetimeWrapper_37_io_in = _T_414 ? 32'h0 : _T_416; // @[package.scala 94:16:@34386.4]
  assign x341_sum_1_clock = clock; // @[:@34393.4]
  assign x341_sum_1_reset = reset; // @[:@34394.4]
  assign x341_sum_1_io_a = x532_sub_1_io_result; // @[Math.scala 151:17:@34395.4]
  assign x341_sum_1_io_b = RetimeWrapper_37_io_out; // @[Math.scala 152:17:@34396.4]
  assign x341_sum_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@34397.4]
  assign RetimeWrapper_38_clock = clock; // @[:@34403.4]
  assign RetimeWrapper_38_reset = reset; // @[:@34404.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34406.4]
  assign RetimeWrapper_38_io_in = $unsigned(_T_776); // @[package.scala 94:16:@34405.4]
  assign RetimeWrapper_39_clock = clock; // @[:@34412.4]
  assign RetimeWrapper_39_reset = reset; // @[:@34413.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34415.4]
  assign RetimeWrapper_39_io_in = ~ x336; // @[package.scala 94:16:@34414.4]
  assign RetimeWrapper_40_clock = clock; // @[:@34424.4]
  assign RetimeWrapper_40_reset = reset; // @[:@34425.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34427.4]
  assign RetimeWrapper_40_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34426.4]
  assign RetimeWrapper_41_clock = clock; // @[:@34445.4]
  assign RetimeWrapper_41_reset = reset; // @[:@34446.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34448.4]
  assign RetimeWrapper_41_io_in = $signed(_T_521) < $signed(32'sh0); // @[package.scala 94:16:@34447.4]
  assign RetimeWrapper_42_clock = clock; // @[:@34460.4]
  assign RetimeWrapper_42_reset = reset; // @[:@34461.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34463.4]
  assign RetimeWrapper_42_io_in = _T_330 ? 32'h0 : _T_332; // @[package.scala 94:16:@34462.4]
  assign x346_sum_1_clock = clock; // @[:@34471.4]
  assign x346_sum_1_reset = reset; // @[:@34472.4]
  assign x346_sum_1_io_a = x532_sub_1_io_result; // @[Math.scala 151:17:@34473.4]
  assign x346_sum_1_io_b = RetimeWrapper_42_io_out; // @[Math.scala 152:17:@34474.4]
  assign x346_sum_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@34475.4]
  assign RetimeWrapper_43_clock = clock; // @[:@34481.4]
  assign RetimeWrapper_43_reset = reset; // @[:@34482.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34484.4]
  assign RetimeWrapper_43_io_in = ~ x344; // @[package.scala 94:16:@34483.4]
  assign RetimeWrapper_44_clock = clock; // @[:@34493.4]
  assign RetimeWrapper_44_reset = reset; // @[:@34494.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34496.4]
  assign RetimeWrapper_44_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34495.4]
  assign RetimeWrapper_45_clock = clock; // @[:@34520.4]
  assign RetimeWrapper_45_reset = reset; // @[:@34521.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34523.4]
  assign RetimeWrapper_45_io_in = _T_608 ? 32'h0 : _T_610; // @[package.scala 94:16:@34522.4]
  assign x351_sum_1_clock = clock; // @[:@34529.4]
  assign x351_sum_1_reset = reset; // @[:@34530.4]
  assign x351_sum_1_io_a = x532_sub_1_io_result; // @[Math.scala 151:17:@34531.4]
  assign x351_sum_1_io_b = RetimeWrapper_45_io_out; // @[Math.scala 152:17:@34532.4]
  assign x351_sum_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@34533.4]
  assign RetimeWrapper_46_clock = clock; // @[:@34539.4]
  assign RetimeWrapper_46_reset = reset; // @[:@34540.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34542.4]
  assign RetimeWrapper_46_io_in = ~ x349; // @[package.scala 94:16:@34541.4]
  assign RetimeWrapper_47_clock = clock; // @[:@34551.4]
  assign RetimeWrapper_47_reset = reset; // @[:@34552.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34554.4]
  assign RetimeWrapper_47_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34553.4]
  assign RetimeWrapper_48_clock = clock; // @[:@34578.4]
  assign RetimeWrapper_48_reset = reset; // @[:@34579.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34581.4]
  assign RetimeWrapper_48_io_in = _T_699 ? 32'h0 : _T_701; // @[package.scala 94:16:@34580.4]
  assign x356_sum_1_clock = clock; // @[:@34587.4]
  assign x356_sum_1_reset = reset; // @[:@34588.4]
  assign x356_sum_1_io_a = x532_sub_1_io_result; // @[Math.scala 151:17:@34589.4]
  assign x356_sum_1_io_b = RetimeWrapper_48_io_out; // @[Math.scala 152:17:@34590.4]
  assign x356_sum_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@34591.4]
  assign RetimeWrapper_49_clock = clock; // @[:@34597.4]
  assign RetimeWrapper_49_reset = reset; // @[:@34598.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34600.4]
  assign RetimeWrapper_49_io_in = ~ x354; // @[package.scala 94:16:@34599.4]
  assign RetimeWrapper_50_clock = clock; // @[:@34609.4]
  assign RetimeWrapper_50_reset = reset; // @[:@34610.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34612.4]
  assign RetimeWrapper_50_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34611.4]
  assign x359_rdrow_1_clock = clock; // @[:@34632.4]
  assign x359_rdrow_1_reset = reset; // @[:@34633.4]
  assign x359_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@34634.4]
  assign x359_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@34635.4]
  assign x359_rdrow_1_io_flow = io_in_x251_TREADY; // @[Math.scala 194:20:@34636.4]
  assign x537_sub_1_clock = clock; // @[:@34704.4]
  assign x537_sub_1_reset = reset; // @[:@34705.4]
  assign x537_sub_1_io_a = _T_1016[31:0]; // @[Math.scala 192:17:@34706.4]
  assign x537_sub_1_io_b = _T_1019[31:0]; // @[Math.scala 193:17:@34707.4]
  assign x537_sub_1_io_flow = io_in_x251_TREADY; // @[Math.scala 194:20:@34708.4]
  assign x367_sum_1_clock = clock; // @[:@34714.4]
  assign x367_sum_1_reset = reset; // @[:@34715.4]
  assign x367_sum_1_io_a = x537_sub_1_io_result; // @[Math.scala 151:17:@34716.4]
  assign x367_sum_1_io_b = RetimeWrapper_37_io_out; // @[Math.scala 152:17:@34717.4]
  assign x367_sum_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@34718.4]
  assign RetimeWrapper_51_clock = clock; // @[:@34724.4]
  assign RetimeWrapper_51_reset = reset; // @[:@34725.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34727.4]
  assign RetimeWrapper_51_io_in = $unsigned(_T_986); // @[package.scala 94:16:@34726.4]
  assign RetimeWrapper_52_clock = clock; // @[:@34733.4]
  assign RetimeWrapper_52_reset = reset; // @[:@34734.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34736.4]
  assign RetimeWrapper_52_io_in = ~ x362; // @[package.scala 94:16:@34735.4]
  assign RetimeWrapper_53_clock = clock; // @[:@34745.4]
  assign RetimeWrapper_53_reset = reset; // @[:@34746.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34748.4]
  assign RetimeWrapper_53_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34747.4]
  assign x372_sum_1_clock = clock; // @[:@34772.4]
  assign x372_sum_1_reset = reset; // @[:@34773.4]
  assign x372_sum_1_io_a = x537_sub_1_io_result; // @[Math.scala 151:17:@34774.4]
  assign x372_sum_1_io_b = RetimeWrapper_42_io_out; // @[Math.scala 152:17:@34775.4]
  assign x372_sum_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@34776.4]
  assign RetimeWrapper_54_clock = clock; // @[:@34782.4]
  assign RetimeWrapper_54_reset = reset; // @[:@34783.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34785.4]
  assign RetimeWrapper_54_io_in = ~ x370; // @[package.scala 94:16:@34784.4]
  assign RetimeWrapper_55_clock = clock; // @[:@34794.4]
  assign RetimeWrapper_55_reset = reset; // @[:@34795.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34797.4]
  assign RetimeWrapper_55_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34796.4]
  assign x377_sum_1_clock = clock; // @[:@34821.4]
  assign x377_sum_1_reset = reset; // @[:@34822.4]
  assign x377_sum_1_io_a = x537_sub_1_io_result; // @[Math.scala 151:17:@34823.4]
  assign x377_sum_1_io_b = RetimeWrapper_45_io_out; // @[Math.scala 152:17:@34824.4]
  assign x377_sum_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@34825.4]
  assign RetimeWrapper_56_clock = clock; // @[:@34831.4]
  assign RetimeWrapper_56_reset = reset; // @[:@34832.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34834.4]
  assign RetimeWrapper_56_io_in = ~ x375; // @[package.scala 94:16:@34833.4]
  assign RetimeWrapper_57_clock = clock; // @[:@34843.4]
  assign RetimeWrapper_57_reset = reset; // @[:@34844.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34846.4]
  assign RetimeWrapper_57_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34845.4]
  assign x382_sum_1_clock = clock; // @[:@34872.4]
  assign x382_sum_1_reset = reset; // @[:@34873.4]
  assign x382_sum_1_io_a = x537_sub_1_io_result; // @[Math.scala 151:17:@34874.4]
  assign x382_sum_1_io_b = RetimeWrapper_48_io_out; // @[Math.scala 152:17:@34875.4]
  assign x382_sum_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@34876.4]
  assign RetimeWrapper_58_clock = clock; // @[:@34882.4]
  assign RetimeWrapper_58_reset = reset; // @[:@34883.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34885.4]
  assign RetimeWrapper_58_io_in = ~ x380; // @[package.scala 94:16:@34884.4]
  assign RetimeWrapper_59_clock = clock; // @[:@34894.4]
  assign RetimeWrapper_59_reset = reset; // @[:@34895.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@34897.4]
  assign RetimeWrapper_59_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@34896.4]
  assign x385_1_clock = clock; // @[:@34917.4]
  assign x385_1_io_a = x285_lb_0_io_rPort_2_output_0; // @[Math.scala 263:17:@34919.4]
  assign x385_1_io_b = 32'h1; // @[Math.scala 264:17:@34920.4]
  assign x385_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@34921.4]
  assign x386_1_clock = clock; // @[:@34929.4]
  assign x386_1_io_a = x285_lb_0_io_rPort_4_output_0; // @[Math.scala 263:17:@34931.4]
  assign x386_1_io_b = 32'h2; // @[Math.scala 264:17:@34932.4]
  assign x386_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@34933.4]
  assign x387_1_clock = clock; // @[:@34941.4]
  assign x387_1_io_a = x285_lb_0_io_rPort_11_output_0; // @[Math.scala 263:17:@34943.4]
  assign x387_1_io_b = 32'h1; // @[Math.scala 264:17:@34944.4]
  assign x387_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@34945.4]
  assign x388_1_clock = clock; // @[:@34953.4]
  assign x388_1_io_a = x285_lb_0_io_rPort_5_output_0; // @[Math.scala 263:17:@34955.4]
  assign x388_1_io_b = 32'h2; // @[Math.scala 264:17:@34956.4]
  assign x388_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@34957.4]
  assign x389_1_clock = clock; // @[:@34965.4]
  assign x389_1_io_a = x285_lb_0_io_rPort_0_output_0; // @[Math.scala 263:17:@34967.4]
  assign x389_1_io_b = 32'h4; // @[Math.scala 264:17:@34968.4]
  assign x389_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@34969.4]
  assign x390_1_clock = clock; // @[:@34977.4]
  assign x390_1_io_a = x285_lb_0_io_rPort_1_output_0; // @[Math.scala 263:17:@34979.4]
  assign x390_1_io_b = 32'h2; // @[Math.scala 264:17:@34980.4]
  assign x390_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@34981.4]
  assign x391_1_clock = clock; // @[:@34989.4]
  assign x391_1_io_a = x285_lb_0_io_rPort_7_output_0; // @[Math.scala 263:17:@34991.4]
  assign x391_1_io_b = 32'h1; // @[Math.scala 264:17:@34992.4]
  assign x391_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@34993.4]
  assign x392_1_clock = clock; // @[:@35001.4]
  assign x392_1_io_a = x285_lb_0_io_rPort_10_output_0; // @[Math.scala 263:17:@35003.4]
  assign x392_1_io_b = 32'h2; // @[Math.scala 264:17:@35004.4]
  assign x392_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35005.4]
  assign x393_1_clock = clock; // @[:@35013.4]
  assign x393_1_io_a = x285_lb_0_io_rPort_8_output_0; // @[Math.scala 263:17:@35015.4]
  assign x393_1_io_b = 32'h1; // @[Math.scala 264:17:@35016.4]
  assign x393_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35017.4]
  assign x394_x7_1_clock = clock; // @[:@35023.4]
  assign x394_x7_1_reset = reset; // @[:@35024.4]
  assign x394_x7_1_io_a = x385_1_io_result; // @[Math.scala 151:17:@35025.4]
  assign x394_x7_1_io_b = x386_1_io_result; // @[Math.scala 152:17:@35026.4]
  assign x394_x7_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35027.4]
  assign x395_x8_1_clock = clock; // @[:@35033.4]
  assign x395_x8_1_reset = reset; // @[:@35034.4]
  assign x395_x8_1_io_a = x387_1_io_result; // @[Math.scala 151:17:@35035.4]
  assign x395_x8_1_io_b = x388_1_io_result; // @[Math.scala 152:17:@35036.4]
  assign x395_x8_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35037.4]
  assign x396_x7_1_clock = clock; // @[:@35043.4]
  assign x396_x7_1_reset = reset; // @[:@35044.4]
  assign x396_x7_1_io_a = x389_1_io_result; // @[Math.scala 151:17:@35045.4]
  assign x396_x7_1_io_b = x390_1_io_result; // @[Math.scala 152:17:@35046.4]
  assign x396_x7_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35047.4]
  assign x397_x8_1_clock = clock; // @[:@35053.4]
  assign x397_x8_1_reset = reset; // @[:@35054.4]
  assign x397_x8_1_io_a = x391_1_io_result; // @[Math.scala 151:17:@35055.4]
  assign x397_x8_1_io_b = x392_1_io_result; // @[Math.scala 152:17:@35056.4]
  assign x397_x8_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35057.4]
  assign x398_x7_1_clock = clock; // @[:@35063.4]
  assign x398_x7_1_reset = reset; // @[:@35064.4]
  assign x398_x7_1_io_a = x394_x7_1_io_result; // @[Math.scala 151:17:@35065.4]
  assign x398_x7_1_io_b = x395_x8_1_io_result; // @[Math.scala 152:17:@35066.4]
  assign x398_x7_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35067.4]
  assign x399_x8_1_clock = clock; // @[:@35073.4]
  assign x399_x8_1_reset = reset; // @[:@35074.4]
  assign x399_x8_1_io_a = x396_x7_1_io_result; // @[Math.scala 151:17:@35075.4]
  assign x399_x8_1_io_b = x397_x8_1_io_result; // @[Math.scala 152:17:@35076.4]
  assign x399_x8_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35077.4]
  assign x400_x7_1_clock = clock; // @[:@35083.4]
  assign x400_x7_1_reset = reset; // @[:@35084.4]
  assign x400_x7_1_io_a = x398_x7_1_io_result; // @[Math.scala 151:17:@35085.4]
  assign x400_x7_1_io_b = x399_x8_1_io_result; // @[Math.scala 152:17:@35086.4]
  assign x400_x7_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35087.4]
  assign RetimeWrapper_60_clock = clock; // @[:@35093.4]
  assign RetimeWrapper_60_reset = reset; // @[:@35094.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35096.4]
  assign RetimeWrapper_60_io_in = x393_1_io_result; // @[package.scala 94:16:@35095.4]
  assign x401_sum_1_clock = clock; // @[:@35102.4]
  assign x401_sum_1_reset = reset; // @[:@35103.4]
  assign x401_sum_1_io_a = x400_x7_1_io_result; // @[Math.scala 151:17:@35104.4]
  assign x401_sum_1_io_b = RetimeWrapper_60_io_out; // @[Math.scala 152:17:@35105.4]
  assign x401_sum_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35106.4]
  assign x402_1_io_b = x401_sum_1_io_result; // @[Math.scala 721:17:@35114.4]
  assign x403_mul_1_clock = clock; // @[:@35123.4]
  assign x403_mul_1_io_a = x402_1_io_result; // @[Math.scala 263:17:@35125.4]
  assign x403_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@35126.4]
  assign x403_mul_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35127.4]
  assign x404_1_io_b = x403_mul_1_io_result; // @[Math.scala 721:17:@35135.4]
  assign x405_1_clock = clock; // @[:@35144.4]
  assign x405_1_io_a = x285_lb_0_io_rPort_4_output_0; // @[Math.scala 263:17:@35146.4]
  assign x405_1_io_b = 32'h1; // @[Math.scala 264:17:@35147.4]
  assign x405_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35148.4]
  assign x406_1_clock = clock; // @[:@35156.4]
  assign x406_1_io_a = x285_lb_0_io_rPort_11_output_0; // @[Math.scala 263:17:@35158.4]
  assign x406_1_io_b = 32'h2; // @[Math.scala 264:17:@35159.4]
  assign x406_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35160.4]
  assign x407_1_clock = clock; // @[:@35168.4]
  assign x407_1_io_a = x285_lb_0_io_rPort_6_output_0; // @[Math.scala 263:17:@35170.4]
  assign x407_1_io_b = 32'h1; // @[Math.scala 264:17:@35171.4]
  assign x407_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35172.4]
  assign x408_1_clock = clock; // @[:@35180.4]
  assign x408_1_io_a = x285_lb_0_io_rPort_0_output_0; // @[Math.scala 263:17:@35182.4]
  assign x408_1_io_b = 32'h2; // @[Math.scala 264:17:@35183.4]
  assign x408_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35184.4]
  assign x409_1_clock = clock; // @[:@35192.4]
  assign x409_1_io_a = x285_lb_0_io_rPort_1_output_0; // @[Math.scala 263:17:@35194.4]
  assign x409_1_io_b = 32'h4; // @[Math.scala 264:17:@35195.4]
  assign x409_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35196.4]
  assign x410_1_clock = clock; // @[:@35204.4]
  assign x410_1_io_a = x285_lb_0_io_rPort_3_output_0; // @[Math.scala 263:17:@35206.4]
  assign x410_1_io_b = 32'h2; // @[Math.scala 264:17:@35207.4]
  assign x410_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35208.4]
  assign x411_1_clock = clock; // @[:@35216.4]
  assign x411_1_io_a = x285_lb_0_io_rPort_10_output_0; // @[Math.scala 263:17:@35218.4]
  assign x411_1_io_b = 32'h1; // @[Math.scala 264:17:@35219.4]
  assign x411_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35220.4]
  assign x412_1_clock = clock; // @[:@35228.4]
  assign x412_1_io_a = x285_lb_0_io_rPort_8_output_0; // @[Math.scala 263:17:@35230.4]
  assign x412_1_io_b = 32'h2; // @[Math.scala 264:17:@35231.4]
  assign x412_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35232.4]
  assign x413_1_clock = clock; // @[:@35240.4]
  assign x413_1_io_a = x285_lb_0_io_rPort_9_output_0; // @[Math.scala 263:17:@35242.4]
  assign x413_1_io_b = 32'h1; // @[Math.scala 264:17:@35243.4]
  assign x413_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35244.4]
  assign x414_x7_1_clock = clock; // @[:@35250.4]
  assign x414_x7_1_reset = reset; // @[:@35251.4]
  assign x414_x7_1_io_a = x405_1_io_result; // @[Math.scala 151:17:@35252.4]
  assign x414_x7_1_io_b = x406_1_io_result; // @[Math.scala 152:17:@35253.4]
  assign x414_x7_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35254.4]
  assign x415_x8_1_clock = clock; // @[:@35260.4]
  assign x415_x8_1_reset = reset; // @[:@35261.4]
  assign x415_x8_1_io_a = x407_1_io_result; // @[Math.scala 151:17:@35262.4]
  assign x415_x8_1_io_b = x408_1_io_result; // @[Math.scala 152:17:@35263.4]
  assign x415_x8_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35264.4]
  assign x416_x7_1_clock = clock; // @[:@35270.4]
  assign x416_x7_1_reset = reset; // @[:@35271.4]
  assign x416_x7_1_io_a = x409_1_io_result; // @[Math.scala 151:17:@35272.4]
  assign x416_x7_1_io_b = x410_1_io_result; // @[Math.scala 152:17:@35273.4]
  assign x416_x7_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35274.4]
  assign x417_x8_1_clock = clock; // @[:@35280.4]
  assign x417_x8_1_reset = reset; // @[:@35281.4]
  assign x417_x8_1_io_a = x411_1_io_result; // @[Math.scala 151:17:@35282.4]
  assign x417_x8_1_io_b = x412_1_io_result; // @[Math.scala 152:17:@35283.4]
  assign x417_x8_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35284.4]
  assign x418_x7_1_clock = clock; // @[:@35290.4]
  assign x418_x7_1_reset = reset; // @[:@35291.4]
  assign x418_x7_1_io_a = x414_x7_1_io_result; // @[Math.scala 151:17:@35292.4]
  assign x418_x7_1_io_b = x415_x8_1_io_result; // @[Math.scala 152:17:@35293.4]
  assign x418_x7_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35294.4]
  assign x419_x8_1_clock = clock; // @[:@35300.4]
  assign x419_x8_1_reset = reset; // @[:@35301.4]
  assign x419_x8_1_io_a = x416_x7_1_io_result; // @[Math.scala 151:17:@35302.4]
  assign x419_x8_1_io_b = x417_x8_1_io_result; // @[Math.scala 152:17:@35303.4]
  assign x419_x8_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35304.4]
  assign x420_x7_1_clock = clock; // @[:@35310.4]
  assign x420_x7_1_reset = reset; // @[:@35311.4]
  assign x420_x7_1_io_a = x418_x7_1_io_result; // @[Math.scala 151:17:@35312.4]
  assign x420_x7_1_io_b = x419_x8_1_io_result; // @[Math.scala 152:17:@35313.4]
  assign x420_x7_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35314.4]
  assign RetimeWrapper_61_clock = clock; // @[:@35320.4]
  assign RetimeWrapper_61_reset = reset; // @[:@35321.4]
  assign RetimeWrapper_61_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35323.4]
  assign RetimeWrapper_61_io_in = x413_1_io_result; // @[package.scala 94:16:@35322.4]
  assign x421_sum_1_clock = clock; // @[:@35329.4]
  assign x421_sum_1_reset = reset; // @[:@35330.4]
  assign x421_sum_1_io_a = x420_x7_1_io_result; // @[Math.scala 151:17:@35331.4]
  assign x421_sum_1_io_b = RetimeWrapper_61_io_out; // @[Math.scala 152:17:@35332.4]
  assign x421_sum_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35333.4]
  assign x422_1_io_b = x421_sum_1_io_result; // @[Math.scala 721:17:@35341.4]
  assign x423_mul_1_clock = clock; // @[:@35350.4]
  assign x423_mul_1_io_a = x422_1_io_result; // @[Math.scala 263:17:@35352.4]
  assign x423_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@35353.4]
  assign x423_mul_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35354.4]
  assign x424_1_io_b = x423_mul_1_io_result; // @[Math.scala 721:17:@35362.4]
  assign RetimeWrapper_62_clock = clock; // @[:@35369.4]
  assign RetimeWrapper_62_reset = reset; // @[:@35370.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35372.4]
  assign RetimeWrapper_62_io_in = x424_1_io_result; // @[package.scala 94:16:@35371.4]
  assign RetimeWrapper_63_clock = clock; // @[:@35378.4]
  assign RetimeWrapper_63_reset = reset; // @[:@35379.4]
  assign RetimeWrapper_63_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35381.4]
  assign RetimeWrapper_63_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@35380.4]
  assign RetimeWrapper_64_clock = clock; // @[:@35387.4]
  assign RetimeWrapper_64_reset = reset; // @[:@35388.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35390.4]
  assign RetimeWrapper_64_io_in = $unsigned(_T_260); // @[package.scala 94:16:@35389.4]
  assign RetimeWrapper_65_clock = clock; // @[:@35396.4]
  assign RetimeWrapper_65_reset = reset; // @[:@35397.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35399.4]
  assign RetimeWrapper_65_io_in = $unsigned(_T_272); // @[package.scala 94:16:@35398.4]
  assign RetimeWrapper_66_clock = clock; // @[:@35405.4]
  assign RetimeWrapper_66_reset = reset; // @[:@35406.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35408.4]
  assign RetimeWrapper_66_io_in = x295_sum_1_io_result; // @[package.scala 94:16:@35407.4]
  assign RetimeWrapper_67_clock = clock; // @[:@35414.4]
  assign RetimeWrapper_67_reset = reset; // @[:@35415.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35417.4]
  assign RetimeWrapper_67_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@35416.4]
  assign RetimeWrapper_68_clock = clock; // @[:@35425.4]
  assign RetimeWrapper_68_reset = reset; // @[:@35426.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35428.4]
  assign RetimeWrapper_68_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35427.4]
  assign RetimeWrapper_69_clock = clock; // @[:@35446.4]
  assign RetimeWrapper_69_reset = reset; // @[:@35447.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35449.4]
  assign RetimeWrapper_69_io_in = x404_1_io_result; // @[package.scala 94:16:@35448.4]
  assign RetimeWrapper_70_clock = clock; // @[:@35455.4]
  assign RetimeWrapper_70_reset = reset; // @[:@35456.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35458.4]
  assign RetimeWrapper_70_io_in = x301_sum_1_io_result; // @[package.scala 94:16:@35457.4]
  assign RetimeWrapper_71_clock = clock; // @[:@35464.4]
  assign RetimeWrapper_71_reset = reset; // @[:@35465.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35467.4]
  assign RetimeWrapper_71_io_in = $unsigned(_T_391); // @[package.scala 94:16:@35466.4]
  assign RetimeWrapper_72_clock = clock; // @[:@35475.4]
  assign RetimeWrapper_72_reset = reset; // @[:@35476.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35478.4]
  assign RetimeWrapper_72_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35477.4]
  assign RetimeWrapper_73_clock = clock; // @[:@35496.4]
  assign RetimeWrapper_73_reset = reset; // @[:@35497.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35499.4]
  assign RetimeWrapper_73_io_in = x301_sum_1_io_result; // @[package.scala 94:16:@35498.4]
  assign RetimeWrapper_74_clock = clock; // @[:@35505.4]
  assign RetimeWrapper_74_reset = reset; // @[:@35506.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35508.4]
  assign RetimeWrapper_74_io_in = ~ x306; // @[package.scala 94:16:@35507.4]
  assign RetimeWrapper_75_clock = clock; // @[:@35514.4]
  assign RetimeWrapper_75_reset = reset; // @[:@35515.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35517.4]
  assign RetimeWrapper_75_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@35516.4]
  assign RetimeWrapper_76_clock = clock; // @[:@35523.4]
  assign RetimeWrapper_76_reset = reset; // @[:@35524.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35526.4]
  assign RetimeWrapper_76_io_in = $unsigned(_T_260); // @[package.scala 94:16:@35525.4]
  assign RetimeWrapper_77_clock = clock; // @[:@35532.4]
  assign RetimeWrapper_77_reset = reset; // @[:@35533.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35535.4]
  assign RetimeWrapper_77_io_in = $unsigned(_T_391); // @[package.scala 94:16:@35534.4]
  assign RetimeWrapper_78_clock = clock; // @[:@35541.4]
  assign RetimeWrapper_78_reset = reset; // @[:@35542.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35544.4]
  assign RetimeWrapper_78_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@35543.4]
  assign RetimeWrapper_79_clock = clock; // @[:@35553.4]
  assign RetimeWrapper_79_reset = reset; // @[:@35554.4]
  assign RetimeWrapper_79_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35556.4]
  assign RetimeWrapper_79_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35555.4]
  assign RetimeWrapper_80_clock = clock; // @[:@35574.4]
  assign RetimeWrapper_80_reset = reset; // @[:@35575.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35577.4]
  assign RetimeWrapper_80_io_in = ~ x311; // @[package.scala 94:16:@35576.4]
  assign RetimeWrapper_81_clock = clock; // @[:@35583.4]
  assign RetimeWrapper_81_reset = reset; // @[:@35584.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35586.4]
  assign RetimeWrapper_81_io_in = $unsigned(_T_272); // @[package.scala 94:16:@35585.4]
  assign RetimeWrapper_82_clock = clock; // @[:@35592.4]
  assign RetimeWrapper_82_reset = reset; // @[:@35593.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35595.4]
  assign RetimeWrapper_82_io_in = x295_sum_1_io_result; // @[package.scala 94:16:@35594.4]
  assign RetimeWrapper_83_clock = clock; // @[:@35604.4]
  assign RetimeWrapper_83_reset = reset; // @[:@35605.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35607.4]
  assign RetimeWrapper_83_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35606.4]
  assign RetimeWrapper_84_clock = clock; // @[:@35625.4]
  assign RetimeWrapper_84_reset = reset; // @[:@35626.4]
  assign RetimeWrapper_84_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35628.4]
  assign RetimeWrapper_84_io_in = x321_sum_1_io_result; // @[package.scala 94:16:@35627.4]
  assign RetimeWrapper_85_clock = clock; // @[:@35634.4]
  assign RetimeWrapper_85_reset = reset; // @[:@35635.4]
  assign RetimeWrapper_85_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35637.4]
  assign RetimeWrapper_85_io_in = $unsigned(_T_585); // @[package.scala 94:16:@35636.4]
  assign RetimeWrapper_86_clock = clock; // @[:@35643.4]
  assign RetimeWrapper_86_reset = reset; // @[:@35644.4]
  assign RetimeWrapper_86_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35646.4]
  assign RetimeWrapper_86_io_in = ~ x317; // @[package.scala 94:16:@35645.4]
  assign RetimeWrapper_87_clock = clock; // @[:@35655.4]
  assign RetimeWrapper_87_reset = reset; // @[:@35656.4]
  assign RetimeWrapper_87_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35658.4]
  assign RetimeWrapper_87_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35657.4]
  assign RetimeWrapper_88_clock = clock; // @[:@35676.4]
  assign RetimeWrapper_88_reset = reset; // @[:@35677.4]
  assign RetimeWrapper_88_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35679.4]
  assign RetimeWrapper_88_io_in = $unsigned(_T_776); // @[package.scala 94:16:@35678.4]
  assign RetimeWrapper_89_clock = clock; // @[:@35685.4]
  assign RetimeWrapper_89_reset = reset; // @[:@35686.4]
  assign RetimeWrapper_89_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35688.4]
  assign RetimeWrapper_89_io_in = x341_sum_1_io_result; // @[package.scala 94:16:@35687.4]
  assign RetimeWrapper_90_clock = clock; // @[:@35694.4]
  assign RetimeWrapper_90_reset = reset; // @[:@35695.4]
  assign RetimeWrapper_90_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35697.4]
  assign RetimeWrapper_90_io_in = ~ x336; // @[package.scala 94:16:@35696.4]
  assign RetimeWrapper_91_clock = clock; // @[:@35706.4]
  assign RetimeWrapper_91_reset = reset; // @[:@35707.4]
  assign RetimeWrapper_91_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35709.4]
  assign RetimeWrapper_91_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35708.4]
  assign RetimeWrapper_92_clock = clock; // @[:@35727.4]
  assign RetimeWrapper_92_reset = reset; // @[:@35728.4]
  assign RetimeWrapper_92_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35730.4]
  assign RetimeWrapper_92_io_in = ~ x344; // @[package.scala 94:16:@35729.4]
  assign RetimeWrapper_93_clock = clock; // @[:@35736.4]
  assign RetimeWrapper_93_reset = reset; // @[:@35737.4]
  assign RetimeWrapper_93_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35739.4]
  assign RetimeWrapper_93_io_in = x346_sum_1_io_result; // @[package.scala 94:16:@35738.4]
  assign RetimeWrapper_94_clock = clock; // @[:@35748.4]
  assign RetimeWrapper_94_reset = reset; // @[:@35749.4]
  assign RetimeWrapper_94_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35751.4]
  assign RetimeWrapper_94_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35750.4]
  assign RetimeWrapper_95_clock = clock; // @[:@35769.4]
  assign RetimeWrapper_95_reset = reset; // @[:@35770.4]
  assign RetimeWrapper_95_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35772.4]
  assign RetimeWrapper_95_io_in = ~ x349; // @[package.scala 94:16:@35771.4]
  assign RetimeWrapper_96_clock = clock; // @[:@35778.4]
  assign RetimeWrapper_96_reset = reset; // @[:@35779.4]
  assign RetimeWrapper_96_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35781.4]
  assign RetimeWrapper_96_io_in = x351_sum_1_io_result; // @[package.scala 94:16:@35780.4]
  assign RetimeWrapper_97_clock = clock; // @[:@35790.4]
  assign RetimeWrapper_97_reset = reset; // @[:@35791.4]
  assign RetimeWrapper_97_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@35793.4]
  assign RetimeWrapper_97_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@35792.4]
  assign x441_1_clock = clock; // @[:@35815.4]
  assign x441_1_io_a = x286_lb2_0_io_rPort_1_output_0; // @[Math.scala 263:17:@35817.4]
  assign x441_1_io_b = 32'h1; // @[Math.scala 264:17:@35818.4]
  assign x441_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35819.4]
  assign x442_1_clock = clock; // @[:@35827.4]
  assign x442_1_io_a = x286_lb2_0_io_rPort_3_output_0; // @[Math.scala 263:17:@35829.4]
  assign x442_1_io_b = 32'h2; // @[Math.scala 264:17:@35830.4]
  assign x442_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35831.4]
  assign x443_1_clock = clock; // @[:@35839.4]
  assign x443_1_io_a = x286_lb2_0_io_rPort_2_output_0; // @[Math.scala 263:17:@35841.4]
  assign x443_1_io_b = 32'h4; // @[Math.scala 264:17:@35842.4]
  assign x443_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35843.4]
  assign x444_1_clock = clock; // @[:@35851.4]
  assign x444_1_io_a = x286_lb2_0_io_rPort_5_output_0; // @[Math.scala 263:17:@35853.4]
  assign x444_1_io_b = 32'h1; // @[Math.scala 264:17:@35854.4]
  assign x444_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35855.4]
  assign x445_x9_1_clock = clock; // @[:@35861.4]
  assign x445_x9_1_reset = reset; // @[:@35862.4]
  assign x445_x9_1_io_a = x441_1_io_result; // @[Math.scala 151:17:@35863.4]
  assign x445_x9_1_io_b = x442_1_io_result; // @[Math.scala 152:17:@35864.4]
  assign x445_x9_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35865.4]
  assign x446_x10_1_clock = clock; // @[:@35873.4]
  assign x446_x10_1_reset = reset; // @[:@35874.4]
  assign x446_x10_1_io_a = x443_1_io_result; // @[Math.scala 151:17:@35875.4]
  assign x446_x10_1_io_b = x444_1_io_result; // @[Math.scala 152:17:@35876.4]
  assign x446_x10_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35877.4]
  assign x447_sum_1_clock = clock; // @[:@35883.4]
  assign x447_sum_1_reset = reset; // @[:@35884.4]
  assign x447_sum_1_io_a = x445_x9_1_io_result; // @[Math.scala 151:17:@35885.4]
  assign x447_sum_1_io_b = x446_x10_1_io_result; // @[Math.scala 152:17:@35886.4]
  assign x447_sum_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35887.4]
  assign x448_1_io_b = x447_sum_1_io_result; // @[Math.scala 721:17:@35895.4]
  assign x449_mul_1_clock = clock; // @[:@35904.4]
  assign x449_mul_1_io_a = x448_1_io_result; // @[Math.scala 263:17:@35906.4]
  assign x449_mul_1_io_b = 32'h10; // @[Math.scala 264:17:@35907.4]
  assign x449_mul_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35908.4]
  assign x450_1_io_b = x449_mul_1_io_result; // @[Math.scala 721:17:@35916.4]
  assign x451_1_clock = clock; // @[:@35925.4]
  assign x451_1_io_a = x286_lb2_0_io_rPort_3_output_0; // @[Math.scala 263:17:@35927.4]
  assign x451_1_io_b = 32'h1; // @[Math.scala 264:17:@35928.4]
  assign x451_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35929.4]
  assign x452_1_clock = clock; // @[:@35937.4]
  assign x452_1_io_a = x286_lb2_0_io_rPort_4_output_0; // @[Math.scala 263:17:@35939.4]
  assign x452_1_io_b = 32'h2; // @[Math.scala 264:17:@35940.4]
  assign x452_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35941.4]
  assign x453_1_clock = clock; // @[:@35949.4]
  assign x453_1_io_a = x286_lb2_0_io_rPort_5_output_0; // @[Math.scala 263:17:@35951.4]
  assign x453_1_io_b = 32'h4; // @[Math.scala 264:17:@35952.4]
  assign x453_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35953.4]
  assign x454_1_clock = clock; // @[:@35961.4]
  assign x454_1_io_a = x286_lb2_0_io_rPort_0_output_0; // @[Math.scala 263:17:@35963.4]
  assign x454_1_io_b = 32'h1; // @[Math.scala 264:17:@35964.4]
  assign x454_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@35965.4]
  assign x455_x9_1_clock = clock; // @[:@35971.4]
  assign x455_x9_1_reset = reset; // @[:@35972.4]
  assign x455_x9_1_io_a = x451_1_io_result; // @[Math.scala 151:17:@35973.4]
  assign x455_x9_1_io_b = x452_1_io_result; // @[Math.scala 152:17:@35974.4]
  assign x455_x9_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35975.4]
  assign x456_x10_1_clock = clock; // @[:@35981.4]
  assign x456_x10_1_reset = reset; // @[:@35982.4]
  assign x456_x10_1_io_a = x453_1_io_result; // @[Math.scala 151:17:@35983.4]
  assign x456_x10_1_io_b = x454_1_io_result; // @[Math.scala 152:17:@35984.4]
  assign x456_x10_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35985.4]
  assign x457_sum_1_clock = clock; // @[:@35991.4]
  assign x457_sum_1_reset = reset; // @[:@35992.4]
  assign x457_sum_1_io_a = x455_x9_1_io_result; // @[Math.scala 151:17:@35993.4]
  assign x457_sum_1_io_b = x456_x10_1_io_result; // @[Math.scala 152:17:@35994.4]
  assign x457_sum_1_io_flow = io_in_x251_TREADY; // @[Math.scala 153:20:@35995.4]
  assign x458_1_io_b = x457_sum_1_io_result; // @[Math.scala 721:17:@36003.4]
  assign x459_mul_1_clock = clock; // @[:@36012.4]
  assign x459_mul_1_io_a = x458_1_io_result; // @[Math.scala 263:17:@36014.4]
  assign x459_mul_1_io_b = 32'h10; // @[Math.scala 264:17:@36015.4]
  assign x459_mul_1_io_flow = io_in_x251_TREADY; // @[Math.scala 265:20:@36016.4]
  assign x460_1_io_b = x459_mul_1_io_result; // @[Math.scala 721:17:@36024.4]
  assign RetimeWrapper_98_clock = clock; // @[:@36037.4]
  assign RetimeWrapper_98_reset = reset; // @[:@36038.4]
  assign RetimeWrapper_98_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@36040.4]
  assign RetimeWrapper_98_io_in = {x450_number,x460_number}; // @[package.scala 94:16:@36039.4]
  assign RetimeWrapper_99_clock = clock; // @[:@36046.4]
  assign RetimeWrapper_99_reset = reset; // @[:@36047.4]
  assign RetimeWrapper_99_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@36049.4]
  assign RetimeWrapper_99_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@36048.4]
  assign RetimeWrapper_100_clock = clock; // @[:@36055.4]
  assign RetimeWrapper_100_reset = reset; // @[:@36056.4]
  assign RetimeWrapper_100_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@36058.4]
  assign RetimeWrapper_100_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@36057.4]
  assign RetimeWrapper_101_clock = clock; // @[:@36064.4]
  assign RetimeWrapper_101_reset = reset; // @[:@36065.4]
  assign RetimeWrapper_101_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@36067.4]
  assign RetimeWrapper_101_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@36066.4]
endmodule
module x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1( // @[:@36085.2]
  input          clock, // @[:@36086.4]
  input          reset, // @[:@36087.4]
  output         io_in_x251_TVALID, // @[:@36088.4]
  input          io_in_x251_TREADY, // @[:@36088.4]
  output [255:0] io_in_x251_TDATA, // @[:@36088.4]
  input          io_in_x250_TVALID, // @[:@36088.4]
  output         io_in_x250_TREADY, // @[:@36088.4]
  input  [255:0] io_in_x250_TDATA, // @[:@36088.4]
  input  [7:0]   io_in_x250_TID, // @[:@36088.4]
  input  [7:0]   io_in_x250_TDEST, // @[:@36088.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@36088.4]
  input          io_sigsIn_smChildAcks_0, // @[:@36088.4]
  output         io_sigsOut_smDoneIn_0, // @[:@36088.4]
  input          io_rr // @[:@36088.4]
);
  wire  x278_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@36122.4]
  wire  x278_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@36122.4]
  wire  x278_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@36122.4]
  wire  x278_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@36122.4]
  wire [12:0] x278_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@36122.4]
  wire [12:0] x278_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@36122.4]
  wire  x278_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@36122.4]
  wire  x278_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@36122.4]
  wire  x278_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@36122.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 32:18:@36182.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 32:18:@36182.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 32:18:@36182.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 32:18:@36182.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 32:18:@36182.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 32:18:@36182.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 32:18:@36182.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 32:18:@36182.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 32:18:@36182.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 32:18:@36182.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 32:18:@36182.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 32:18:@36182.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@36210.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@36210.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@36210.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@36210.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@36210.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@36252.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@36252.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@36252.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@36252.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@36252.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@36260.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@36260.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@36260.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@36260.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@36260.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 713:24:@36294.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 713:24:@36294.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x251_TVALID; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 713:24:@36294.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x251_TREADY; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 713:24:@36294.4]
  wire [255:0] x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x251_TDATA; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 713:24:@36294.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x250_TREADY; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 713:24:@36294.4]
  wire [255:0] x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x250_TDATA; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 713:24:@36294.4]
  wire [7:0] x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x250_TID; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 713:24:@36294.4]
  wire [7:0] x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x250_TDEST; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 713:24:@36294.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 713:24:@36294.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 713:24:@36294.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 713:24:@36294.4]
  wire [31:0] x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 713:24:@36294.4]
  wire [31:0] x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 713:24:@36294.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 713:24:@36294.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 713:24:@36294.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 713:24:@36294.4]
  wire  _T_240; // @[package.scala 96:25:@36215.4 package.scala 96:25:@36216.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x466_outr_UnitPipe.scala 69:66:@36221.4]
  wire  _T_253; // @[package.scala 96:25:@36257.4 package.scala 96:25:@36258.4]
  wire  _T_259; // @[package.scala 96:25:@36265.4 package.scala 96:25:@36266.4]
  wire  _T_262; // @[SpatialBlocks.scala 138:93:@36268.4]
  wire  x465_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@36269.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:36:@36277.4]
  wire  _T_265; // @[SpatialBlocks.scala 157:78:@36278.4]
  wire  _T_272; // @[SpatialBlocks.scala 159:58:@36290.4]
  x258_ctrchain x278_ctrchain ( // @[SpatialBlocks.scala 37:22:@36122.4]
    .clock(x278_ctrchain_clock),
    .reset(x278_ctrchain_reset),
    .io_input_reset(x278_ctrchain_io_input_reset),
    .io_input_enable(x278_ctrchain_io_input_enable),
    .io_output_counts_1(x278_ctrchain_io_output_counts_1),
    .io_output_counts_0(x278_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x278_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x278_ctrchain_io_output_oobs_1),
    .io_output_done(x278_ctrchain_io_output_done)
  );
  x465_inr_Foreach_SAMPLER_BOX_sm x465_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 32:18:@36182.4]
    .clock(x465_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x465_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x465_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x465_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x465_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x465_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x465_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x465_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x465_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x465_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x465_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x465_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@36210.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@36252.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@36260.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1 x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 713:24:@36294.4]
    .clock(x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x251_TVALID(x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x251_TVALID),
    .io_in_x251_TREADY(x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x251_TREADY),
    .io_in_x251_TDATA(x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x251_TDATA),
    .io_in_x250_TREADY(x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x250_TREADY),
    .io_in_x250_TDATA(x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x250_TDATA),
    .io_in_x250_TID(x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x250_TID),
    .io_in_x250_TDEST(x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x250_TDEST),
    .io_sigsIn_backpressure(x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_240 = RetimeWrapper_io_out; // @[package.scala 96:25:@36215.4 package.scala 96:25:@36216.4]
  assign x465_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x250_TVALID | x465_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x466_outr_UnitPipe.scala 69:66:@36221.4]
  assign _T_253 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@36257.4 package.scala 96:25:@36258.4]
  assign _T_259 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@36265.4 package.scala 96:25:@36266.4]
  assign _T_262 = ~ _T_259; // @[SpatialBlocks.scala 138:93:@36268.4]
  assign x465_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_253 & _T_262; // @[SpatialBlocks.scala 138:90:@36269.4]
  assign _T_264 = x465_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@36277.4]
  assign _T_265 = ~ x465_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@36278.4]
  assign _T_272 = x465_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@36290.4]
  assign io_in_x251_TVALID = x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x251_TVALID; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 48:23:@36353.4]
  assign io_in_x251_TDATA = x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x251_TDATA; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 48:23:@36351.4]
  assign io_in_x250_TREADY = x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x250_TREADY; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 49:23:@36361.4]
  assign io_sigsOut_smDoneIn_0 = x465_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@36275.4]
  assign x278_ctrchain_clock = clock; // @[:@36123.4]
  assign x278_ctrchain_reset = reset; // @[:@36124.4]
  assign x278_ctrchain_io_input_reset = x465_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@36293.4]
  assign x278_ctrchain_io_input_enable = _T_272 & x465_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@36245.4 SpatialBlocks.scala 159:42:@36292.4]
  assign x465_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@36183.4]
  assign x465_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@36184.4]
  assign x465_inr_Foreach_SAMPLER_BOX_sm_io_enable = x465_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x465_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@36272.4]
  assign x465_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_240 : 1'h0; // @[sm_x466_outr_UnitPipe.scala 67:50:@36218.4]
  assign x465_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@36274.4]
  assign x465_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x251_TREADY | x465_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@36246.4]
  assign x465_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x466_outr_UnitPipe.scala 71:48:@36224.4]
  assign RetimeWrapper_clock = clock; // @[:@36211.4]
  assign RetimeWrapper_reset = reset; // @[:@36212.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@36214.4]
  assign RetimeWrapper_io_in = x278_ctrchain_io_output_done; // @[package.scala 94:16:@36213.4]
  assign RetimeWrapper_1_clock = clock; // @[:@36253.4]
  assign RetimeWrapper_1_reset = reset; // @[:@36254.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@36256.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@36255.4]
  assign RetimeWrapper_2_clock = clock; // @[:@36261.4]
  assign RetimeWrapper_2_reset = reset; // @[:@36262.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@36264.4]
  assign RetimeWrapper_2_io_in = x465_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@36263.4]
  assign x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@36295.4]
  assign x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@36296.4]
  assign x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x251_TREADY = io_in_x251_TREADY; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 48:23:@36352.4]
  assign x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x250_TDATA = io_in_x250_TDATA; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 49:23:@36360.4]
  assign x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x250_TID = io_in_x250_TID; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 49:23:@36356.4]
  assign x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x250_TDEST = io_in_x250_TDEST; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 49:23:@36355.4]
  assign x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x251_TREADY | x465_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 718:22:@36379.4]
  assign x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_264 & _T_265; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 718:22:@36377.4]
  assign x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x465_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 718:22:@36375.4]
  assign x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x278_ctrchain_io_output_counts_1[12]}},x278_ctrchain_io_output_counts_1}; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 718:22:@36370.4]
  assign x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x278_ctrchain_io_output_counts_0[12]}},x278_ctrchain_io_output_counts_0}; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 718:22:@36369.4]
  assign x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x278_ctrchain_io_output_oobs_0; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 718:22:@36367.4]
  assign x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x278_ctrchain_io_output_oobs_1; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 718:22:@36368.4]
  assign x465_inr_Foreach_SAMPLER_BOX_kernelx465_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x465_inr_Foreach_SAMPLER_BOX.scala 717:18:@36363.4]
endmodule
module x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1( // @[:@36393.2]
  input          clock, // @[:@36394.4]
  input          reset, // @[:@36395.4]
  output         io_in_x251_TVALID, // @[:@36396.4]
  input          io_in_x251_TREADY, // @[:@36396.4]
  output [255:0] io_in_x251_TDATA, // @[:@36396.4]
  input          io_in_x250_TVALID, // @[:@36396.4]
  output         io_in_x250_TREADY, // @[:@36396.4]
  input  [255:0] io_in_x250_TDATA, // @[:@36396.4]
  input  [7:0]   io_in_x250_TID, // @[:@36396.4]
  input  [7:0]   io_in_x250_TDEST, // @[:@36396.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@36396.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@36396.4]
  input          io_sigsIn_smChildAcks_0, // @[:@36396.4]
  input          io_sigsIn_smChildAcks_1, // @[:@36396.4]
  output         io_sigsOut_smDoneIn_0, // @[:@36396.4]
  output         io_sigsOut_smDoneIn_1, // @[:@36396.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@36396.4]
  output         io_sigsOut_smCtrCopyDone_1, // @[:@36396.4]
  input          io_rr // @[:@36396.4]
);
  wire  x253_fifoinraw_0_clock; // @[m_x253_fifoinraw_0.scala 27:17:@36410.4]
  wire  x253_fifoinraw_0_reset; // @[m_x253_fifoinraw_0.scala 27:17:@36410.4]
  wire  x254_fifoinpacked_0_clock; // @[m_x254_fifoinpacked_0.scala 27:17:@36434.4]
  wire  x254_fifoinpacked_0_reset; // @[m_x254_fifoinpacked_0.scala 27:17:@36434.4]
  wire  x254_fifoinpacked_0_io_wPort_0_en_0; // @[m_x254_fifoinpacked_0.scala 27:17:@36434.4]
  wire  x254_fifoinpacked_0_io_full; // @[m_x254_fifoinpacked_0.scala 27:17:@36434.4]
  wire  x254_fifoinpacked_0_io_active_0_in; // @[m_x254_fifoinpacked_0.scala 27:17:@36434.4]
  wire  x254_fifoinpacked_0_io_active_0_out; // @[m_x254_fifoinpacked_0.scala 27:17:@36434.4]
  wire  x255_fifooutraw_0_clock; // @[m_x255_fifooutraw_0.scala 27:17:@36458.4]
  wire  x255_fifooutraw_0_reset; // @[m_x255_fifooutraw_0.scala 27:17:@36458.4]
  wire  x258_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@36482.4]
  wire  x258_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@36482.4]
  wire  x258_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@36482.4]
  wire  x258_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@36482.4]
  wire [12:0] x258_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@36482.4]
  wire [12:0] x258_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@36482.4]
  wire  x258_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@36482.4]
  wire  x258_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@36482.4]
  wire  x258_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@36482.4]
  wire  x274_inr_Foreach_sm_clock; // @[sm_x274_inr_Foreach.scala 32:18:@36542.4]
  wire  x274_inr_Foreach_sm_reset; // @[sm_x274_inr_Foreach.scala 32:18:@36542.4]
  wire  x274_inr_Foreach_sm_io_enable; // @[sm_x274_inr_Foreach.scala 32:18:@36542.4]
  wire  x274_inr_Foreach_sm_io_done; // @[sm_x274_inr_Foreach.scala 32:18:@36542.4]
  wire  x274_inr_Foreach_sm_io_doneLatch; // @[sm_x274_inr_Foreach.scala 32:18:@36542.4]
  wire  x274_inr_Foreach_sm_io_ctrDone; // @[sm_x274_inr_Foreach.scala 32:18:@36542.4]
  wire  x274_inr_Foreach_sm_io_datapathEn; // @[sm_x274_inr_Foreach.scala 32:18:@36542.4]
  wire  x274_inr_Foreach_sm_io_ctrInc; // @[sm_x274_inr_Foreach.scala 32:18:@36542.4]
  wire  x274_inr_Foreach_sm_io_ctrRst; // @[sm_x274_inr_Foreach.scala 32:18:@36542.4]
  wire  x274_inr_Foreach_sm_io_parentAck; // @[sm_x274_inr_Foreach.scala 32:18:@36542.4]
  wire  x274_inr_Foreach_sm_io_backpressure; // @[sm_x274_inr_Foreach.scala 32:18:@36542.4]
  wire  x274_inr_Foreach_sm_io_break; // @[sm_x274_inr_Foreach.scala 32:18:@36542.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@36570.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@36570.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@36570.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@36570.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@36570.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@36616.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@36616.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@36616.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@36616.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@36616.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@36624.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@36624.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@36624.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@36624.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@36624.4]
  wire  x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_clock; // @[sm_x274_inr_Foreach.scala 98:24:@36659.4]
  wire  x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_reset; // @[sm_x274_inr_Foreach.scala 98:24:@36659.4]
  wire  x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_in_x254_fifoinpacked_0_wPort_0_en_0; // @[sm_x274_inr_Foreach.scala 98:24:@36659.4]
  wire  x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_in_x254_fifoinpacked_0_full; // @[sm_x274_inr_Foreach.scala 98:24:@36659.4]
  wire  x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_in_x254_fifoinpacked_0_active_0_in; // @[sm_x274_inr_Foreach.scala 98:24:@36659.4]
  wire  x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_in_x254_fifoinpacked_0_active_0_out; // @[sm_x274_inr_Foreach.scala 98:24:@36659.4]
  wire  x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x274_inr_Foreach.scala 98:24:@36659.4]
  wire  x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x274_inr_Foreach.scala 98:24:@36659.4]
  wire  x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x274_inr_Foreach.scala 98:24:@36659.4]
  wire [31:0] x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x274_inr_Foreach.scala 98:24:@36659.4]
  wire [31:0] x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x274_inr_Foreach.scala 98:24:@36659.4]
  wire  x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x274_inr_Foreach.scala 98:24:@36659.4]
  wire  x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x274_inr_Foreach.scala 98:24:@36659.4]
  wire  x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_rr; // @[sm_x274_inr_Foreach.scala 98:24:@36659.4]
  wire  x466_outr_UnitPipe_sm_clock; // @[sm_x466_outr_UnitPipe.scala 32:18:@36791.4]
  wire  x466_outr_UnitPipe_sm_reset; // @[sm_x466_outr_UnitPipe.scala 32:18:@36791.4]
  wire  x466_outr_UnitPipe_sm_io_enable; // @[sm_x466_outr_UnitPipe.scala 32:18:@36791.4]
  wire  x466_outr_UnitPipe_sm_io_done; // @[sm_x466_outr_UnitPipe.scala 32:18:@36791.4]
  wire  x466_outr_UnitPipe_sm_io_rst; // @[sm_x466_outr_UnitPipe.scala 32:18:@36791.4]
  wire  x466_outr_UnitPipe_sm_io_ctrDone; // @[sm_x466_outr_UnitPipe.scala 32:18:@36791.4]
  wire  x466_outr_UnitPipe_sm_io_ctrInc; // @[sm_x466_outr_UnitPipe.scala 32:18:@36791.4]
  wire  x466_outr_UnitPipe_sm_io_parentAck; // @[sm_x466_outr_UnitPipe.scala 32:18:@36791.4]
  wire  x466_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x466_outr_UnitPipe.scala 32:18:@36791.4]
  wire  x466_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x466_outr_UnitPipe.scala 32:18:@36791.4]
  wire  x466_outr_UnitPipe_sm_io_childAck_0; // @[sm_x466_outr_UnitPipe.scala 32:18:@36791.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@36848.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@36848.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@36848.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@36848.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@36848.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@36856.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@36856.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@36856.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@36856.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@36856.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_clock; // @[sm_x466_outr_UnitPipe.scala 76:24:@36886.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_reset; // @[sm_x466_outr_UnitPipe.scala 76:24:@36886.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x251_TVALID; // @[sm_x466_outr_UnitPipe.scala 76:24:@36886.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x251_TREADY; // @[sm_x466_outr_UnitPipe.scala 76:24:@36886.4]
  wire [255:0] x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x251_TDATA; // @[sm_x466_outr_UnitPipe.scala 76:24:@36886.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x250_TVALID; // @[sm_x466_outr_UnitPipe.scala 76:24:@36886.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x250_TREADY; // @[sm_x466_outr_UnitPipe.scala 76:24:@36886.4]
  wire [255:0] x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x250_TDATA; // @[sm_x466_outr_UnitPipe.scala 76:24:@36886.4]
  wire [7:0] x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x250_TID; // @[sm_x466_outr_UnitPipe.scala 76:24:@36886.4]
  wire [7:0] x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x250_TDEST; // @[sm_x466_outr_UnitPipe.scala 76:24:@36886.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x466_outr_UnitPipe.scala 76:24:@36886.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x466_outr_UnitPipe.scala 76:24:@36886.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x466_outr_UnitPipe.scala 76:24:@36886.4]
  wire  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_rr; // @[sm_x466_outr_UnitPipe.scala 76:24:@36886.4]
  wire  _T_254; // @[package.scala 96:25:@36575.4 package.scala 96:25:@36576.4]
  wire  _T_260; // @[implicits.scala 47:10:@36579.4]
  wire  _T_261; // @[sm_x467_outr_UnitPipe.scala 70:41:@36580.4]
  wire  _T_262; // @[sm_x467_outr_UnitPipe.scala 70:78:@36581.4]
  wire  _T_263; // @[sm_x467_outr_UnitPipe.scala 70:76:@36582.4]
  wire  _T_275; // @[package.scala 96:25:@36621.4 package.scala 96:25:@36622.4]
  wire  _T_281; // @[package.scala 96:25:@36629.4 package.scala 96:25:@36630.4]
  wire  _T_284; // @[SpatialBlocks.scala 138:93:@36632.4]
  wire  _T_286; // @[SpatialBlocks.scala 157:36:@36641.4]
  wire  _T_287; // @[SpatialBlocks.scala 157:78:@36642.4]
  wire  _T_354; // @[package.scala 100:49:@36819.4]
  reg  _T_357; // @[package.scala 48:56:@36820.4]
  reg [31:0] _RAND_0;
  wire  _T_371; // @[package.scala 96:25:@36853.4 package.scala 96:25:@36854.4]
  wire  _T_377; // @[package.scala 96:25:@36861.4 package.scala 96:25:@36862.4]
  wire  _T_380; // @[SpatialBlocks.scala 138:93:@36864.4]
  x253_fifoinraw_0 x253_fifoinraw_0 ( // @[m_x253_fifoinraw_0.scala 27:17:@36410.4]
    .clock(x253_fifoinraw_0_clock),
    .reset(x253_fifoinraw_0_reset)
  );
  x254_fifoinpacked_0 x254_fifoinpacked_0 ( // @[m_x254_fifoinpacked_0.scala 27:17:@36434.4]
    .clock(x254_fifoinpacked_0_clock),
    .reset(x254_fifoinpacked_0_reset),
    .io_wPort_0_en_0(x254_fifoinpacked_0_io_wPort_0_en_0),
    .io_full(x254_fifoinpacked_0_io_full),
    .io_active_0_in(x254_fifoinpacked_0_io_active_0_in),
    .io_active_0_out(x254_fifoinpacked_0_io_active_0_out)
  );
  x253_fifoinraw_0 x255_fifooutraw_0 ( // @[m_x255_fifooutraw_0.scala 27:17:@36458.4]
    .clock(x255_fifooutraw_0_clock),
    .reset(x255_fifooutraw_0_reset)
  );
  x258_ctrchain x258_ctrchain ( // @[SpatialBlocks.scala 37:22:@36482.4]
    .clock(x258_ctrchain_clock),
    .reset(x258_ctrchain_reset),
    .io_input_reset(x258_ctrchain_io_input_reset),
    .io_input_enable(x258_ctrchain_io_input_enable),
    .io_output_counts_1(x258_ctrchain_io_output_counts_1),
    .io_output_counts_0(x258_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x258_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x258_ctrchain_io_output_oobs_1),
    .io_output_done(x258_ctrchain_io_output_done)
  );
  x274_inr_Foreach_sm x274_inr_Foreach_sm ( // @[sm_x274_inr_Foreach.scala 32:18:@36542.4]
    .clock(x274_inr_Foreach_sm_clock),
    .reset(x274_inr_Foreach_sm_reset),
    .io_enable(x274_inr_Foreach_sm_io_enable),
    .io_done(x274_inr_Foreach_sm_io_done),
    .io_doneLatch(x274_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x274_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x274_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x274_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x274_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x274_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x274_inr_Foreach_sm_io_backpressure),
    .io_break(x274_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@36570.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@36616.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@36624.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x274_inr_Foreach_kernelx274_inr_Foreach_concrete1 x274_inr_Foreach_kernelx274_inr_Foreach_concrete1 ( // @[sm_x274_inr_Foreach.scala 98:24:@36659.4]
    .clock(x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_clock),
    .reset(x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_reset),
    .io_in_x254_fifoinpacked_0_wPort_0_en_0(x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_in_x254_fifoinpacked_0_wPort_0_en_0),
    .io_in_x254_fifoinpacked_0_full(x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_in_x254_fifoinpacked_0_full),
    .io_in_x254_fifoinpacked_0_active_0_in(x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_in_x254_fifoinpacked_0_active_0_in),
    .io_in_x254_fifoinpacked_0_active_0_out(x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_in_x254_fifoinpacked_0_active_0_out),
    .io_sigsIn_backpressure(x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_rr)
  );
  RootController_sm x466_outr_UnitPipe_sm ( // @[sm_x466_outr_UnitPipe.scala 32:18:@36791.4]
    .clock(x466_outr_UnitPipe_sm_clock),
    .reset(x466_outr_UnitPipe_sm_reset),
    .io_enable(x466_outr_UnitPipe_sm_io_enable),
    .io_done(x466_outr_UnitPipe_sm_io_done),
    .io_rst(x466_outr_UnitPipe_sm_io_rst),
    .io_ctrDone(x466_outr_UnitPipe_sm_io_ctrDone),
    .io_ctrInc(x466_outr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x466_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x466_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x466_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x466_outr_UnitPipe_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@36848.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@36856.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1 x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1 ( // @[sm_x466_outr_UnitPipe.scala 76:24:@36886.4]
    .clock(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_clock),
    .reset(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_reset),
    .io_in_x251_TVALID(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x251_TVALID),
    .io_in_x251_TREADY(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x251_TREADY),
    .io_in_x251_TDATA(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x251_TDATA),
    .io_in_x250_TVALID(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x250_TVALID),
    .io_in_x250_TREADY(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x250_TREADY),
    .io_in_x250_TDATA(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x250_TDATA),
    .io_in_x250_TID(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x250_TID),
    .io_in_x250_TDEST(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x250_TDEST),
    .io_sigsIn_smEnableOuts_0(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_254 = RetimeWrapper_io_out; // @[package.scala 96:25:@36575.4 package.scala 96:25:@36576.4]
  assign _T_260 = x254_fifoinpacked_0_io_full; // @[implicits.scala 47:10:@36579.4]
  assign _T_261 = ~ _T_260; // @[sm_x467_outr_UnitPipe.scala 70:41:@36580.4]
  assign _T_262 = ~ x254_fifoinpacked_0_io_active_0_out; // @[sm_x467_outr_UnitPipe.scala 70:78:@36581.4]
  assign _T_263 = _T_261 | _T_262; // @[sm_x467_outr_UnitPipe.scala 70:76:@36582.4]
  assign _T_275 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@36621.4 package.scala 96:25:@36622.4]
  assign _T_281 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@36629.4 package.scala 96:25:@36630.4]
  assign _T_284 = ~ _T_281; // @[SpatialBlocks.scala 138:93:@36632.4]
  assign _T_286 = x274_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@36641.4]
  assign _T_287 = ~ x274_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@36642.4]
  assign _T_354 = x466_outr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@36819.4]
  assign _T_371 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@36853.4 package.scala 96:25:@36854.4]
  assign _T_377 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@36861.4 package.scala 96:25:@36862.4]
  assign _T_380 = ~ _T_377; // @[SpatialBlocks.scala 138:93:@36864.4]
  assign io_in_x251_TVALID = x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x251_TVALID; // @[sm_x466_outr_UnitPipe.scala 48:23:@36943.4]
  assign io_in_x251_TDATA = x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x251_TDATA; // @[sm_x466_outr_UnitPipe.scala 48:23:@36941.4]
  assign io_in_x250_TREADY = x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x250_TREADY; // @[sm_x466_outr_UnitPipe.scala 49:23:@36951.4]
  assign io_sigsOut_smDoneIn_0 = x274_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@36639.4]
  assign io_sigsOut_smDoneIn_1 = x466_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@36871.4]
  assign io_sigsOut_smCtrCopyDone_0 = x274_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@36658.4]
  assign io_sigsOut_smCtrCopyDone_1 = x466_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@36885.4]
  assign x253_fifoinraw_0_clock = clock; // @[:@36411.4]
  assign x253_fifoinraw_0_reset = reset; // @[:@36412.4]
  assign x254_fifoinpacked_0_clock = clock; // @[:@36435.4]
  assign x254_fifoinpacked_0_reset = reset; // @[:@36436.4]
  assign x254_fifoinpacked_0_io_wPort_0_en_0 = x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_in_x254_fifoinpacked_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@36719.4]
  assign x254_fifoinpacked_0_io_active_0_in = x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_in_x254_fifoinpacked_0_active_0_in; // @[MemInterfaceType.scala 167:86:@36718.4]
  assign x255_fifooutraw_0_clock = clock; // @[:@36459.4]
  assign x255_fifooutraw_0_reset = reset; // @[:@36460.4]
  assign x258_ctrchain_clock = clock; // @[:@36483.4]
  assign x258_ctrchain_reset = reset; // @[:@36484.4]
  assign x258_ctrchain_io_input_reset = x274_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@36657.4]
  assign x258_ctrchain_io_input_enable = x274_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@36609.4 SpatialBlocks.scala 159:42:@36656.4]
  assign x274_inr_Foreach_sm_clock = clock; // @[:@36543.4]
  assign x274_inr_Foreach_sm_reset = reset; // @[:@36544.4]
  assign x274_inr_Foreach_sm_io_enable = _T_275 & _T_284; // @[SpatialBlocks.scala 140:18:@36636.4]
  assign x274_inr_Foreach_sm_io_ctrDone = io_rr ? _T_254 : 1'h0; // @[sm_x467_outr_UnitPipe.scala 69:38:@36578.4]
  assign x274_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@36638.4]
  assign x274_inr_Foreach_sm_io_backpressure = _T_263 | x274_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@36610.4]
  assign x274_inr_Foreach_sm_io_break = 1'h0; // @[sm_x467_outr_UnitPipe.scala 73:36:@36588.4]
  assign RetimeWrapper_clock = clock; // @[:@36571.4]
  assign RetimeWrapper_reset = reset; // @[:@36572.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@36574.4]
  assign RetimeWrapper_io_in = x258_ctrchain_io_output_done; // @[package.scala 94:16:@36573.4]
  assign RetimeWrapper_1_clock = clock; // @[:@36617.4]
  assign RetimeWrapper_1_reset = reset; // @[:@36618.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@36620.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@36619.4]
  assign RetimeWrapper_2_clock = clock; // @[:@36625.4]
  assign RetimeWrapper_2_reset = reset; // @[:@36626.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@36628.4]
  assign RetimeWrapper_2_io_in = x274_inr_Foreach_sm_io_done; // @[package.scala 94:16:@36627.4]
  assign x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_clock = clock; // @[:@36660.4]
  assign x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_reset = reset; // @[:@36661.4]
  assign x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_in_x254_fifoinpacked_0_full = x254_fifoinpacked_0_io_full; // @[MemInterfaceType.scala 159:15:@36713.4]
  assign x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_in_x254_fifoinpacked_0_active_0_out = x254_fifoinpacked_0_io_active_0_out; // @[MemInterfaceType.scala 158:75:@36712.4]
  assign x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_263 | x274_inr_Foreach_sm_io_doneLatch; // @[sm_x274_inr_Foreach.scala 103:22:@36742.4]
  assign x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_286 & _T_287; // @[sm_x274_inr_Foreach.scala 103:22:@36740.4]
  assign x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_break = x274_inr_Foreach_sm_io_break; // @[sm_x274_inr_Foreach.scala 103:22:@36738.4]
  assign x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x258_ctrchain_io_output_counts_1[12]}},x258_ctrchain_io_output_counts_1}; // @[sm_x274_inr_Foreach.scala 103:22:@36733.4]
  assign x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x258_ctrchain_io_output_counts_0[12]}},x258_ctrchain_io_output_counts_0}; // @[sm_x274_inr_Foreach.scala 103:22:@36732.4]
  assign x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x258_ctrchain_io_output_oobs_0; // @[sm_x274_inr_Foreach.scala 103:22:@36730.4]
  assign x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x258_ctrchain_io_output_oobs_1; // @[sm_x274_inr_Foreach.scala 103:22:@36731.4]
  assign x274_inr_Foreach_kernelx274_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x274_inr_Foreach.scala 102:18:@36726.4]
  assign x466_outr_UnitPipe_sm_clock = clock; // @[:@36792.4]
  assign x466_outr_UnitPipe_sm_reset = reset; // @[:@36793.4]
  assign x466_outr_UnitPipe_sm_io_enable = _T_371 & _T_380; // @[SpatialBlocks.scala 140:18:@36868.4]
  assign x466_outr_UnitPipe_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 134:15:@36843.4]
  assign x466_outr_UnitPipe_sm_io_ctrDone = x466_outr_UnitPipe_sm_io_ctrInc & _T_357; // @[sm_x467_outr_UnitPipe.scala 78:40:@36823.4]
  assign x466_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@36870.4]
  assign x466_outr_UnitPipe_sm_io_doneIn_0 = x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@36840.4]
  assign RetimeWrapper_3_clock = clock; // @[:@36849.4]
  assign RetimeWrapper_3_reset = reset; // @[:@36850.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@36852.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@36851.4]
  assign RetimeWrapper_4_clock = clock; // @[:@36857.4]
  assign RetimeWrapper_4_reset = reset; // @[:@36858.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@36860.4]
  assign RetimeWrapper_4_io_in = x466_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@36859.4]
  assign x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_clock = clock; // @[:@36887.4]
  assign x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_reset = reset; // @[:@36888.4]
  assign x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x251_TREADY = io_in_x251_TREADY; // @[sm_x466_outr_UnitPipe.scala 48:23:@36942.4]
  assign x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x250_TVALID = io_in_x250_TVALID; // @[sm_x466_outr_UnitPipe.scala 49:23:@36952.4]
  assign x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x250_TDATA = io_in_x250_TDATA; // @[sm_x466_outr_UnitPipe.scala 49:23:@36950.4]
  assign x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x250_TID = io_in_x250_TID; // @[sm_x466_outr_UnitPipe.scala 49:23:@36946.4]
  assign x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_in_x250_TDEST = io_in_x250_TDEST; // @[sm_x466_outr_UnitPipe.scala 49:23:@36945.4]
  assign x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x466_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x466_outr_UnitPipe.scala 81:22:@36961.4]
  assign x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x466_outr_UnitPipe_sm_io_childAck_0; // @[sm_x466_outr_UnitPipe.scala 81:22:@36959.4]
  assign x466_outr_UnitPipe_kernelx466_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x466_outr_UnitPipe.scala 80:18:@36953.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_357 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_357 <= 1'h0;
    end else begin
      _T_357 <= _T_354;
    end
  end
endmodule
module x489_outr_UnitPipe_sm( // @[:@37450.2]
  input   clock, // @[:@37451.4]
  input   reset, // @[:@37452.4]
  input   io_enable, // @[:@37453.4]
  output  io_done, // @[:@37453.4]
  input   io_parentAck, // @[:@37453.4]
  input   io_doneIn_0, // @[:@37453.4]
  input   io_doneIn_1, // @[:@37453.4]
  input   io_doneIn_2, // @[:@37453.4]
  output  io_enableOut_0, // @[:@37453.4]
  output  io_enableOut_1, // @[:@37453.4]
  output  io_enableOut_2, // @[:@37453.4]
  output  io_childAck_0, // @[:@37453.4]
  output  io_childAck_1, // @[:@37453.4]
  output  io_childAck_2, // @[:@37453.4]
  input   io_ctrCopyDone_0, // @[:@37453.4]
  input   io_ctrCopyDone_1, // @[:@37453.4]
  input   io_ctrCopyDone_2 // @[:@37453.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@37456.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@37456.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@37456.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@37456.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@37456.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@37456.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@37459.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@37459.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@37459.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@37459.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@37459.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@37459.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@37462.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@37462.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@37462.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@37462.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@37462.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@37462.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@37465.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@37465.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@37465.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@37465.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@37465.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@37465.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@37468.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@37468.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@37468.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@37468.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@37468.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@37468.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@37471.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@37471.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@37471.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@37471.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@37471.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@37471.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@37512.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@37512.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@37512.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@37512.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@37512.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@37512.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@37515.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@37515.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@37515.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@37515.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@37515.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@37515.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@37518.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@37518.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@37518.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@37518.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@37518.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@37518.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@37569.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@37569.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@37569.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@37569.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@37569.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@37583.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@37583.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@37583.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@37583.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@37583.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@37601.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@37601.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@37601.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@37601.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@37601.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@37638.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@37638.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@37638.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@37638.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@37638.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@37652.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@37652.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@37652.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@37652.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@37652.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@37670.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@37670.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@37670.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@37670.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@37670.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@37707.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@37707.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@37707.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@37707.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@37707.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@37721.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@37721.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@37721.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@37721.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@37721.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@37739.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@37739.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@37739.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@37739.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@37739.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@37796.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@37796.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@37796.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@37796.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@37796.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@37813.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@37813.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@37813.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@37813.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@37813.4]
  wire  _T_77; // @[Controllers.scala 80:47:@37474.4]
  wire  allDone; // @[Controllers.scala 80:47:@37475.4]
  wire  _T_151; // @[Controllers.scala 165:35:@37553.4]
  wire  _T_153; // @[Controllers.scala 165:60:@37554.4]
  wire  _T_154; // @[Controllers.scala 165:58:@37555.4]
  wire  _T_156; // @[Controllers.scala 165:76:@37556.4]
  wire  _T_157; // @[Controllers.scala 165:74:@37557.4]
  wire  _T_161; // @[Controllers.scala 165:109:@37560.4]
  wire  _T_164; // @[Controllers.scala 165:141:@37562.4]
  wire  _T_172; // @[package.scala 96:25:@37574.4 package.scala 96:25:@37575.4]
  wire  _T_176; // @[Controllers.scala 167:54:@37577.4]
  wire  _T_177; // @[Controllers.scala 167:52:@37578.4]
  wire  _T_184; // @[package.scala 96:25:@37588.4 package.scala 96:25:@37589.4]
  wire  _T_202; // @[package.scala 96:25:@37606.4 package.scala 96:25:@37607.4]
  wire  _T_206; // @[Controllers.scala 169:67:@37609.4]
  wire  _T_207; // @[Controllers.scala 169:86:@37610.4]
  wire  _T_219; // @[Controllers.scala 165:35:@37622.4]
  wire  _T_221; // @[Controllers.scala 165:60:@37623.4]
  wire  _T_222; // @[Controllers.scala 165:58:@37624.4]
  wire  _T_224; // @[Controllers.scala 165:76:@37625.4]
  wire  _T_225; // @[Controllers.scala 165:74:@37626.4]
  wire  _T_229; // @[Controllers.scala 165:109:@37629.4]
  wire  _T_232; // @[Controllers.scala 165:141:@37631.4]
  wire  _T_240; // @[package.scala 96:25:@37643.4 package.scala 96:25:@37644.4]
  wire  _T_244; // @[Controllers.scala 167:54:@37646.4]
  wire  _T_245; // @[Controllers.scala 167:52:@37647.4]
  wire  _T_252; // @[package.scala 96:25:@37657.4 package.scala 96:25:@37658.4]
  wire  _T_270; // @[package.scala 96:25:@37675.4 package.scala 96:25:@37676.4]
  wire  _T_274; // @[Controllers.scala 169:67:@37678.4]
  wire  _T_275; // @[Controllers.scala 169:86:@37679.4]
  wire  _T_287; // @[Controllers.scala 165:35:@37691.4]
  wire  _T_289; // @[Controllers.scala 165:60:@37692.4]
  wire  _T_290; // @[Controllers.scala 165:58:@37693.4]
  wire  _T_292; // @[Controllers.scala 165:76:@37694.4]
  wire  _T_293; // @[Controllers.scala 165:74:@37695.4]
  wire  _T_297; // @[Controllers.scala 165:109:@37698.4]
  wire  _T_300; // @[Controllers.scala 165:141:@37700.4]
  wire  _T_308; // @[package.scala 96:25:@37712.4 package.scala 96:25:@37713.4]
  wire  _T_312; // @[Controllers.scala 167:54:@37715.4]
  wire  _T_313; // @[Controllers.scala 167:52:@37716.4]
  wire  _T_320; // @[package.scala 96:25:@37726.4 package.scala 96:25:@37727.4]
  wire  _T_338; // @[package.scala 96:25:@37744.4 package.scala 96:25:@37745.4]
  wire  _T_342; // @[Controllers.scala 169:67:@37747.4]
  wire  _T_343; // @[Controllers.scala 169:86:@37748.4]
  wire  _T_358; // @[Controllers.scala 213:68:@37766.4]
  wire  _T_360; // @[Controllers.scala 213:90:@37768.4]
  wire  _T_362; // @[Controllers.scala 213:132:@37770.4]
  wire  _T_366; // @[Controllers.scala 213:68:@37775.4]
  wire  _T_368; // @[Controllers.scala 213:90:@37777.4]
  wire  _T_374; // @[Controllers.scala 213:68:@37783.4]
  wire  _T_376; // @[Controllers.scala 213:90:@37785.4]
  wire  _T_383; // @[package.scala 100:49:@37791.4]
  reg  _T_386; // @[package.scala 48:56:@37792.4]
  reg [31:0] _RAND_0;
  wire  _T_387; // @[package.scala 100:41:@37794.4]
  reg  _T_400; // @[package.scala 48:56:@37810.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@37456.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@37459.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@37462.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@37465.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@37468.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@37471.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@37512.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@37515.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@37518.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@37569.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@37583.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@37601.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@37638.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@37652.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@37670.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@37707.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@37721.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@37739.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@37796.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@37813.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@37474.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@37475.4]
  assign _T_151 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@37553.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@37554.4]
  assign _T_154 = _T_151 & _T_153; // @[Controllers.scala 165:58:@37555.4]
  assign _T_156 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@37556.4]
  assign _T_157 = _T_154 & _T_156; // @[Controllers.scala 165:74:@37557.4]
  assign _T_161 = _T_157 & io_enable; // @[Controllers.scala 165:109:@37560.4]
  assign _T_164 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@37562.4]
  assign _T_172 = RetimeWrapper_io_out; // @[package.scala 96:25:@37574.4 package.scala 96:25:@37575.4]
  assign _T_176 = _T_172 == 1'h0; // @[Controllers.scala 167:54:@37577.4]
  assign _T_177 = io_doneIn_0 | _T_176; // @[Controllers.scala 167:52:@37578.4]
  assign _T_184 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@37588.4 package.scala 96:25:@37589.4]
  assign _T_202 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@37606.4 package.scala 96:25:@37607.4]
  assign _T_206 = _T_202 == 1'h0; // @[Controllers.scala 169:67:@37609.4]
  assign _T_207 = _T_206 & io_enable; // @[Controllers.scala 169:86:@37610.4]
  assign _T_219 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@37622.4]
  assign _T_221 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@37623.4]
  assign _T_222 = _T_219 & _T_221; // @[Controllers.scala 165:58:@37624.4]
  assign _T_224 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@37625.4]
  assign _T_225 = _T_222 & _T_224; // @[Controllers.scala 165:74:@37626.4]
  assign _T_229 = _T_225 & io_enable; // @[Controllers.scala 165:109:@37629.4]
  assign _T_232 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@37631.4]
  assign _T_240 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@37643.4 package.scala 96:25:@37644.4]
  assign _T_244 = _T_240 == 1'h0; // @[Controllers.scala 167:54:@37646.4]
  assign _T_245 = io_doneIn_1 | _T_244; // @[Controllers.scala 167:52:@37647.4]
  assign _T_252 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@37657.4 package.scala 96:25:@37658.4]
  assign _T_270 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@37675.4 package.scala 96:25:@37676.4]
  assign _T_274 = _T_270 == 1'h0; // @[Controllers.scala 169:67:@37678.4]
  assign _T_275 = _T_274 & io_enable; // @[Controllers.scala 169:86:@37679.4]
  assign _T_287 = ~ iterDone_2_io_output; // @[Controllers.scala 165:35:@37691.4]
  assign _T_289 = io_doneIn_2 == 1'h0; // @[Controllers.scala 165:60:@37692.4]
  assign _T_290 = _T_287 & _T_289; // @[Controllers.scala 165:58:@37693.4]
  assign _T_292 = done_2_io_output == 1'h0; // @[Controllers.scala 165:76:@37694.4]
  assign _T_293 = _T_290 & _T_292; // @[Controllers.scala 165:74:@37695.4]
  assign _T_297 = _T_293 & io_enable; // @[Controllers.scala 165:109:@37698.4]
  assign _T_300 = io_ctrCopyDone_2 == 1'h0; // @[Controllers.scala 165:141:@37700.4]
  assign _T_308 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@37712.4 package.scala 96:25:@37713.4]
  assign _T_312 = _T_308 == 1'h0; // @[Controllers.scala 167:54:@37715.4]
  assign _T_313 = io_doneIn_2 | _T_312; // @[Controllers.scala 167:52:@37716.4]
  assign _T_320 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@37726.4 package.scala 96:25:@37727.4]
  assign _T_338 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@37744.4 package.scala 96:25:@37745.4]
  assign _T_342 = _T_338 == 1'h0; // @[Controllers.scala 169:67:@37747.4]
  assign _T_343 = _T_342 & io_enable; // @[Controllers.scala 169:86:@37748.4]
  assign _T_358 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@37766.4]
  assign _T_360 = _T_358 & _T_151; // @[Controllers.scala 213:90:@37768.4]
  assign _T_362 = ~ allDone; // @[Controllers.scala 213:132:@37770.4]
  assign _T_366 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@37775.4]
  assign _T_368 = _T_366 & _T_219; // @[Controllers.scala 213:90:@37777.4]
  assign _T_374 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@37783.4]
  assign _T_376 = _T_374 & _T_287; // @[Controllers.scala 213:90:@37785.4]
  assign _T_383 = allDone == 1'h0; // @[package.scala 100:49:@37791.4]
  assign _T_387 = allDone & _T_386; // @[package.scala 100:41:@37794.4]
  assign io_done = RetimeWrapper_10_io_out; // @[Controllers.scala 245:13:@37820.4]
  assign io_enableOut_0 = _T_360 & _T_362; // @[Controllers.scala 213:55:@37774.4]
  assign io_enableOut_1 = _T_368 & _T_362; // @[Controllers.scala 213:55:@37782.4]
  assign io_enableOut_2 = _T_376 & _T_362; // @[Controllers.scala 213:55:@37790.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@37761.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@37763.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@37765.4]
  assign active_0_clock = clock; // @[:@37457.4]
  assign active_0_reset = reset; // @[:@37458.4]
  assign active_0_io_input_set = _T_161 & _T_164; // @[Controllers.scala 165:32:@37564.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@37568.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@37478.4]
  assign active_1_clock = clock; // @[:@37460.4]
  assign active_1_reset = reset; // @[:@37461.4]
  assign active_1_io_input_set = _T_229 & _T_232; // @[Controllers.scala 165:32:@37633.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@37637.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@37479.4]
  assign active_2_clock = clock; // @[:@37463.4]
  assign active_2_reset = reset; // @[:@37464.4]
  assign active_2_io_input_set = _T_297 & _T_300; // @[Controllers.scala 165:32:@37702.4]
  assign active_2_io_input_reset = io_ctrCopyDone_2 | io_parentAck; // @[Controllers.scala 166:34:@37706.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@37480.4]
  assign done_0_clock = clock; // @[:@37466.4]
  assign done_0_reset = reset; // @[:@37467.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_207; // @[Controllers.scala 169:30:@37614.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@37492.4 Controllers.scala 170:32:@37621.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@37481.4]
  assign done_1_clock = clock; // @[:@37469.4]
  assign done_1_reset = reset; // @[:@37470.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_275; // @[Controllers.scala 169:30:@37683.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@37501.4 Controllers.scala 170:32:@37690.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@37482.4]
  assign done_2_clock = clock; // @[:@37472.4]
  assign done_2_reset = reset; // @[:@37473.4]
  assign done_2_io_input_set = io_ctrCopyDone_2 | _T_343; // @[Controllers.scala 169:30:@37752.4]
  assign done_2_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@37510.4 Controllers.scala 170:32:@37759.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@37483.4]
  assign iterDone_0_clock = clock; // @[:@37513.4]
  assign iterDone_0_reset = reset; // @[:@37514.4]
  assign iterDone_0_io_input_set = _T_177 & io_enable; // @[Controllers.scala 167:34:@37582.4]
  assign iterDone_0_io_input_reset = _T_184 | io_parentAck; // @[Controllers.scala 92:37:@37532.4 Controllers.scala 168:36:@37598.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@37521.4]
  assign iterDone_1_clock = clock; // @[:@37516.4]
  assign iterDone_1_reset = reset; // @[:@37517.4]
  assign iterDone_1_io_input_set = _T_245 & io_enable; // @[Controllers.scala 167:34:@37651.4]
  assign iterDone_1_io_input_reset = _T_252 | io_parentAck; // @[Controllers.scala 92:37:@37541.4 Controllers.scala 168:36:@37667.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@37522.4]
  assign iterDone_2_clock = clock; // @[:@37519.4]
  assign iterDone_2_reset = reset; // @[:@37520.4]
  assign iterDone_2_io_input_set = _T_313 & io_enable; // @[Controllers.scala 167:34:@37720.4]
  assign iterDone_2_io_input_reset = _T_320 | io_parentAck; // @[Controllers.scala 92:37:@37550.4 Controllers.scala 168:36:@37736.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@37523.4]
  assign RetimeWrapper_clock = clock; // @[:@37570.4]
  assign RetimeWrapper_reset = reset; // @[:@37571.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@37573.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@37572.4]
  assign RetimeWrapper_1_clock = clock; // @[:@37584.4]
  assign RetimeWrapper_1_reset = reset; // @[:@37585.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@37587.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@37586.4]
  assign RetimeWrapper_2_clock = clock; // @[:@37602.4]
  assign RetimeWrapper_2_reset = reset; // @[:@37603.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@37605.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@37604.4]
  assign RetimeWrapper_3_clock = clock; // @[:@37639.4]
  assign RetimeWrapper_3_reset = reset; // @[:@37640.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@37642.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@37641.4]
  assign RetimeWrapper_4_clock = clock; // @[:@37653.4]
  assign RetimeWrapper_4_reset = reset; // @[:@37654.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@37656.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@37655.4]
  assign RetimeWrapper_5_clock = clock; // @[:@37671.4]
  assign RetimeWrapper_5_reset = reset; // @[:@37672.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@37674.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@37673.4]
  assign RetimeWrapper_6_clock = clock; // @[:@37708.4]
  assign RetimeWrapper_6_reset = reset; // @[:@37709.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@37711.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@37710.4]
  assign RetimeWrapper_7_clock = clock; // @[:@37722.4]
  assign RetimeWrapper_7_reset = reset; // @[:@37723.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@37725.4]
  assign RetimeWrapper_7_io_in = io_doneIn_2; // @[package.scala 94:16:@37724.4]
  assign RetimeWrapper_8_clock = clock; // @[:@37740.4]
  assign RetimeWrapper_8_reset = reset; // @[:@37741.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@37743.4]
  assign RetimeWrapper_8_io_in = 1'h1; // @[package.scala 94:16:@37742.4]
  assign RetimeWrapper_9_clock = clock; // @[:@37797.4]
  assign RetimeWrapper_9_reset = reset; // @[:@37798.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@37800.4]
  assign RetimeWrapper_9_io_in = _T_387 | io_parentAck; // @[package.scala 94:16:@37799.4]
  assign RetimeWrapper_10_clock = clock; // @[:@37814.4]
  assign RetimeWrapper_10_reset = reset; // @[:@37815.4]
  assign RetimeWrapper_10_io_flow = io_enable; // @[package.scala 95:18:@37817.4]
  assign RetimeWrapper_10_io_in = allDone & _T_400; // @[package.scala 94:16:@37816.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_386 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_400 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_386 <= 1'h0;
    end else begin
      _T_386 <= _T_383;
    end
    if (reset) begin
      _T_400 <= 1'h0;
    end else begin
      _T_400 <= _T_383;
    end
  end
endmodule
module x475_inr_UnitPipe_sm( // @[:@37993.2]
  input   clock, // @[:@37994.4]
  input   reset, // @[:@37995.4]
  input   io_enable, // @[:@37996.4]
  output  io_done, // @[:@37996.4]
  output  io_doneLatch, // @[:@37996.4]
  input   io_ctrDone, // @[:@37996.4]
  output  io_datapathEn, // @[:@37996.4]
  output  io_ctrInc, // @[:@37996.4]
  input   io_parentAck, // @[:@37996.4]
  input   io_backpressure // @[:@37996.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@37998.4]
  wire  active_reset; // @[Controllers.scala 261:22:@37998.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@37998.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@37998.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@37998.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@37998.4]
  wire  done_clock; // @[Controllers.scala 262:20:@38001.4]
  wire  done_reset; // @[Controllers.scala 262:20:@38001.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@38001.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@38001.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@38001.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@38001.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@38055.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@38055.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@38055.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@38055.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@38055.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@38063.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@38063.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@38063.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@38063.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@38063.4]
  wire  _T_80; // @[Controllers.scala 264:48:@38006.4]
  wire  _T_81; // @[Controllers.scala 264:46:@38007.4]
  wire  _T_82; // @[Controllers.scala 264:62:@38008.4]
  wire  _T_83; // @[Controllers.scala 264:60:@38009.4]
  wire  _T_100; // @[package.scala 100:49:@38026.4]
  reg  _T_103; // @[package.scala 48:56:@38027.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 100:49:@38035.4]
  wire  _T_116; // @[Controllers.scala 283:41:@38043.4]
  wire  _T_117; // @[Controllers.scala 283:59:@38044.4]
  wire  _T_119; // @[Controllers.scala 284:37:@38047.4]
  reg  _T_125; // @[package.scala 48:56:@38051.4]
  reg [31:0] _RAND_1;
  reg  _T_142; // @[Controllers.scala 291:31:@38073.4]
  reg [31:0] _RAND_2;
  reg  _T_149; // @[package.scala 48:56:@38076.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:41:@38078.4]
  wire  _T_152; // @[Controllers.scala 292:61:@38079.4]
  wire  _T_153; // @[Controllers.scala 292:24:@38080.4]
  SRFF active ( // @[Controllers.scala 261:22:@37998.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@38001.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@38055.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@38063.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@38006.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@38007.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@38008.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@38009.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@38026.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 100:49:@38035.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@38043.4]
  assign _T_117 = _T_116 & io_enable; // @[Controllers.scala 283:59:@38044.4]
  assign _T_119 = active_io_output & io_enable; // @[Controllers.scala 284:37:@38047.4]
  assign _T_150 = done_io_output & _T_149; // @[package.scala 100:41:@38078.4]
  assign _T_152 = _T_150 ? 1'h1 : _T_142; // @[Controllers.scala 292:61:@38079.4]
  assign _T_153 = io_parentAck ? 1'h0 : _T_152; // @[Controllers.scala 292:24:@38080.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@38054.4]
  assign io_doneLatch = _T_142; // @[Controllers.scala 293:18:@38082.4]
  assign io_datapathEn = _T_117 & io_backpressure; // @[Controllers.scala 283:21:@38046.4]
  assign io_ctrInc = _T_119 & io_backpressure; // @[Controllers.scala 284:17:@38049.4]
  assign active_clock = clock; // @[:@37999.4]
  assign active_reset = reset; // @[:@38000.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@38011.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@38015.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@38016.4]
  assign done_clock = clock; // @[:@38002.4]
  assign done_reset = reset; // @[:@38003.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@38031.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@38024.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@38025.4]
  assign RetimeWrapper_clock = clock; // @[:@38056.4]
  assign RetimeWrapper_reset = reset; // @[:@38057.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@38059.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@38058.4]
  assign RetimeWrapper_1_clock = clock; // @[:@38064.4]
  assign RetimeWrapper_1_reset = reset; // @[:@38065.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@38067.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 94:16:@38066.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_125 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_142 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_149 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_142 <= 1'h0;
      end else begin
        if (_T_150) begin
          _T_142 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_108;
    end
  end
endmodule
module x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1( // @[:@38157.2]
  output        io_in_x468_valid, // @[:@38160.4]
  output [63:0] io_in_x468_bits_addr, // @[:@38160.4]
  output [31:0] io_in_x468_bits_size, // @[:@38160.4]
  input  [63:0] io_in_x248_outdram_number, // @[:@38160.4]
  input         io_sigsIn_backpressure, // @[:@38160.4]
  input         io_sigsIn_datapathEn, // @[:@38160.4]
  input         io_rr // @[:@38160.4]
);
  wire [96:0] x472_tuple; // @[Cat.scala 30:58:@38174.4]
  wire  _T_135; // @[implicits.scala 55:10:@38177.4]
  assign x472_tuple = {33'h7e9000,io_in_x248_outdram_number}; // @[Cat.scala 30:58:@38174.4]
  assign _T_135 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@38177.4]
  assign io_in_x468_valid = _T_135 & io_sigsIn_backpressure; // @[sm_x475_inr_UnitPipe.scala 65:18:@38180.4]
  assign io_in_x468_bits_addr = x472_tuple[63:0]; // @[sm_x475_inr_UnitPipe.scala 66:22:@38182.4]
  assign io_in_x468_bits_size = x472_tuple[95:64]; // @[sm_x475_inr_UnitPipe.scala 67:22:@38184.4]
endmodule
module FF_13( // @[:@38186.2]
  input         clock, // @[:@38187.4]
  input         reset, // @[:@38188.4]
  output [22:0] io_rPort_0_output_0, // @[:@38189.4]
  input  [22:0] io_wPort_0_data_0, // @[:@38189.4]
  input         io_wPort_0_reset, // @[:@38189.4]
  input         io_wPort_0_en_0 // @[:@38189.4]
);
  reg [22:0] ff; // @[MemPrimitives.scala 321:19:@38204.4]
  reg [31:0] _RAND_0;
  wire [22:0] _T_68; // @[MemPrimitives.scala 325:32:@38206.4]
  wire [22:0] _T_69; // @[MemPrimitives.scala 325:12:@38207.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@38206.4]
  assign _T_69 = io_wPort_0_reset ? 23'h0 : _T_68; // @[MemPrimitives.scala 325:12:@38207.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@38209.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[22:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 23'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 23'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_5( // @[:@38224.2]
  input         clock, // @[:@38225.4]
  input         reset, // @[:@38226.4]
  input         io_input_reset, // @[:@38227.4]
  input         io_input_enable, // @[:@38227.4]
  output [22:0] io_output_count_0, // @[:@38227.4]
  output        io_output_oobs_0, // @[:@38227.4]
  output        io_output_done // @[:@38227.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@38240.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@38240.4]
  wire [22:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@38240.4]
  wire [22:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@38240.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@38240.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@38240.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@38256.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@38256.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@38256.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@38256.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@38256.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@38256.4]
  wire  _T_36; // @[Counter.scala 264:45:@38259.4]
  wire [22:0] _T_48; // @[Counter.scala 287:52:@38284.4]
  wire [23:0] _T_50; // @[Counter.scala 291:33:@38285.4]
  wire [22:0] _T_51; // @[Counter.scala 291:33:@38286.4]
  wire [22:0] _T_52; // @[Counter.scala 291:33:@38287.4]
  wire  _T_57; // @[Counter.scala 293:18:@38289.4]
  wire [22:0] _T_68; // @[Counter.scala 299:115:@38297.4]
  wire [22:0] _T_71; // @[Counter.scala 299:152:@38300.4]
  wire [22:0] _T_72; // @[Counter.scala 299:74:@38301.4]
  wire  _T_75; // @[Counter.scala 322:102:@38305.4]
  wire  _T_77; // @[Counter.scala 322:130:@38306.4]
  FF_13 bases_0 ( // @[Counter.scala 261:53:@38240.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@38256.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@38259.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@38284.4]
  assign _T_50 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@38285.4]
  assign _T_51 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@38286.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@38287.4]
  assign _T_57 = $signed(_T_52) >= $signed(23'sh1fa400); // @[Counter.scala 293:18:@38289.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@38297.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@38300.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@38301.4]
  assign _T_75 = $signed(_T_48) < $signed(23'sh0); // @[Counter.scala 322:102:@38305.4]
  assign _T_77 = $signed(_T_48) >= $signed(23'sh1fa400); // @[Counter.scala 322:130:@38306.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@38304.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@38308.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@38310.4]
  assign bases_0_clock = clock; // @[:@38241.4]
  assign bases_0_reset = reset; // @[:@38242.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 23'h0 : _T_72; // @[Counter.scala 299:31:@38303.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@38282.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@38283.4]
  assign SRFF_clock = clock; // @[:@38257.4]
  assign SRFF_reset = reset; // @[:@38258.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@38261.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@38263.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@38264.4]
endmodule
module x477_ctrchain( // @[:@38315.2]
  input         clock, // @[:@38316.4]
  input         reset, // @[:@38317.4]
  input         io_input_reset, // @[:@38318.4]
  input         io_input_enable, // @[:@38318.4]
  output [22:0] io_output_counts_0, // @[:@38318.4]
  output        io_output_oobs_0, // @[:@38318.4]
  output        io_output_done // @[:@38318.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@38320.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@38320.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@38320.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@38320.4]
  wire [22:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@38320.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@38320.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@38320.4]
  reg  wasDone; // @[Counter.scala 542:24:@38329.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 546:69:@38335.4]
  wire  _T_47; // @[Counter.scala 546:80:@38336.4]
  reg  doneLatch; // @[Counter.scala 550:26:@38341.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 551:48:@38342.4]
  wire  _T_55; // @[Counter.scala 551:19:@38343.4]
  SingleCounter_5 ctrs_0 ( // @[Counter.scala 513:46:@38320.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 546:69:@38335.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 546:80:@38336.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@38342.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 551:19:@38343.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@38345.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@38347.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 546:18:@38338.4]
  assign ctrs_0_clock = clock; // @[:@38321.4]
  assign ctrs_0_reset = reset; // @[:@38322.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@38326.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@38327.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x484_inr_Foreach_sm( // @[:@38535.2]
  input   clock, // @[:@38536.4]
  input   reset, // @[:@38537.4]
  input   io_enable, // @[:@38538.4]
  output  io_done, // @[:@38538.4]
  output  io_doneLatch, // @[:@38538.4]
  input   io_ctrDone, // @[:@38538.4]
  output  io_datapathEn, // @[:@38538.4]
  output  io_ctrInc, // @[:@38538.4]
  output  io_ctrRst, // @[:@38538.4]
  input   io_parentAck, // @[:@38538.4]
  input   io_backpressure, // @[:@38538.4]
  input   io_break // @[:@38538.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@38540.4]
  wire  active_reset; // @[Controllers.scala 261:22:@38540.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@38540.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@38540.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@38540.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@38540.4]
  wire  done_clock; // @[Controllers.scala 262:20:@38543.4]
  wire  done_reset; // @[Controllers.scala 262:20:@38543.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@38543.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@38543.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@38543.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@38543.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@38577.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@38577.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@38577.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@38577.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@38577.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@38599.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@38599.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@38599.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@38599.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@38599.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@38611.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@38611.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@38611.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@38611.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@38611.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@38619.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@38619.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@38619.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@38619.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@38619.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@38635.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@38635.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@38635.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@38635.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@38635.4]
  wire  _T_80; // @[Controllers.scala 264:48:@38548.4]
  wire  _T_81; // @[Controllers.scala 264:46:@38549.4]
  wire  _T_82; // @[Controllers.scala 264:62:@38550.4]
  wire  _T_83; // @[Controllers.scala 264:60:@38551.4]
  wire  _T_100; // @[package.scala 100:49:@38568.4]
  reg  _T_103; // @[package.scala 48:56:@38569.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@38582.4 package.scala 96:25:@38583.4]
  wire  _T_110; // @[package.scala 100:49:@38584.4]
  reg  _T_113; // @[package.scala 48:56:@38585.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@38587.4]
  wire  _T_118; // @[Controllers.scala 283:41:@38592.4]
  wire  _T_119; // @[Controllers.scala 283:59:@38593.4]
  wire  _T_121; // @[Controllers.scala 284:37:@38596.4]
  wire  _T_124; // @[package.scala 96:25:@38604.4 package.scala 96:25:@38605.4]
  wire  _T_126; // @[package.scala 100:49:@38606.4]
  reg  _T_129; // @[package.scala 48:56:@38607.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@38629.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@38631.4]
  reg  _T_153; // @[package.scala 48:56:@38632.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@38640.4 package.scala 96:25:@38641.4]
  wire  _T_158; // @[Controllers.scala 292:61:@38642.4]
  wire  _T_159; // @[Controllers.scala 292:24:@38643.4]
  SRFF active ( // @[Controllers.scala 261:22:@38540.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@38543.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@38577.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@38599.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@38611.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@38619.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@38635.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@38548.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@38549.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@38550.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@38551.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@38568.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@38582.4 package.scala 96:25:@38583.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@38584.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@38587.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@38592.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@38593.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@38596.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@38604.4 package.scala 96:25:@38605.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@38606.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@38631.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@38640.4 package.scala 96:25:@38641.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@38642.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@38643.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@38610.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@38645.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@38595.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@38598.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@38590.4]
  assign active_clock = clock; // @[:@38541.4]
  assign active_reset = reset; // @[:@38542.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@38553.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@38557.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@38558.4]
  assign done_clock = clock; // @[:@38544.4]
  assign done_reset = reset; // @[:@38545.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@38573.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@38566.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@38567.4]
  assign RetimeWrapper_clock = clock; // @[:@38578.4]
  assign RetimeWrapper_reset = reset; // @[:@38579.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@38581.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@38580.4]
  assign RetimeWrapper_1_clock = clock; // @[:@38600.4]
  assign RetimeWrapper_1_reset = reset; // @[:@38601.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@38603.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@38602.4]
  assign RetimeWrapper_2_clock = clock; // @[:@38612.4]
  assign RetimeWrapper_2_reset = reset; // @[:@38613.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@38615.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@38614.4]
  assign RetimeWrapper_3_clock = clock; // @[:@38620.4]
  assign RetimeWrapper_3_reset = reset; // @[:@38621.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@38623.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@38622.4]
  assign RetimeWrapper_4_clock = clock; // @[:@38636.4]
  assign RetimeWrapper_4_reset = reset; // @[:@38637.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@38639.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@38638.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x484_inr_Foreach_kernelx484_inr_Foreach_concrete1( // @[:@38852.2]
  input         clock, // @[:@38853.4]
  input         reset, // @[:@38854.4]
  output [20:0] io_in_x252_outbuf_0_rPort_0_ofs_0, // @[:@38855.4]
  output        io_in_x252_outbuf_0_rPort_0_en_0, // @[:@38855.4]
  output        io_in_x252_outbuf_0_rPort_0_backpressure, // @[:@38855.4]
  input  [31:0] io_in_x252_outbuf_0_rPort_0_output_0, // @[:@38855.4]
  output        io_in_x469_valid, // @[:@38855.4]
  output [31:0] io_in_x469_bits_wdata_0, // @[:@38855.4]
  output        io_in_x469_bits_wstrb, // @[:@38855.4]
  input         io_sigsIn_backpressure, // @[:@38855.4]
  input         io_sigsIn_datapathEn, // @[:@38855.4]
  input         io_sigsIn_break, // @[:@38855.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@38855.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@38855.4]
  input         io_rr // @[:@38855.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@38882.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@38882.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@38911.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@38911.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@38911.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@38911.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@38911.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@38920.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@38920.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@38920.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@38920.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@38920.4]
  wire  b479; // @[sm_x484_inr_Foreach.scala 62:18:@38890.4]
  wire  _T_274; // @[sm_x484_inr_Foreach.scala 67:129:@38894.4]
  wire  _T_278; // @[implicits.scala 55:10:@38897.4]
  wire  _T_279; // @[sm_x484_inr_Foreach.scala 67:146:@38898.4]
  wire [32:0] x482_tuple; // @[Cat.scala 30:58:@38908.4]
  wire  _T_290; // @[package.scala 96:25:@38925.4 package.scala 96:25:@38926.4]
  wire  _T_292; // @[implicits.scala 55:10:@38927.4]
  wire  x621_b479_D2; // @[package.scala 96:25:@38916.4 package.scala 96:25:@38917.4]
  wire  _T_293; // @[sm_x484_inr_Foreach.scala 74:112:@38928.4]
  wire [31:0] b478_number; // @[Math.scala 723:22:@38887.4 Math.scala 724:14:@38888.4]
  _ _ ( // @[Math.scala 720:24:@38882.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@38911.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@38920.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign b479 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x484_inr_Foreach.scala 62:18:@38890.4]
  assign _T_274 = ~ io_sigsIn_break; // @[sm_x484_inr_Foreach.scala 67:129:@38894.4]
  assign _T_278 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@38897.4]
  assign _T_279 = _T_274 & _T_278; // @[sm_x484_inr_Foreach.scala 67:146:@38898.4]
  assign x482_tuple = {1'h1,io_in_x252_outbuf_0_rPort_0_output_0}; // @[Cat.scala 30:58:@38908.4]
  assign _T_290 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@38925.4 package.scala 96:25:@38926.4]
  assign _T_292 = io_rr ? _T_290 : 1'h0; // @[implicits.scala 55:10:@38927.4]
  assign x621_b479_D2 = RetimeWrapper_io_out; // @[package.scala 96:25:@38916.4 package.scala 96:25:@38917.4]
  assign _T_293 = _T_292 & x621_b479_D2; // @[sm_x484_inr_Foreach.scala 74:112:@38928.4]
  assign b478_number = __io_result; // @[Math.scala 723:22:@38887.4 Math.scala 724:14:@38888.4]
  assign io_in_x252_outbuf_0_rPort_0_ofs_0 = b478_number[20:0]; // @[MemInterfaceType.scala 107:54:@38901.4]
  assign io_in_x252_outbuf_0_rPort_0_en_0 = _T_279 & b479; // @[MemInterfaceType.scala 110:79:@38903.4]
  assign io_in_x252_outbuf_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@38902.4]
  assign io_in_x469_valid = _T_293 & io_sigsIn_backpressure; // @[sm_x484_inr_Foreach.scala 74:18:@38930.4]
  assign io_in_x469_bits_wdata_0 = x482_tuple[31:0]; // @[sm_x484_inr_Foreach.scala 75:26:@38932.4]
  assign io_in_x469_bits_wstrb = x482_tuple[32]; // @[sm_x484_inr_Foreach.scala 76:23:@38934.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@38885.4]
  assign RetimeWrapper_clock = clock; // @[:@38912.4]
  assign RetimeWrapper_reset = reset; // @[:@38913.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38915.4]
  assign RetimeWrapper_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@38914.4]
  assign RetimeWrapper_1_clock = clock; // @[:@38921.4]
  assign RetimeWrapper_1_reset = reset; // @[:@38922.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@38924.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@38923.4]
endmodule
module x488_inr_UnitPipe_sm( // @[:@39090.2]
  input   clock, // @[:@39091.4]
  input   reset, // @[:@39092.4]
  input   io_enable, // @[:@39093.4]
  output  io_done, // @[:@39093.4]
  output  io_doneLatch, // @[:@39093.4]
  input   io_ctrDone, // @[:@39093.4]
  output  io_datapathEn, // @[:@39093.4]
  output  io_ctrInc, // @[:@39093.4]
  input   io_parentAck // @[:@39093.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@39095.4]
  wire  active_reset; // @[Controllers.scala 261:22:@39095.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@39095.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@39095.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@39095.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@39095.4]
  wire  done_clock; // @[Controllers.scala 262:20:@39098.4]
  wire  done_reset; // @[Controllers.scala 262:20:@39098.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@39098.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@39098.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@39098.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@39098.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@39132.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@39132.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@39132.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@39132.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@39132.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@39154.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@39154.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@39154.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@39154.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@39154.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@39166.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@39166.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@39166.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@39166.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@39166.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@39174.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@39174.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@39174.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@39174.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@39174.4]
  wire  _T_80; // @[Controllers.scala 264:48:@39103.4]
  wire  _T_81; // @[Controllers.scala 264:46:@39104.4]
  wire  _T_82; // @[Controllers.scala 264:62:@39105.4]
  wire  _T_100; // @[package.scala 100:49:@39123.4]
  reg  _T_103; // @[package.scala 48:56:@39124.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@39147.4]
  wire  _T_124; // @[package.scala 96:25:@39159.4 package.scala 96:25:@39160.4]
  wire  _T_126; // @[package.scala 100:49:@39161.4]
  reg  _T_129; // @[package.scala 48:56:@39162.4]
  reg [31:0] _RAND_1;
  reg  _T_146; // @[Controllers.scala 291:31:@39184.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@39186.4]
  reg  _T_153; // @[package.scala 48:56:@39187.4]
  reg [31:0] _RAND_3;
  wire  _T_154; // @[package.scala 100:41:@39189.4]
  wire  _T_156; // @[Controllers.scala 292:61:@39190.4]
  wire  _T_157; // @[Controllers.scala 292:24:@39191.4]
  SRFF active ( // @[Controllers.scala 261:22:@39095.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@39098.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@39132.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@39154.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@39166.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@39174.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@39103.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@39104.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@39105.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@39123.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@39147.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@39159.4 package.scala 96:25:@39160.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@39161.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@39186.4]
  assign _T_154 = done_io_output & _T_153; // @[package.scala 100:41:@39189.4]
  assign _T_156 = _T_154 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@39190.4]
  assign _T_157 = io_parentAck ? 1'h0 : _T_156; // @[Controllers.scala 292:24:@39191.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@39165.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@39193.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@39150.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@39153.4]
  assign active_clock = clock; // @[:@39096.4]
  assign active_reset = reset; // @[:@39097.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@39108.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@39112.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@39113.4]
  assign done_clock = clock; // @[:@39099.4]
  assign done_reset = reset; // @[:@39100.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@39128.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@39121.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@39122.4]
  assign RetimeWrapper_clock = clock; // @[:@39133.4]
  assign RetimeWrapper_reset = reset; // @[:@39134.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@39136.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@39135.4]
  assign RetimeWrapper_1_clock = clock; // @[:@39155.4]
  assign RetimeWrapper_1_reset = reset; // @[:@39156.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@39158.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@39157.4]
  assign RetimeWrapper_2_clock = clock; // @[:@39167.4]
  assign RetimeWrapper_2_reset = reset; // @[:@39168.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@39170.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@39169.4]
  assign RetimeWrapper_3_clock = clock; // @[:@39175.4]
  assign RetimeWrapper_3_reset = reset; // @[:@39176.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@39178.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@39177.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_154) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x488_inr_UnitPipe_kernelx488_inr_UnitPipe_concrete1( // @[:@39268.2]
  output  io_in_x470_ready, // @[:@39271.4]
  input   io_sigsIn_datapathEn // @[:@39271.4]
);
  assign io_in_x470_ready = io_sigsIn_datapathEn; // @[sm_x488_inr_UnitPipe.scala 57:18:@39283.4]
endmodule
module x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1( // @[:@39286.2]
  input         clock, // @[:@39287.4]
  input         reset, // @[:@39288.4]
  input         io_in_x468_ready, // @[:@39289.4]
  output        io_in_x468_valid, // @[:@39289.4]
  output [63:0] io_in_x468_bits_addr, // @[:@39289.4]
  output [31:0] io_in_x468_bits_size, // @[:@39289.4]
  input  [63:0] io_in_x248_outdram_number, // @[:@39289.4]
  output [20:0] io_in_x252_outbuf_0_rPort_0_ofs_0, // @[:@39289.4]
  output        io_in_x252_outbuf_0_rPort_0_en_0, // @[:@39289.4]
  output        io_in_x252_outbuf_0_rPort_0_backpressure, // @[:@39289.4]
  input  [31:0] io_in_x252_outbuf_0_rPort_0_output_0, // @[:@39289.4]
  output        io_in_x470_ready, // @[:@39289.4]
  input         io_in_x470_valid, // @[:@39289.4]
  input         io_in_x469_ready, // @[:@39289.4]
  output        io_in_x469_valid, // @[:@39289.4]
  output [31:0] io_in_x469_bits_wdata_0, // @[:@39289.4]
  output        io_in_x469_bits_wstrb, // @[:@39289.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@39289.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@39289.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@39289.4]
  input         io_sigsIn_smChildAcks_0, // @[:@39289.4]
  input         io_sigsIn_smChildAcks_1, // @[:@39289.4]
  input         io_sigsIn_smChildAcks_2, // @[:@39289.4]
  output        io_sigsOut_smDoneIn_0, // @[:@39289.4]
  output        io_sigsOut_smDoneIn_1, // @[:@39289.4]
  output        io_sigsOut_smDoneIn_2, // @[:@39289.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@39289.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@39289.4]
  output        io_sigsOut_smCtrCopyDone_2, // @[:@39289.4]
  input         io_rr // @[:@39289.4]
);
  wire  x475_inr_UnitPipe_sm_clock; // @[sm_x475_inr_UnitPipe.scala 33:18:@39356.4]
  wire  x475_inr_UnitPipe_sm_reset; // @[sm_x475_inr_UnitPipe.scala 33:18:@39356.4]
  wire  x475_inr_UnitPipe_sm_io_enable; // @[sm_x475_inr_UnitPipe.scala 33:18:@39356.4]
  wire  x475_inr_UnitPipe_sm_io_done; // @[sm_x475_inr_UnitPipe.scala 33:18:@39356.4]
  wire  x475_inr_UnitPipe_sm_io_doneLatch; // @[sm_x475_inr_UnitPipe.scala 33:18:@39356.4]
  wire  x475_inr_UnitPipe_sm_io_ctrDone; // @[sm_x475_inr_UnitPipe.scala 33:18:@39356.4]
  wire  x475_inr_UnitPipe_sm_io_datapathEn; // @[sm_x475_inr_UnitPipe.scala 33:18:@39356.4]
  wire  x475_inr_UnitPipe_sm_io_ctrInc; // @[sm_x475_inr_UnitPipe.scala 33:18:@39356.4]
  wire  x475_inr_UnitPipe_sm_io_parentAck; // @[sm_x475_inr_UnitPipe.scala 33:18:@39356.4]
  wire  x475_inr_UnitPipe_sm_io_backpressure; // @[sm_x475_inr_UnitPipe.scala 33:18:@39356.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@39413.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@39413.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@39413.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@39413.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@39413.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@39421.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@39421.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@39421.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@39421.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@39421.4]
  wire  x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_in_x468_valid; // @[sm_x475_inr_UnitPipe.scala 69:24:@39451.4]
  wire [63:0] x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_in_x468_bits_addr; // @[sm_x475_inr_UnitPipe.scala 69:24:@39451.4]
  wire [31:0] x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_in_x468_bits_size; // @[sm_x475_inr_UnitPipe.scala 69:24:@39451.4]
  wire [63:0] x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_in_x248_outdram_number; // @[sm_x475_inr_UnitPipe.scala 69:24:@39451.4]
  wire  x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x475_inr_UnitPipe.scala 69:24:@39451.4]
  wire  x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x475_inr_UnitPipe.scala 69:24:@39451.4]
  wire  x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_rr; // @[sm_x475_inr_UnitPipe.scala 69:24:@39451.4]
  wire  x477_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@39519.4]
  wire  x477_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@39519.4]
  wire  x477_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@39519.4]
  wire  x477_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@39519.4]
  wire [22:0] x477_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@39519.4]
  wire  x477_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@39519.4]
  wire  x477_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@39519.4]
  wire  x484_inr_Foreach_sm_clock; // @[sm_x484_inr_Foreach.scala 33:18:@39572.4]
  wire  x484_inr_Foreach_sm_reset; // @[sm_x484_inr_Foreach.scala 33:18:@39572.4]
  wire  x484_inr_Foreach_sm_io_enable; // @[sm_x484_inr_Foreach.scala 33:18:@39572.4]
  wire  x484_inr_Foreach_sm_io_done; // @[sm_x484_inr_Foreach.scala 33:18:@39572.4]
  wire  x484_inr_Foreach_sm_io_doneLatch; // @[sm_x484_inr_Foreach.scala 33:18:@39572.4]
  wire  x484_inr_Foreach_sm_io_ctrDone; // @[sm_x484_inr_Foreach.scala 33:18:@39572.4]
  wire  x484_inr_Foreach_sm_io_datapathEn; // @[sm_x484_inr_Foreach.scala 33:18:@39572.4]
  wire  x484_inr_Foreach_sm_io_ctrInc; // @[sm_x484_inr_Foreach.scala 33:18:@39572.4]
  wire  x484_inr_Foreach_sm_io_ctrRst; // @[sm_x484_inr_Foreach.scala 33:18:@39572.4]
  wire  x484_inr_Foreach_sm_io_parentAck; // @[sm_x484_inr_Foreach.scala 33:18:@39572.4]
  wire  x484_inr_Foreach_sm_io_backpressure; // @[sm_x484_inr_Foreach.scala 33:18:@39572.4]
  wire  x484_inr_Foreach_sm_io_break; // @[sm_x484_inr_Foreach.scala 33:18:@39572.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@39600.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@39600.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@39600.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@39600.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@39600.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@39640.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@39640.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@39640.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@39640.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@39640.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@39648.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@39648.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@39648.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@39648.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@39648.4]
  wire  x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_clock; // @[sm_x484_inr_Foreach.scala 78:24:@39683.4]
  wire  x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_reset; // @[sm_x484_inr_Foreach.scala 78:24:@39683.4]
  wire [20:0] x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x252_outbuf_0_rPort_0_ofs_0; // @[sm_x484_inr_Foreach.scala 78:24:@39683.4]
  wire  x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x252_outbuf_0_rPort_0_en_0; // @[sm_x484_inr_Foreach.scala 78:24:@39683.4]
  wire  x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x252_outbuf_0_rPort_0_backpressure; // @[sm_x484_inr_Foreach.scala 78:24:@39683.4]
  wire [31:0] x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x252_outbuf_0_rPort_0_output_0; // @[sm_x484_inr_Foreach.scala 78:24:@39683.4]
  wire  x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x469_valid; // @[sm_x484_inr_Foreach.scala 78:24:@39683.4]
  wire [31:0] x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x469_bits_wdata_0; // @[sm_x484_inr_Foreach.scala 78:24:@39683.4]
  wire  x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x469_bits_wstrb; // @[sm_x484_inr_Foreach.scala 78:24:@39683.4]
  wire  x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x484_inr_Foreach.scala 78:24:@39683.4]
  wire  x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x484_inr_Foreach.scala 78:24:@39683.4]
  wire  x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x484_inr_Foreach.scala 78:24:@39683.4]
  wire [31:0] x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x484_inr_Foreach.scala 78:24:@39683.4]
  wire  x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x484_inr_Foreach.scala 78:24:@39683.4]
  wire  x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_rr; // @[sm_x484_inr_Foreach.scala 78:24:@39683.4]
  wire  x488_inr_UnitPipe_sm_clock; // @[sm_x488_inr_UnitPipe.scala 32:18:@39803.4]
  wire  x488_inr_UnitPipe_sm_reset; // @[sm_x488_inr_UnitPipe.scala 32:18:@39803.4]
  wire  x488_inr_UnitPipe_sm_io_enable; // @[sm_x488_inr_UnitPipe.scala 32:18:@39803.4]
  wire  x488_inr_UnitPipe_sm_io_done; // @[sm_x488_inr_UnitPipe.scala 32:18:@39803.4]
  wire  x488_inr_UnitPipe_sm_io_doneLatch; // @[sm_x488_inr_UnitPipe.scala 32:18:@39803.4]
  wire  x488_inr_UnitPipe_sm_io_ctrDone; // @[sm_x488_inr_UnitPipe.scala 32:18:@39803.4]
  wire  x488_inr_UnitPipe_sm_io_datapathEn; // @[sm_x488_inr_UnitPipe.scala 32:18:@39803.4]
  wire  x488_inr_UnitPipe_sm_io_ctrInc; // @[sm_x488_inr_UnitPipe.scala 32:18:@39803.4]
  wire  x488_inr_UnitPipe_sm_io_parentAck; // @[sm_x488_inr_UnitPipe.scala 32:18:@39803.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@39860.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@39860.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@39860.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@39860.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@39860.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@39868.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@39868.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@39868.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@39868.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@39868.4]
  wire  x488_inr_UnitPipe_kernelx488_inr_UnitPipe_concrete1_io_in_x470_ready; // @[sm_x488_inr_UnitPipe.scala 60:24:@39898.4]
  wire  x488_inr_UnitPipe_kernelx488_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x488_inr_UnitPipe.scala 60:24:@39898.4]
  wire  _T_359; // @[package.scala 100:49:@39384.4]
  reg  _T_362; // @[package.scala 48:56:@39385.4]
  reg [31:0] _RAND_0;
  wire  _T_375; // @[package.scala 96:25:@39418.4 package.scala 96:25:@39419.4]
  wire  _T_381; // @[package.scala 96:25:@39426.4 package.scala 96:25:@39427.4]
  wire  _T_384; // @[SpatialBlocks.scala 138:93:@39429.4]
  wire  _T_454; // @[package.scala 96:25:@39605.4 package.scala 96:25:@39606.4]
  wire  _T_468; // @[package.scala 96:25:@39645.4 package.scala 96:25:@39646.4]
  wire  _T_474; // @[package.scala 96:25:@39653.4 package.scala 96:25:@39654.4]
  wire  _T_477; // @[SpatialBlocks.scala 138:93:@39656.4]
  wire  _T_479; // @[SpatialBlocks.scala 157:36:@39665.4]
  wire  _T_480; // @[SpatialBlocks.scala 157:78:@39666.4]
  wire  _T_547; // @[package.scala 100:49:@39831.4]
  reg  _T_550; // @[package.scala 48:56:@39832.4]
  reg [31:0] _RAND_1;
  wire  x488_inr_UnitPipe_sigsIn_forwardpressure; // @[sm_x489_outr_UnitPipe.scala 101:55:@39838.4]
  wire  _T_563; // @[package.scala 96:25:@39865.4 package.scala 96:25:@39866.4]
  wire  _T_569; // @[package.scala 96:25:@39873.4 package.scala 96:25:@39874.4]
  wire  _T_572; // @[SpatialBlocks.scala 138:93:@39876.4]
  wire  x488_inr_UnitPipe_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@39877.4]
  x475_inr_UnitPipe_sm x475_inr_UnitPipe_sm ( // @[sm_x475_inr_UnitPipe.scala 33:18:@39356.4]
    .clock(x475_inr_UnitPipe_sm_clock),
    .reset(x475_inr_UnitPipe_sm_reset),
    .io_enable(x475_inr_UnitPipe_sm_io_enable),
    .io_done(x475_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x475_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x475_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x475_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x475_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x475_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x475_inr_UnitPipe_sm_io_backpressure)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@39413.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@39421.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1 x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1 ( // @[sm_x475_inr_UnitPipe.scala 69:24:@39451.4]
    .io_in_x468_valid(x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_in_x468_valid),
    .io_in_x468_bits_addr(x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_in_x468_bits_addr),
    .io_in_x468_bits_size(x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_in_x468_bits_size),
    .io_in_x248_outdram_number(x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_in_x248_outdram_number),
    .io_sigsIn_backpressure(x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_rr(x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_rr)
  );
  x477_ctrchain x477_ctrchain ( // @[SpatialBlocks.scala 37:22:@39519.4]
    .clock(x477_ctrchain_clock),
    .reset(x477_ctrchain_reset),
    .io_input_reset(x477_ctrchain_io_input_reset),
    .io_input_enable(x477_ctrchain_io_input_enable),
    .io_output_counts_0(x477_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x477_ctrchain_io_output_oobs_0),
    .io_output_done(x477_ctrchain_io_output_done)
  );
  x484_inr_Foreach_sm x484_inr_Foreach_sm ( // @[sm_x484_inr_Foreach.scala 33:18:@39572.4]
    .clock(x484_inr_Foreach_sm_clock),
    .reset(x484_inr_Foreach_sm_reset),
    .io_enable(x484_inr_Foreach_sm_io_enable),
    .io_done(x484_inr_Foreach_sm_io_done),
    .io_doneLatch(x484_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x484_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x484_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x484_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x484_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x484_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x484_inr_Foreach_sm_io_backpressure),
    .io_break(x484_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@39600.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@39640.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@39648.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x484_inr_Foreach_kernelx484_inr_Foreach_concrete1 x484_inr_Foreach_kernelx484_inr_Foreach_concrete1 ( // @[sm_x484_inr_Foreach.scala 78:24:@39683.4]
    .clock(x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_clock),
    .reset(x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_reset),
    .io_in_x252_outbuf_0_rPort_0_ofs_0(x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x252_outbuf_0_rPort_0_ofs_0),
    .io_in_x252_outbuf_0_rPort_0_en_0(x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x252_outbuf_0_rPort_0_en_0),
    .io_in_x252_outbuf_0_rPort_0_backpressure(x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x252_outbuf_0_rPort_0_backpressure),
    .io_in_x252_outbuf_0_rPort_0_output_0(x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x252_outbuf_0_rPort_0_output_0),
    .io_in_x469_valid(x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x469_valid),
    .io_in_x469_bits_wdata_0(x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x469_bits_wdata_0),
    .io_in_x469_bits_wstrb(x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x469_bits_wstrb),
    .io_sigsIn_backpressure(x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_rr)
  );
  x488_inr_UnitPipe_sm x488_inr_UnitPipe_sm ( // @[sm_x488_inr_UnitPipe.scala 32:18:@39803.4]
    .clock(x488_inr_UnitPipe_sm_clock),
    .reset(x488_inr_UnitPipe_sm_reset),
    .io_enable(x488_inr_UnitPipe_sm_io_enable),
    .io_done(x488_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x488_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x488_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x488_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x488_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x488_inr_UnitPipe_sm_io_parentAck)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@39860.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@39868.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x488_inr_UnitPipe_kernelx488_inr_UnitPipe_concrete1 x488_inr_UnitPipe_kernelx488_inr_UnitPipe_concrete1 ( // @[sm_x488_inr_UnitPipe.scala 60:24:@39898.4]
    .io_in_x470_ready(x488_inr_UnitPipe_kernelx488_inr_UnitPipe_concrete1_io_in_x470_ready),
    .io_sigsIn_datapathEn(x488_inr_UnitPipe_kernelx488_inr_UnitPipe_concrete1_io_sigsIn_datapathEn)
  );
  assign _T_359 = x475_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@39384.4]
  assign _T_375 = RetimeWrapper_io_out; // @[package.scala 96:25:@39418.4 package.scala 96:25:@39419.4]
  assign _T_381 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@39426.4 package.scala 96:25:@39427.4]
  assign _T_384 = ~ _T_381; // @[SpatialBlocks.scala 138:93:@39429.4]
  assign _T_454 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@39605.4 package.scala 96:25:@39606.4]
  assign _T_468 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@39645.4 package.scala 96:25:@39646.4]
  assign _T_474 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@39653.4 package.scala 96:25:@39654.4]
  assign _T_477 = ~ _T_474; // @[SpatialBlocks.scala 138:93:@39656.4]
  assign _T_479 = x484_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@39665.4]
  assign _T_480 = ~ x484_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@39666.4]
  assign _T_547 = x488_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@39831.4]
  assign x488_inr_UnitPipe_sigsIn_forwardpressure = io_in_x470_valid | x488_inr_UnitPipe_sm_io_doneLatch; // @[sm_x489_outr_UnitPipe.scala 101:55:@39838.4]
  assign _T_563 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@39865.4 package.scala 96:25:@39866.4]
  assign _T_569 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@39873.4 package.scala 96:25:@39874.4]
  assign _T_572 = ~ _T_569; // @[SpatialBlocks.scala 138:93:@39876.4]
  assign x488_inr_UnitPipe_sigsIn_baseEn = _T_563 & _T_572; // @[SpatialBlocks.scala 138:90:@39877.4]
  assign io_in_x468_valid = x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_in_x468_valid; // @[sm_x475_inr_UnitPipe.scala 49:23:@39489.4]
  assign io_in_x468_bits_addr = x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_in_x468_bits_addr; // @[sm_x475_inr_UnitPipe.scala 49:23:@39488.4]
  assign io_in_x468_bits_size = x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_in_x468_bits_size; // @[sm_x475_inr_UnitPipe.scala 49:23:@39487.4]
  assign io_in_x252_outbuf_0_rPort_0_ofs_0 = x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x252_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@39734.4]
  assign io_in_x252_outbuf_0_rPort_0_en_0 = x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x252_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@39733.4]
  assign io_in_x252_outbuf_0_rPort_0_backpressure = x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x252_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@39732.4]
  assign io_in_x470_ready = x488_inr_UnitPipe_kernelx488_inr_UnitPipe_concrete1_io_in_x470_ready; // @[sm_x488_inr_UnitPipe.scala 46:23:@39934.4]
  assign io_in_x469_valid = x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x469_valid; // @[sm_x484_inr_Foreach.scala 50:23:@39738.4]
  assign io_in_x469_bits_wdata_0 = x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x469_bits_wdata_0; // @[sm_x484_inr_Foreach.scala 50:23:@39737.4]
  assign io_in_x469_bits_wstrb = x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x469_bits_wstrb; // @[sm_x484_inr_Foreach.scala 50:23:@39736.4]
  assign io_sigsOut_smDoneIn_0 = x475_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@39436.4]
  assign io_sigsOut_smDoneIn_1 = x484_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@39663.4]
  assign io_sigsOut_smDoneIn_2 = x488_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@39883.4]
  assign io_sigsOut_smCtrCopyDone_0 = x475_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@39450.4]
  assign io_sigsOut_smCtrCopyDone_1 = x484_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@39682.4]
  assign io_sigsOut_smCtrCopyDone_2 = x488_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@39897.4]
  assign x475_inr_UnitPipe_sm_clock = clock; // @[:@39357.4]
  assign x475_inr_UnitPipe_sm_reset = reset; // @[:@39358.4]
  assign x475_inr_UnitPipe_sm_io_enable = _T_375 & _T_384; // @[SpatialBlocks.scala 140:18:@39433.4]
  assign x475_inr_UnitPipe_sm_io_ctrDone = x475_inr_UnitPipe_sm_io_ctrInc & _T_362; // @[sm_x489_outr_UnitPipe.scala 77:39:@39388.4]
  assign x475_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@39435.4]
  assign x475_inr_UnitPipe_sm_io_backpressure = io_in_x468_ready | x475_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@39407.4]
  assign RetimeWrapper_clock = clock; // @[:@39414.4]
  assign RetimeWrapper_reset = reset; // @[:@39415.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@39417.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@39416.4]
  assign RetimeWrapper_1_clock = clock; // @[:@39422.4]
  assign RetimeWrapper_1_reset = reset; // @[:@39423.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@39425.4]
  assign RetimeWrapper_1_io_in = x475_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@39424.4]
  assign x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_in_x248_outdram_number = io_in_x248_outdram_number; // @[sm_x475_inr_UnitPipe.scala 50:31:@39491.4]
  assign x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x468_ready | x475_inr_UnitPipe_sm_io_doneLatch; // @[sm_x475_inr_UnitPipe.scala 74:22:@39506.4]
  assign x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x475_inr_UnitPipe_sm_io_datapathEn; // @[sm_x475_inr_UnitPipe.scala 74:22:@39504.4]
  assign x475_inr_UnitPipe_kernelx475_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x475_inr_UnitPipe.scala 73:18:@39492.4]
  assign x477_ctrchain_clock = clock; // @[:@39520.4]
  assign x477_ctrchain_reset = reset; // @[:@39521.4]
  assign x477_ctrchain_io_input_reset = x484_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@39681.4]
  assign x477_ctrchain_io_input_enable = x484_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@39633.4 SpatialBlocks.scala 159:42:@39680.4]
  assign x484_inr_Foreach_sm_clock = clock; // @[:@39573.4]
  assign x484_inr_Foreach_sm_reset = reset; // @[:@39574.4]
  assign x484_inr_Foreach_sm_io_enable = _T_468 & _T_477; // @[SpatialBlocks.scala 140:18:@39660.4]
  assign x484_inr_Foreach_sm_io_ctrDone = io_rr ? _T_454 : 1'h0; // @[sm_x489_outr_UnitPipe.scala 90:38:@39608.4]
  assign x484_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@39662.4]
  assign x484_inr_Foreach_sm_io_backpressure = io_in_x469_ready | x484_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@39634.4]
  assign x484_inr_Foreach_sm_io_break = 1'h0; // @[sm_x489_outr_UnitPipe.scala 94:36:@39614.4]
  assign RetimeWrapper_2_clock = clock; // @[:@39601.4]
  assign RetimeWrapper_2_reset = reset; // @[:@39602.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@39604.4]
  assign RetimeWrapper_2_io_in = x477_ctrchain_io_output_done; // @[package.scala 94:16:@39603.4]
  assign RetimeWrapper_3_clock = clock; // @[:@39641.4]
  assign RetimeWrapper_3_reset = reset; // @[:@39642.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@39644.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@39643.4]
  assign RetimeWrapper_4_clock = clock; // @[:@39649.4]
  assign RetimeWrapper_4_reset = reset; // @[:@39650.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@39652.4]
  assign RetimeWrapper_4_io_in = x484_inr_Foreach_sm_io_done; // @[package.scala 94:16:@39651.4]
  assign x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_clock = clock; // @[:@39684.4]
  assign x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_reset = reset; // @[:@39685.4]
  assign x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_in_x252_outbuf_0_rPort_0_output_0 = io_in_x252_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@39731.4]
  assign x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x469_ready | x484_inr_Foreach_sm_io_doneLatch; // @[sm_x484_inr_Foreach.scala 83:22:@39754.4]
  assign x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_479 & _T_480; // @[sm_x484_inr_Foreach.scala 83:22:@39752.4]
  assign x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_sigsIn_break = x484_inr_Foreach_sm_io_break; // @[sm_x484_inr_Foreach.scala 83:22:@39750.4]
  assign x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{9{x477_ctrchain_io_output_counts_0[22]}},x477_ctrchain_io_output_counts_0}; // @[sm_x484_inr_Foreach.scala 83:22:@39745.4]
  assign x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x477_ctrchain_io_output_oobs_0; // @[sm_x484_inr_Foreach.scala 83:22:@39744.4]
  assign x484_inr_Foreach_kernelx484_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x484_inr_Foreach.scala 82:18:@39740.4]
  assign x488_inr_UnitPipe_sm_clock = clock; // @[:@39804.4]
  assign x488_inr_UnitPipe_sm_reset = reset; // @[:@39805.4]
  assign x488_inr_UnitPipe_sm_io_enable = x488_inr_UnitPipe_sigsIn_baseEn & x488_inr_UnitPipe_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@39880.4]
  assign x488_inr_UnitPipe_sm_io_ctrDone = x488_inr_UnitPipe_sm_io_ctrInc & _T_550; // @[sm_x489_outr_UnitPipe.scala 99:39:@39835.4]
  assign x488_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 142:21:@39882.4]
  assign RetimeWrapper_5_clock = clock; // @[:@39861.4]
  assign RetimeWrapper_5_reset = reset; // @[:@39862.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@39864.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@39863.4]
  assign RetimeWrapper_6_clock = clock; // @[:@39869.4]
  assign RetimeWrapper_6_reset = reset; // @[:@39870.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@39872.4]
  assign RetimeWrapper_6_io_in = x488_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@39871.4]
  assign x488_inr_UnitPipe_kernelx488_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x488_inr_UnitPipe_sm_io_datapathEn; // @[sm_x488_inr_UnitPipe.scala 65:22:@39947.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_362 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_550 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_362 <= 1'h0;
    end else begin
      _T_362 <= _T_359;
    end
    if (reset) begin
      _T_550 <= 1'h0;
    end else begin
      _T_550 <= _T_547;
    end
  end
endmodule
module x538_kernelx538_concrete1( // @[:@39963.2]
  input          clock, // @[:@39964.4]
  input          reset, // @[:@39965.4]
  input          io_in_x468_ready, // @[:@39966.4]
  output         io_in_x468_valid, // @[:@39966.4]
  output [63:0]  io_in_x468_bits_addr, // @[:@39966.4]
  output [31:0]  io_in_x468_bits_size, // @[:@39966.4]
  input  [63:0]  io_in_x248_outdram_number, // @[:@39966.4]
  output [20:0]  io_in_x252_outbuf_0_rPort_0_ofs_0, // @[:@39966.4]
  output         io_in_x252_outbuf_0_rPort_0_en_0, // @[:@39966.4]
  output         io_in_x252_outbuf_0_rPort_0_backpressure, // @[:@39966.4]
  input  [31:0]  io_in_x252_outbuf_0_rPort_0_output_0, // @[:@39966.4]
  output         io_in_x251_TVALID, // @[:@39966.4]
  input          io_in_x251_TREADY, // @[:@39966.4]
  output [255:0] io_in_x251_TDATA, // @[:@39966.4]
  output         io_in_x470_ready, // @[:@39966.4]
  input          io_in_x470_valid, // @[:@39966.4]
  input          io_in_x250_TVALID, // @[:@39966.4]
  output         io_in_x250_TREADY, // @[:@39966.4]
  input  [255:0] io_in_x250_TDATA, // @[:@39966.4]
  input  [7:0]   io_in_x250_TID, // @[:@39966.4]
  input  [7:0]   io_in_x250_TDEST, // @[:@39966.4]
  input          io_in_x469_ready, // @[:@39966.4]
  output         io_in_x469_valid, // @[:@39966.4]
  output [31:0]  io_in_x469_bits_wdata_0, // @[:@39966.4]
  output         io_in_x469_bits_wstrb, // @[:@39966.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@39966.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@39966.4]
  input          io_sigsIn_smChildAcks_0, // @[:@39966.4]
  input          io_sigsIn_smChildAcks_1, // @[:@39966.4]
  output         io_sigsOut_smDoneIn_0, // @[:@39966.4]
  output         io_sigsOut_smDoneIn_1, // @[:@39966.4]
  input          io_rr // @[:@39966.4]
);
  wire  x467_outr_UnitPipe_sm_clock; // @[sm_x467_outr_UnitPipe.scala 32:18:@40039.4]
  wire  x467_outr_UnitPipe_sm_reset; // @[sm_x467_outr_UnitPipe.scala 32:18:@40039.4]
  wire  x467_outr_UnitPipe_sm_io_enable; // @[sm_x467_outr_UnitPipe.scala 32:18:@40039.4]
  wire  x467_outr_UnitPipe_sm_io_done; // @[sm_x467_outr_UnitPipe.scala 32:18:@40039.4]
  wire  x467_outr_UnitPipe_sm_io_parentAck; // @[sm_x467_outr_UnitPipe.scala 32:18:@40039.4]
  wire  x467_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x467_outr_UnitPipe.scala 32:18:@40039.4]
  wire  x467_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x467_outr_UnitPipe.scala 32:18:@40039.4]
  wire  x467_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x467_outr_UnitPipe.scala 32:18:@40039.4]
  wire  x467_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x467_outr_UnitPipe.scala 32:18:@40039.4]
  wire  x467_outr_UnitPipe_sm_io_childAck_0; // @[sm_x467_outr_UnitPipe.scala 32:18:@40039.4]
  wire  x467_outr_UnitPipe_sm_io_childAck_1; // @[sm_x467_outr_UnitPipe.scala 32:18:@40039.4]
  wire  x467_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x467_outr_UnitPipe.scala 32:18:@40039.4]
  wire  x467_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x467_outr_UnitPipe.scala 32:18:@40039.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@40101.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@40101.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@40101.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@40101.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@40101.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@40109.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@40109.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@40109.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@40109.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@40109.4]
  wire  x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_clock; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire  x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_reset; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire  x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x251_TVALID; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire  x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x251_TREADY; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire [255:0] x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x251_TDATA; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire  x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x250_TVALID; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire  x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x250_TREADY; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire [255:0] x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x250_TDATA; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire [7:0] x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x250_TID; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire [7:0] x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x250_TDEST; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire  x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire  x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire  x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire  x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire  x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire  x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire  x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire  x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire  x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_rr; // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
  wire  x489_outr_UnitPipe_sm_clock; // @[sm_x489_outr_UnitPipe.scala 36:18:@40318.4]
  wire  x489_outr_UnitPipe_sm_reset; // @[sm_x489_outr_UnitPipe.scala 36:18:@40318.4]
  wire  x489_outr_UnitPipe_sm_io_enable; // @[sm_x489_outr_UnitPipe.scala 36:18:@40318.4]
  wire  x489_outr_UnitPipe_sm_io_done; // @[sm_x489_outr_UnitPipe.scala 36:18:@40318.4]
  wire  x489_outr_UnitPipe_sm_io_parentAck; // @[sm_x489_outr_UnitPipe.scala 36:18:@40318.4]
  wire  x489_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x489_outr_UnitPipe.scala 36:18:@40318.4]
  wire  x489_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x489_outr_UnitPipe.scala 36:18:@40318.4]
  wire  x489_outr_UnitPipe_sm_io_doneIn_2; // @[sm_x489_outr_UnitPipe.scala 36:18:@40318.4]
  wire  x489_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x489_outr_UnitPipe.scala 36:18:@40318.4]
  wire  x489_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x489_outr_UnitPipe.scala 36:18:@40318.4]
  wire  x489_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x489_outr_UnitPipe.scala 36:18:@40318.4]
  wire  x489_outr_UnitPipe_sm_io_childAck_0; // @[sm_x489_outr_UnitPipe.scala 36:18:@40318.4]
  wire  x489_outr_UnitPipe_sm_io_childAck_1; // @[sm_x489_outr_UnitPipe.scala 36:18:@40318.4]
  wire  x489_outr_UnitPipe_sm_io_childAck_2; // @[sm_x489_outr_UnitPipe.scala 36:18:@40318.4]
  wire  x489_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x489_outr_UnitPipe.scala 36:18:@40318.4]
  wire  x489_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x489_outr_UnitPipe.scala 36:18:@40318.4]
  wire  x489_outr_UnitPipe_sm_io_ctrCopyDone_2; // @[sm_x489_outr_UnitPipe.scala 36:18:@40318.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@40390.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@40390.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@40390.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@40390.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@40390.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@40398.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@40398.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@40398.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@40398.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@40398.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_clock; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_reset; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x468_ready; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x468_valid; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire [63:0] x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x468_bits_addr; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire [31:0] x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x468_bits_size; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire [63:0] x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x248_outdram_number; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire [20:0] x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x252_outbuf_0_rPort_0_ofs_0; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x252_outbuf_0_rPort_0_en_0; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x252_outbuf_0_rPort_0_backpressure; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire [31:0] x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x252_outbuf_0_rPort_0_output_0; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x470_ready; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x470_valid; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x469_ready; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x469_valid; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire [31:0] x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x469_bits_wdata_0; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x469_bits_wstrb; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_rr; // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
  wire  _T_408; // @[package.scala 96:25:@40106.4 package.scala 96:25:@40107.4]
  wire  _T_414; // @[package.scala 96:25:@40114.4 package.scala 96:25:@40115.4]
  wire  _T_417; // @[SpatialBlocks.scala 138:93:@40117.4]
  wire  _T_508; // @[package.scala 96:25:@40395.4 package.scala 96:25:@40396.4]
  wire  _T_514; // @[package.scala 96:25:@40403.4 package.scala 96:25:@40404.4]
  wire  _T_517; // @[SpatialBlocks.scala 138:93:@40406.4]
  x467_outr_UnitPipe_sm x467_outr_UnitPipe_sm ( // @[sm_x467_outr_UnitPipe.scala 32:18:@40039.4]
    .clock(x467_outr_UnitPipe_sm_clock),
    .reset(x467_outr_UnitPipe_sm_reset),
    .io_enable(x467_outr_UnitPipe_sm_io_enable),
    .io_done(x467_outr_UnitPipe_sm_io_done),
    .io_parentAck(x467_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x467_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x467_outr_UnitPipe_sm_io_doneIn_1),
    .io_enableOut_0(x467_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x467_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x467_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x467_outr_UnitPipe_sm_io_childAck_1),
    .io_ctrCopyDone_0(x467_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x467_outr_UnitPipe_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@40101.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@40109.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1 x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1 ( // @[sm_x467_outr_UnitPipe.scala 87:24:@40140.4]
    .clock(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_clock),
    .reset(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_reset),
    .io_in_x251_TVALID(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x251_TVALID),
    .io_in_x251_TREADY(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x251_TREADY),
    .io_in_x251_TDATA(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x251_TDATA),
    .io_in_x250_TVALID(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x250_TVALID),
    .io_in_x250_TREADY(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x250_TREADY),
    .io_in_x250_TDATA(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x250_TDATA),
    .io_in_x250_TID(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x250_TID),
    .io_in_x250_TDEST(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x250_TDEST),
    .io_sigsIn_smEnableOuts_0(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_rr)
  );
  x489_outr_UnitPipe_sm x489_outr_UnitPipe_sm ( // @[sm_x489_outr_UnitPipe.scala 36:18:@40318.4]
    .clock(x489_outr_UnitPipe_sm_clock),
    .reset(x489_outr_UnitPipe_sm_reset),
    .io_enable(x489_outr_UnitPipe_sm_io_enable),
    .io_done(x489_outr_UnitPipe_sm_io_done),
    .io_parentAck(x489_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x489_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x489_outr_UnitPipe_sm_io_doneIn_1),
    .io_doneIn_2(x489_outr_UnitPipe_sm_io_doneIn_2),
    .io_enableOut_0(x489_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x489_outr_UnitPipe_sm_io_enableOut_1),
    .io_enableOut_2(x489_outr_UnitPipe_sm_io_enableOut_2),
    .io_childAck_0(x489_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x489_outr_UnitPipe_sm_io_childAck_1),
    .io_childAck_2(x489_outr_UnitPipe_sm_io_childAck_2),
    .io_ctrCopyDone_0(x489_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x489_outr_UnitPipe_sm_io_ctrCopyDone_1),
    .io_ctrCopyDone_2(x489_outr_UnitPipe_sm_io_ctrCopyDone_2)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@40390.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@40398.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1 x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1 ( // @[sm_x489_outr_UnitPipe.scala 108:24:@40430.4]
    .clock(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_clock),
    .reset(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_reset),
    .io_in_x468_ready(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x468_ready),
    .io_in_x468_valid(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x468_valid),
    .io_in_x468_bits_addr(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x468_bits_addr),
    .io_in_x468_bits_size(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x468_bits_size),
    .io_in_x248_outdram_number(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x248_outdram_number),
    .io_in_x252_outbuf_0_rPort_0_ofs_0(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x252_outbuf_0_rPort_0_ofs_0),
    .io_in_x252_outbuf_0_rPort_0_en_0(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x252_outbuf_0_rPort_0_en_0),
    .io_in_x252_outbuf_0_rPort_0_backpressure(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x252_outbuf_0_rPort_0_backpressure),
    .io_in_x252_outbuf_0_rPort_0_output_0(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x252_outbuf_0_rPort_0_output_0),
    .io_in_x470_ready(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x470_ready),
    .io_in_x470_valid(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x470_valid),
    .io_in_x469_ready(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x469_ready),
    .io_in_x469_valid(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x469_valid),
    .io_in_x469_bits_wdata_0(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x469_bits_wdata_0),
    .io_in_x469_bits_wstrb(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x469_bits_wstrb),
    .io_sigsIn_smEnableOuts_0(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smCtrCopyDone_0(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_sigsOut_smCtrCopyDone_2(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2),
    .io_rr(x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_408 = RetimeWrapper_io_out; // @[package.scala 96:25:@40106.4 package.scala 96:25:@40107.4]
  assign _T_414 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@40114.4 package.scala 96:25:@40115.4]
  assign _T_417 = ~ _T_414; // @[SpatialBlocks.scala 138:93:@40117.4]
  assign _T_508 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@40395.4 package.scala 96:25:@40396.4]
  assign _T_514 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@40403.4 package.scala 96:25:@40404.4]
  assign _T_517 = ~ _T_514; // @[SpatialBlocks.scala 138:93:@40406.4]
  assign io_in_x468_valid = x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x468_valid; // @[sm_x489_outr_UnitPipe.scala 58:23:@40512.4]
  assign io_in_x468_bits_addr = x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x468_bits_addr; // @[sm_x489_outr_UnitPipe.scala 58:23:@40511.4]
  assign io_in_x468_bits_size = x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x468_bits_size; // @[sm_x489_outr_UnitPipe.scala 58:23:@40510.4]
  assign io_in_x252_outbuf_0_rPort_0_ofs_0 = x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x252_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@40518.4]
  assign io_in_x252_outbuf_0_rPort_0_en_0 = x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x252_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@40517.4]
  assign io_in_x252_outbuf_0_rPort_0_backpressure = x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x252_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@40516.4]
  assign io_in_x251_TVALID = x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x251_TVALID; // @[sm_x467_outr_UnitPipe.scala 48:23:@40209.4]
  assign io_in_x251_TDATA = x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x251_TDATA; // @[sm_x467_outr_UnitPipe.scala 48:23:@40207.4]
  assign io_in_x470_ready = x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x470_ready; // @[sm_x489_outr_UnitPipe.scala 61:23:@40522.4]
  assign io_in_x250_TREADY = x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x250_TREADY; // @[sm_x467_outr_UnitPipe.scala 49:23:@40217.4]
  assign io_in_x469_valid = x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x469_valid; // @[sm_x489_outr_UnitPipe.scala 62:23:@40525.4]
  assign io_in_x469_bits_wdata_0 = x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x469_bits_wdata_0; // @[sm_x489_outr_UnitPipe.scala 62:23:@40524.4]
  assign io_in_x469_bits_wstrb = x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x469_bits_wstrb; // @[sm_x489_outr_UnitPipe.scala 62:23:@40523.4]
  assign io_sigsOut_smDoneIn_0 = x467_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@40124.4]
  assign io_sigsOut_smDoneIn_1 = x489_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@40413.4]
  assign x467_outr_UnitPipe_sm_clock = clock; // @[:@40040.4]
  assign x467_outr_UnitPipe_sm_reset = reset; // @[:@40041.4]
  assign x467_outr_UnitPipe_sm_io_enable = _T_408 & _T_417; // @[SpatialBlocks.scala 140:18:@40121.4]
  assign x467_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@40123.4]
  assign x467_outr_UnitPipe_sm_io_doneIn_0 = x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@40091.4]
  assign x467_outr_UnitPipe_sm_io_doneIn_1 = x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@40092.4]
  assign x467_outr_UnitPipe_sm_io_ctrCopyDone_0 = x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@40138.4]
  assign x467_outr_UnitPipe_sm_io_ctrCopyDone_1 = x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@40139.4]
  assign RetimeWrapper_clock = clock; // @[:@40102.4]
  assign RetimeWrapper_reset = reset; // @[:@40103.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@40105.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@40104.4]
  assign RetimeWrapper_1_clock = clock; // @[:@40110.4]
  assign RetimeWrapper_1_reset = reset; // @[:@40111.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@40113.4]
  assign RetimeWrapper_1_io_in = x467_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@40112.4]
  assign x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_clock = clock; // @[:@40141.4]
  assign x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_reset = reset; // @[:@40142.4]
  assign x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x251_TREADY = io_in_x251_TREADY; // @[sm_x467_outr_UnitPipe.scala 48:23:@40208.4]
  assign x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x250_TVALID = io_in_x250_TVALID; // @[sm_x467_outr_UnitPipe.scala 49:23:@40218.4]
  assign x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x250_TDATA = io_in_x250_TDATA; // @[sm_x467_outr_UnitPipe.scala 49:23:@40216.4]
  assign x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x250_TID = io_in_x250_TID; // @[sm_x467_outr_UnitPipe.scala 49:23:@40212.4]
  assign x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_in_x250_TDEST = io_in_x250_TDEST; // @[sm_x467_outr_UnitPipe.scala 49:23:@40211.4]
  assign x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x467_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x467_outr_UnitPipe.scala 92:22:@40234.4]
  assign x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x467_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x467_outr_UnitPipe.scala 92:22:@40235.4]
  assign x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x467_outr_UnitPipe_sm_io_childAck_0; // @[sm_x467_outr_UnitPipe.scala 92:22:@40230.4]
  assign x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x467_outr_UnitPipe_sm_io_childAck_1; // @[sm_x467_outr_UnitPipe.scala 92:22:@40231.4]
  assign x467_outr_UnitPipe_kernelx467_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x467_outr_UnitPipe.scala 91:18:@40219.4]
  assign x489_outr_UnitPipe_sm_clock = clock; // @[:@40319.4]
  assign x489_outr_UnitPipe_sm_reset = reset; // @[:@40320.4]
  assign x489_outr_UnitPipe_sm_io_enable = _T_508 & _T_517; // @[SpatialBlocks.scala 140:18:@40410.4]
  assign x489_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@40412.4]
  assign x489_outr_UnitPipe_sm_io_doneIn_0 = x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@40378.4]
  assign x489_outr_UnitPipe_sm_io_doneIn_1 = x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@40379.4]
  assign x489_outr_UnitPipe_sm_io_doneIn_2 = x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:67:@40380.4]
  assign x489_outr_UnitPipe_sm_io_ctrCopyDone_0 = x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@40427.4]
  assign x489_outr_UnitPipe_sm_io_ctrCopyDone_1 = x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@40428.4]
  assign x489_outr_UnitPipe_sm_io_ctrCopyDone_2 = x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[SpatialBlocks.scala 161:90:@40429.4]
  assign RetimeWrapper_2_clock = clock; // @[:@40391.4]
  assign RetimeWrapper_2_reset = reset; // @[:@40392.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@40394.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@40393.4]
  assign RetimeWrapper_3_clock = clock; // @[:@40399.4]
  assign RetimeWrapper_3_reset = reset; // @[:@40400.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@40402.4]
  assign RetimeWrapper_3_io_in = x489_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@40401.4]
  assign x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_clock = clock; // @[:@40431.4]
  assign x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_reset = reset; // @[:@40432.4]
  assign x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x468_ready = io_in_x468_ready; // @[sm_x489_outr_UnitPipe.scala 58:23:@40513.4]
  assign x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x248_outdram_number = io_in_x248_outdram_number; // @[sm_x489_outr_UnitPipe.scala 59:31:@40514.4]
  assign x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x252_outbuf_0_rPort_0_output_0 = io_in_x252_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@40515.4]
  assign x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x470_valid = io_in_x470_valid; // @[sm_x489_outr_UnitPipe.scala 61:23:@40521.4]
  assign x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_in_x469_ready = io_in_x469_ready; // @[sm_x489_outr_UnitPipe.scala 62:23:@40526.4]
  assign x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x489_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x489_outr_UnitPipe.scala 113:22:@40549.4]
  assign x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x489_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x489_outr_UnitPipe.scala 113:22:@40550.4]
  assign x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2 = x489_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x489_outr_UnitPipe.scala 113:22:@40551.4]
  assign x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x489_outr_UnitPipe_sm_io_childAck_0; // @[sm_x489_outr_UnitPipe.scala 113:22:@40543.4]
  assign x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x489_outr_UnitPipe_sm_io_childAck_1; // @[sm_x489_outr_UnitPipe.scala 113:22:@40544.4]
  assign x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2 = x489_outr_UnitPipe_sm_io_childAck_2; // @[sm_x489_outr_UnitPipe.scala 113:22:@40545.4]
  assign x489_outr_UnitPipe_kernelx489_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x489_outr_UnitPipe.scala 112:18:@40527.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@40579.2]
  input          clock, // @[:@40580.4]
  input          reset, // @[:@40581.4]
  input          io_in_x468_ready, // @[:@40582.4]
  output         io_in_x468_valid, // @[:@40582.4]
  output [63:0]  io_in_x468_bits_addr, // @[:@40582.4]
  output [31:0]  io_in_x468_bits_size, // @[:@40582.4]
  input  [63:0]  io_in_x248_outdram_number, // @[:@40582.4]
  output         io_in_x251_TVALID, // @[:@40582.4]
  input          io_in_x251_TREADY, // @[:@40582.4]
  output [255:0] io_in_x251_TDATA, // @[:@40582.4]
  output         io_in_x470_ready, // @[:@40582.4]
  input          io_in_x470_valid, // @[:@40582.4]
  input          io_in_x250_TVALID, // @[:@40582.4]
  output         io_in_x250_TREADY, // @[:@40582.4]
  input  [255:0] io_in_x250_TDATA, // @[:@40582.4]
  input  [7:0]   io_in_x250_TID, // @[:@40582.4]
  input  [7:0]   io_in_x250_TDEST, // @[:@40582.4]
  input          io_in_x469_ready, // @[:@40582.4]
  output         io_in_x469_valid, // @[:@40582.4]
  output [31:0]  io_in_x469_bits_wdata_0, // @[:@40582.4]
  output         io_in_x469_bits_wstrb, // @[:@40582.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@40582.4]
  input          io_sigsIn_smChildAcks_0, // @[:@40582.4]
  output         io_sigsOut_smDoneIn_0, // @[:@40582.4]
  input          io_rr // @[:@40582.4]
);
  wire  x252_outbuf_0_clock; // @[m_x252_outbuf_0.scala 27:17:@40592.4]
  wire  x252_outbuf_0_reset; // @[m_x252_outbuf_0.scala 27:17:@40592.4]
  wire [20:0] x252_outbuf_0_io_rPort_0_ofs_0; // @[m_x252_outbuf_0.scala 27:17:@40592.4]
  wire  x252_outbuf_0_io_rPort_0_en_0; // @[m_x252_outbuf_0.scala 27:17:@40592.4]
  wire  x252_outbuf_0_io_rPort_0_backpressure; // @[m_x252_outbuf_0.scala 27:17:@40592.4]
  wire [31:0] x252_outbuf_0_io_rPort_0_output_0; // @[m_x252_outbuf_0.scala 27:17:@40592.4]
  wire  x538_sm_clock; // @[sm_x538.scala 37:18:@40650.4]
  wire  x538_sm_reset; // @[sm_x538.scala 37:18:@40650.4]
  wire  x538_sm_io_enable; // @[sm_x538.scala 37:18:@40650.4]
  wire  x538_sm_io_done; // @[sm_x538.scala 37:18:@40650.4]
  wire  x538_sm_io_ctrDone; // @[sm_x538.scala 37:18:@40650.4]
  wire  x538_sm_io_ctrInc; // @[sm_x538.scala 37:18:@40650.4]
  wire  x538_sm_io_parentAck; // @[sm_x538.scala 37:18:@40650.4]
  wire  x538_sm_io_doneIn_0; // @[sm_x538.scala 37:18:@40650.4]
  wire  x538_sm_io_doneIn_1; // @[sm_x538.scala 37:18:@40650.4]
  wire  x538_sm_io_enableOut_0; // @[sm_x538.scala 37:18:@40650.4]
  wire  x538_sm_io_enableOut_1; // @[sm_x538.scala 37:18:@40650.4]
  wire  x538_sm_io_childAck_0; // @[sm_x538.scala 37:18:@40650.4]
  wire  x538_sm_io_childAck_1; // @[sm_x538.scala 37:18:@40650.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@40717.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@40717.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@40717.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@40717.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@40717.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@40725.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@40725.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@40725.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@40725.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@40725.4]
  wire  x538_kernelx538_concrete1_clock; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_reset; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_in_x468_ready; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_in_x468_valid; // @[sm_x538.scala 102:24:@40754.4]
  wire [63:0] x538_kernelx538_concrete1_io_in_x468_bits_addr; // @[sm_x538.scala 102:24:@40754.4]
  wire [31:0] x538_kernelx538_concrete1_io_in_x468_bits_size; // @[sm_x538.scala 102:24:@40754.4]
  wire [63:0] x538_kernelx538_concrete1_io_in_x248_outdram_number; // @[sm_x538.scala 102:24:@40754.4]
  wire [20:0] x538_kernelx538_concrete1_io_in_x252_outbuf_0_rPort_0_ofs_0; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_in_x252_outbuf_0_rPort_0_en_0; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_in_x252_outbuf_0_rPort_0_backpressure; // @[sm_x538.scala 102:24:@40754.4]
  wire [31:0] x538_kernelx538_concrete1_io_in_x252_outbuf_0_rPort_0_output_0; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_in_x251_TVALID; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_in_x251_TREADY; // @[sm_x538.scala 102:24:@40754.4]
  wire [255:0] x538_kernelx538_concrete1_io_in_x251_TDATA; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_in_x470_ready; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_in_x470_valid; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_in_x250_TVALID; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_in_x250_TREADY; // @[sm_x538.scala 102:24:@40754.4]
  wire [255:0] x538_kernelx538_concrete1_io_in_x250_TDATA; // @[sm_x538.scala 102:24:@40754.4]
  wire [7:0] x538_kernelx538_concrete1_io_in_x250_TID; // @[sm_x538.scala 102:24:@40754.4]
  wire [7:0] x538_kernelx538_concrete1_io_in_x250_TDEST; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_in_x469_ready; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_in_x469_valid; // @[sm_x538.scala 102:24:@40754.4]
  wire [31:0] x538_kernelx538_concrete1_io_in_x469_bits_wdata_0; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_in_x469_bits_wstrb; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x538.scala 102:24:@40754.4]
  wire  x538_kernelx538_concrete1_io_rr; // @[sm_x538.scala 102:24:@40754.4]
  wire  _T_266; // @[package.scala 100:49:@40683.4]
  reg  _T_269; // @[package.scala 48:56:@40684.4]
  reg [31:0] _RAND_0;
  wire  _T_283; // @[package.scala 96:25:@40722.4 package.scala 96:25:@40723.4]
  wire  _T_289; // @[package.scala 96:25:@40730.4 package.scala 96:25:@40731.4]
  wire  _T_292; // @[SpatialBlocks.scala 138:93:@40733.4]
  x252_outbuf_0 x252_outbuf_0 ( // @[m_x252_outbuf_0.scala 27:17:@40592.4]
    .clock(x252_outbuf_0_clock),
    .reset(x252_outbuf_0_reset),
    .io_rPort_0_ofs_0(x252_outbuf_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x252_outbuf_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x252_outbuf_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x252_outbuf_0_io_rPort_0_output_0)
  );
  x538_sm x538_sm ( // @[sm_x538.scala 37:18:@40650.4]
    .clock(x538_sm_clock),
    .reset(x538_sm_reset),
    .io_enable(x538_sm_io_enable),
    .io_done(x538_sm_io_done),
    .io_ctrDone(x538_sm_io_ctrDone),
    .io_ctrInc(x538_sm_io_ctrInc),
    .io_parentAck(x538_sm_io_parentAck),
    .io_doneIn_0(x538_sm_io_doneIn_0),
    .io_doneIn_1(x538_sm_io_doneIn_1),
    .io_enableOut_0(x538_sm_io_enableOut_0),
    .io_enableOut_1(x538_sm_io_enableOut_1),
    .io_childAck_0(x538_sm_io_childAck_0),
    .io_childAck_1(x538_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@40717.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@40725.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x538_kernelx538_concrete1 x538_kernelx538_concrete1 ( // @[sm_x538.scala 102:24:@40754.4]
    .clock(x538_kernelx538_concrete1_clock),
    .reset(x538_kernelx538_concrete1_reset),
    .io_in_x468_ready(x538_kernelx538_concrete1_io_in_x468_ready),
    .io_in_x468_valid(x538_kernelx538_concrete1_io_in_x468_valid),
    .io_in_x468_bits_addr(x538_kernelx538_concrete1_io_in_x468_bits_addr),
    .io_in_x468_bits_size(x538_kernelx538_concrete1_io_in_x468_bits_size),
    .io_in_x248_outdram_number(x538_kernelx538_concrete1_io_in_x248_outdram_number),
    .io_in_x252_outbuf_0_rPort_0_ofs_0(x538_kernelx538_concrete1_io_in_x252_outbuf_0_rPort_0_ofs_0),
    .io_in_x252_outbuf_0_rPort_0_en_0(x538_kernelx538_concrete1_io_in_x252_outbuf_0_rPort_0_en_0),
    .io_in_x252_outbuf_0_rPort_0_backpressure(x538_kernelx538_concrete1_io_in_x252_outbuf_0_rPort_0_backpressure),
    .io_in_x252_outbuf_0_rPort_0_output_0(x538_kernelx538_concrete1_io_in_x252_outbuf_0_rPort_0_output_0),
    .io_in_x251_TVALID(x538_kernelx538_concrete1_io_in_x251_TVALID),
    .io_in_x251_TREADY(x538_kernelx538_concrete1_io_in_x251_TREADY),
    .io_in_x251_TDATA(x538_kernelx538_concrete1_io_in_x251_TDATA),
    .io_in_x470_ready(x538_kernelx538_concrete1_io_in_x470_ready),
    .io_in_x470_valid(x538_kernelx538_concrete1_io_in_x470_valid),
    .io_in_x250_TVALID(x538_kernelx538_concrete1_io_in_x250_TVALID),
    .io_in_x250_TREADY(x538_kernelx538_concrete1_io_in_x250_TREADY),
    .io_in_x250_TDATA(x538_kernelx538_concrete1_io_in_x250_TDATA),
    .io_in_x250_TID(x538_kernelx538_concrete1_io_in_x250_TID),
    .io_in_x250_TDEST(x538_kernelx538_concrete1_io_in_x250_TDEST),
    .io_in_x469_ready(x538_kernelx538_concrete1_io_in_x469_ready),
    .io_in_x469_valid(x538_kernelx538_concrete1_io_in_x469_valid),
    .io_in_x469_bits_wdata_0(x538_kernelx538_concrete1_io_in_x469_bits_wdata_0),
    .io_in_x469_bits_wstrb(x538_kernelx538_concrete1_io_in_x469_bits_wstrb),
    .io_sigsIn_smEnableOuts_0(x538_kernelx538_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x538_kernelx538_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x538_kernelx538_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x538_kernelx538_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x538_kernelx538_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x538_kernelx538_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(x538_kernelx538_concrete1_io_rr)
  );
  assign _T_266 = x538_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@40683.4]
  assign _T_283 = RetimeWrapper_io_out; // @[package.scala 96:25:@40722.4 package.scala 96:25:@40723.4]
  assign _T_289 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@40730.4 package.scala 96:25:@40731.4]
  assign _T_292 = ~ _T_289; // @[SpatialBlocks.scala 138:93:@40733.4]
  assign io_in_x468_valid = x538_kernelx538_concrete1_io_in_x468_valid; // @[sm_x538.scala 63:23:@40835.4]
  assign io_in_x468_bits_addr = x538_kernelx538_concrete1_io_in_x468_bits_addr; // @[sm_x538.scala 63:23:@40834.4]
  assign io_in_x468_bits_size = x538_kernelx538_concrete1_io_in_x468_bits_size; // @[sm_x538.scala 63:23:@40833.4]
  assign io_in_x251_TVALID = x538_kernelx538_concrete1_io_in_x251_TVALID; // @[sm_x538.scala 66:23:@40851.4]
  assign io_in_x251_TDATA = x538_kernelx538_concrete1_io_in_x251_TDATA; // @[sm_x538.scala 66:23:@40849.4]
  assign io_in_x470_ready = x538_kernelx538_concrete1_io_in_x470_ready; // @[sm_x538.scala 67:23:@40854.4]
  assign io_in_x250_TREADY = x538_kernelx538_concrete1_io_in_x250_TREADY; // @[sm_x538.scala 68:23:@40862.4]
  assign io_in_x469_valid = x538_kernelx538_concrete1_io_in_x469_valid; // @[sm_x538.scala 69:23:@40866.4]
  assign io_in_x469_bits_wdata_0 = x538_kernelx538_concrete1_io_in_x469_bits_wdata_0; // @[sm_x538.scala 69:23:@40865.4]
  assign io_in_x469_bits_wstrb = x538_kernelx538_concrete1_io_in_x469_bits_wstrb; // @[sm_x538.scala 69:23:@40864.4]
  assign io_sigsOut_smDoneIn_0 = x538_sm_io_done; // @[SpatialBlocks.scala 156:53:@40740.4]
  assign x252_outbuf_0_clock = clock; // @[:@40593.4]
  assign x252_outbuf_0_reset = reset; // @[:@40594.4]
  assign x252_outbuf_0_io_rPort_0_ofs_0 = x538_kernelx538_concrete1_io_in_x252_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@40841.4]
  assign x252_outbuf_0_io_rPort_0_en_0 = x538_kernelx538_concrete1_io_in_x252_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@40840.4]
  assign x252_outbuf_0_io_rPort_0_backpressure = x538_kernelx538_concrete1_io_in_x252_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@40839.4]
  assign x538_sm_clock = clock; // @[:@40651.4]
  assign x538_sm_reset = reset; // @[:@40652.4]
  assign x538_sm_io_enable = _T_283 & _T_292; // @[SpatialBlocks.scala 140:18:@40737.4]
  assign x538_sm_io_ctrDone = x538_sm_io_ctrInc & _T_269; // @[sm_RootController.scala 82:26:@40687.4]
  assign x538_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@40739.4]
  assign x538_sm_io_doneIn_0 = x538_kernelx538_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@40707.4]
  assign x538_sm_io_doneIn_1 = x538_kernelx538_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@40708.4]
  assign RetimeWrapper_clock = clock; // @[:@40718.4]
  assign RetimeWrapper_reset = reset; // @[:@40719.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@40721.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@40720.4]
  assign RetimeWrapper_1_clock = clock; // @[:@40726.4]
  assign RetimeWrapper_1_reset = reset; // @[:@40727.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@40729.4]
  assign RetimeWrapper_1_io_in = x538_sm_io_done; // @[package.scala 94:16:@40728.4]
  assign x538_kernelx538_concrete1_clock = clock; // @[:@40755.4]
  assign x538_kernelx538_concrete1_reset = reset; // @[:@40756.4]
  assign x538_kernelx538_concrete1_io_in_x468_ready = io_in_x468_ready; // @[sm_x538.scala 63:23:@40836.4]
  assign x538_kernelx538_concrete1_io_in_x248_outdram_number = io_in_x248_outdram_number; // @[sm_x538.scala 64:31:@40837.4]
  assign x538_kernelx538_concrete1_io_in_x252_outbuf_0_rPort_0_output_0 = x252_outbuf_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@40838.4]
  assign x538_kernelx538_concrete1_io_in_x251_TREADY = io_in_x251_TREADY; // @[sm_x538.scala 66:23:@40850.4]
  assign x538_kernelx538_concrete1_io_in_x470_valid = io_in_x470_valid; // @[sm_x538.scala 67:23:@40853.4]
  assign x538_kernelx538_concrete1_io_in_x250_TVALID = io_in_x250_TVALID; // @[sm_x538.scala 68:23:@40863.4]
  assign x538_kernelx538_concrete1_io_in_x250_TDATA = io_in_x250_TDATA; // @[sm_x538.scala 68:23:@40861.4]
  assign x538_kernelx538_concrete1_io_in_x250_TID = io_in_x250_TID; // @[sm_x538.scala 68:23:@40857.4]
  assign x538_kernelx538_concrete1_io_in_x250_TDEST = io_in_x250_TDEST; // @[sm_x538.scala 68:23:@40856.4]
  assign x538_kernelx538_concrete1_io_in_x469_ready = io_in_x469_ready; // @[sm_x538.scala 69:23:@40867.4]
  assign x538_kernelx538_concrete1_io_sigsIn_smEnableOuts_0 = x538_sm_io_enableOut_0; // @[sm_x538.scala 107:22:@40878.4]
  assign x538_kernelx538_concrete1_io_sigsIn_smEnableOuts_1 = x538_sm_io_enableOut_1; // @[sm_x538.scala 107:22:@40879.4]
  assign x538_kernelx538_concrete1_io_sigsIn_smChildAcks_0 = x538_sm_io_childAck_0; // @[sm_x538.scala 107:22:@40874.4]
  assign x538_kernelx538_concrete1_io_sigsIn_smChildAcks_1 = x538_sm_io_childAck_1; // @[sm_x538.scala 107:22:@40875.4]
  assign x538_kernelx538_concrete1_io_rr = io_rr; // @[sm_x538.scala 106:18:@40868.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_269 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_269 <= 1'h0;
    end else begin
      _T_269 <= _T_266;
    end
  end
endmodule
module AccelUnit( // @[:@40901.2]
  input          clock, // @[:@40902.4]
  input          reset, // @[:@40903.4]
  input          io_enable, // @[:@40904.4]
  output         io_done, // @[:@40904.4]
  input          io_reset, // @[:@40904.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@40904.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@40904.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@40904.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@40904.4]
  output         io_memStreams_loads_0_data_ready, // @[:@40904.4]
  input          io_memStreams_loads_0_data_valid, // @[:@40904.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@40904.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@40904.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@40904.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@40904.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@40904.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@40904.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@40904.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@40904.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@40904.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@40904.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@40904.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@40904.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@40904.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@40904.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@40904.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@40904.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@40904.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@40904.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@40904.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@40904.4]
  input          io_memStreams_stores_0_data_ready, // @[:@40904.4]
  output         io_memStreams_stores_0_data_valid, // @[:@40904.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@40904.4]
  output         io_memStreams_stores_0_data_bits_wstrb, // @[:@40904.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@40904.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@40904.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@40904.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@40904.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@40904.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@40904.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@40904.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@40904.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@40904.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@40904.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@40904.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@40904.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@40904.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@40904.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@40904.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@40904.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@40904.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@40904.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@40904.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@40904.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@40904.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@40904.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@40904.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@40904.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@40904.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@40904.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@40904.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@40904.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@40904.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@40904.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@40904.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@40904.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@40904.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@40904.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@40904.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@40904.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@40904.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@40904.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@40904.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@40904.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@40904.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@40904.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@40904.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@40904.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@40904.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@40904.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@40904.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@40904.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@40904.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@40904.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@40904.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@40904.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@40904.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@40904.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@40904.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@40904.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@40904.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@40904.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@40904.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@40904.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@40904.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@40904.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@40904.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@40904.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@40904.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@40904.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@40904.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@40904.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@40904.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@40904.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@40904.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@40904.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@40904.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@40904.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@40904.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@40904.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@40904.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@40904.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@40904.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@40904.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@40904.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@40904.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@40904.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@40904.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@40904.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@40904.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@40904.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@40904.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@40904.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@40904.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@40904.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@40904.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@40904.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@40904.4]
  output         io_heap_0_req_valid, // @[:@40904.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@40904.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@40904.4]
  input          io_heap_0_resp_valid, // @[:@40904.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@40904.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@40904.4]
  input  [63:0]  io_argIns_0, // @[:@40904.4]
  input  [63:0]  io_argIns_1, // @[:@40904.4]
  input          io_argOuts_0_port_ready, // @[:@40904.4]
  output         io_argOuts_0_port_valid, // @[:@40904.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@40904.4]
  input  [63:0]  io_argOuts_0_echo // @[:@40904.4]
);
  wire  SingleCounter_clock; // @[Main.scala 40:32:@41052.4]
  wire  SingleCounter_reset; // @[Main.scala 40:32:@41052.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 40:32:@41052.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 40:32:@41052.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@41070.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@41070.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@41070.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@41070.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@41070.4]
  wire  SRFF_clock; // @[Main.scala 44:28:@41079.4]
  wire  SRFF_reset; // @[Main.scala 44:28:@41079.4]
  wire  SRFF_io_input_set; // @[Main.scala 44:28:@41079.4]
  wire  SRFF_io_input_reset; // @[Main.scala 44:28:@41079.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 44:28:@41079.4]
  wire  SRFF_io_output; // @[Main.scala 44:28:@41079.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 36:18:@41118.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 36:18:@41118.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 36:18:@41118.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 36:18:@41118.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 36:18:@41118.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 36:18:@41118.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 36:18:@41118.4]
  wire  RootController_sm_io_parentAck; // @[sm_RootController.scala 36:18:@41118.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 36:18:@41118.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 36:18:@41118.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 36:18:@41118.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@41150.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@41150.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@41150.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@41150.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@41150.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 91:24:@41212.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 91:24:@41212.4]
  wire  RootController_kernelRootController_concrete1_io_in_x468_ready; // @[sm_RootController.scala 91:24:@41212.4]
  wire  RootController_kernelRootController_concrete1_io_in_x468_valid; // @[sm_RootController.scala 91:24:@41212.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x468_bits_addr; // @[sm_RootController.scala 91:24:@41212.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x468_bits_size; // @[sm_RootController.scala 91:24:@41212.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x248_outdram_number; // @[sm_RootController.scala 91:24:@41212.4]
  wire  RootController_kernelRootController_concrete1_io_in_x251_TVALID; // @[sm_RootController.scala 91:24:@41212.4]
  wire  RootController_kernelRootController_concrete1_io_in_x251_TREADY; // @[sm_RootController.scala 91:24:@41212.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x251_TDATA; // @[sm_RootController.scala 91:24:@41212.4]
  wire  RootController_kernelRootController_concrete1_io_in_x470_ready; // @[sm_RootController.scala 91:24:@41212.4]
  wire  RootController_kernelRootController_concrete1_io_in_x470_valid; // @[sm_RootController.scala 91:24:@41212.4]
  wire  RootController_kernelRootController_concrete1_io_in_x250_TVALID; // @[sm_RootController.scala 91:24:@41212.4]
  wire  RootController_kernelRootController_concrete1_io_in_x250_TREADY; // @[sm_RootController.scala 91:24:@41212.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x250_TDATA; // @[sm_RootController.scala 91:24:@41212.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x250_TID; // @[sm_RootController.scala 91:24:@41212.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x250_TDEST; // @[sm_RootController.scala 91:24:@41212.4]
  wire  RootController_kernelRootController_concrete1_io_in_x469_ready; // @[sm_RootController.scala 91:24:@41212.4]
  wire  RootController_kernelRootController_concrete1_io_in_x469_valid; // @[sm_RootController.scala 91:24:@41212.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x469_bits_wdata_0; // @[sm_RootController.scala 91:24:@41212.4]
  wire  RootController_kernelRootController_concrete1_io_in_x469_bits_wstrb; // @[sm_RootController.scala 91:24:@41212.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 91:24:@41212.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 91:24:@41212.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 91:24:@41212.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 91:24:@41212.4]
  wire  _T_599; // @[package.scala 96:25:@41075.4 package.scala 96:25:@41076.4]
  wire  _T_664; // @[Main.scala 46:50:@41146.4]
  wire  _T_665; // @[Main.scala 46:59:@41147.4]
  wire  _T_677; // @[package.scala 100:49:@41167.4]
  reg  _T_680; // @[package.scala 48:56:@41168.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 40:32:@41052.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@41070.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 44:28:@41079.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 36:18:@41118.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_parentAck(RootController_sm_io_parentAck),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@41150.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 91:24:@41212.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x468_ready(RootController_kernelRootController_concrete1_io_in_x468_ready),
    .io_in_x468_valid(RootController_kernelRootController_concrete1_io_in_x468_valid),
    .io_in_x468_bits_addr(RootController_kernelRootController_concrete1_io_in_x468_bits_addr),
    .io_in_x468_bits_size(RootController_kernelRootController_concrete1_io_in_x468_bits_size),
    .io_in_x248_outdram_number(RootController_kernelRootController_concrete1_io_in_x248_outdram_number),
    .io_in_x251_TVALID(RootController_kernelRootController_concrete1_io_in_x251_TVALID),
    .io_in_x251_TREADY(RootController_kernelRootController_concrete1_io_in_x251_TREADY),
    .io_in_x251_TDATA(RootController_kernelRootController_concrete1_io_in_x251_TDATA),
    .io_in_x470_ready(RootController_kernelRootController_concrete1_io_in_x470_ready),
    .io_in_x470_valid(RootController_kernelRootController_concrete1_io_in_x470_valid),
    .io_in_x250_TVALID(RootController_kernelRootController_concrete1_io_in_x250_TVALID),
    .io_in_x250_TREADY(RootController_kernelRootController_concrete1_io_in_x250_TREADY),
    .io_in_x250_TDATA(RootController_kernelRootController_concrete1_io_in_x250_TDATA),
    .io_in_x250_TID(RootController_kernelRootController_concrete1_io_in_x250_TID),
    .io_in_x250_TDEST(RootController_kernelRootController_concrete1_io_in_x250_TDEST),
    .io_in_x469_ready(RootController_kernelRootController_concrete1_io_in_x469_ready),
    .io_in_x469_valid(RootController_kernelRootController_concrete1_io_in_x469_valid),
    .io_in_x469_bits_wdata_0(RootController_kernelRootController_concrete1_io_in_x469_bits_wdata_0),
    .io_in_x469_bits_wstrb(RootController_kernelRootController_concrete1_io_in_x469_bits_wstrb),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@41075.4 package.scala 96:25:@41076.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 46:50:@41146.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 46:59:@41147.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@41167.4]
  assign io_done = SRFF_io_output; // @[Main.scala 53:23:@41166.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x468_valid; // @[sm_RootController.scala 60:23:@41275.4]
  assign io_memStreams_stores_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x468_bits_addr; // @[sm_RootController.scala 60:23:@41274.4]
  assign io_memStreams_stores_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x468_bits_size; // @[sm_RootController.scala 60:23:@41273.4]
  assign io_memStreams_stores_0_data_valid = RootController_kernelRootController_concrete1_io_in_x469_valid; // @[sm_RootController.scala 65:23:@41301.4]
  assign io_memStreams_stores_0_data_bits_wdata_0 = RootController_kernelRootController_concrete1_io_in_x469_bits_wdata_0; // @[sm_RootController.scala 65:23:@41300.4]
  assign io_memStreams_stores_0_data_bits_wstrb = RootController_kernelRootController_concrete1_io_in_x469_bits_wstrb; // @[sm_RootController.scala 65:23:@41299.4]
  assign io_memStreams_stores_0_wresp_ready = RootController_kernelRootController_concrete1_io_in_x470_ready; // @[sm_RootController.scala 63:23:@41289.4]
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x250_TREADY; // @[sm_RootController.scala 64:23:@41297.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x251_TVALID; // @[sm_RootController.scala 62:23:@41286.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x251_TDATA; // @[sm_RootController.scala 62:23:@41284.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 62:23:@41283.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 62:23:@41282.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 62:23:@41281.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 62:23:@41280.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 62:23:@41279.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 62:23:@41278.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@41053.4]
  assign SingleCounter_reset = reset; // @[:@41054.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 41:79:@41068.4]
  assign RetimeWrapper_clock = clock; // @[:@41071.4]
  assign RetimeWrapper_reset = reset; // @[:@41072.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@41074.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@41073.4]
  assign SRFF_clock = clock; // @[:@41080.4]
  assign SRFF_reset = reset; // @[:@41081.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 62:29:@41330.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 51:31:@41164.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 52:36:@41165.4]
  assign RootController_sm_clock = clock; // @[:@41119.4]
  assign RootController_sm_reset = reset; // @[:@41120.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 50:33:@41163.4 SpatialBlocks.scala 140:18:@41197.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@41191.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 54:34:@41171.4]
  assign RootController_sm_io_parentAck = 1'h0; // @[Main.scala 49:36:@41159.4 SpatialBlocks.scala 142:21:@41199.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@41188.4]
  assign RetimeWrapper_1_clock = clock; // @[:@41151.4]
  assign RetimeWrapper_1_reset = reset; // @[:@41152.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@41154.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@41153.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@41213.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@41214.4]
  assign RootController_kernelRootController_concrete1_io_in_x468_ready = io_memStreams_stores_0_cmd_ready; // @[sm_RootController.scala 60:23:@41276.4]
  assign RootController_kernelRootController_concrete1_io_in_x248_outdram_number = io_argIns_1; // @[sm_RootController.scala 61:31:@41277.4]
  assign RootController_kernelRootController_concrete1_io_in_x251_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 62:23:@41285.4]
  assign RootController_kernelRootController_concrete1_io_in_x470_valid = io_memStreams_stores_0_wresp_valid; // @[sm_RootController.scala 63:23:@41288.4]
  assign RootController_kernelRootController_concrete1_io_in_x250_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 64:23:@41298.4]
  assign RootController_kernelRootController_concrete1_io_in_x250_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 64:23:@41296.4]
  assign RootController_kernelRootController_concrete1_io_in_x250_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 64:23:@41292.4]
  assign RootController_kernelRootController_concrete1_io_in_x250_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 64:23:@41291.4]
  assign RootController_kernelRootController_concrete1_io_in_x469_ready = io_memStreams_stores_0_data_ready; // @[sm_RootController.scala 65:23:@41302.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 96:22:@41311.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 96:22:@41309.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 95:18:@41303.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module Counter( // @[:@41332.2]
  input        clock, // @[:@41333.4]
  input        reset, // @[:@41334.4]
  input        io_enable, // @[:@41335.4]
  output [5:0] io_out, // @[:@41335.4]
  output [5:0] io_next // @[:@41335.4]
);
  reg [5:0] count; // @[Counter.scala 15:22:@41337.4]
  reg [31:0] _RAND_0;
  wire [6:0] _T_17; // @[Counter.scala 17:24:@41338.4]
  wire [5:0] newCount; // @[Counter.scala 17:24:@41339.4]
  wire [5:0] _GEN_0; // @[Counter.scala 21:26:@41344.6]
  assign _T_17 = count + 6'h1; // @[Counter.scala 17:24:@41338.4]
  assign newCount = count + 6'h1; // @[Counter.scala 17:24:@41339.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@41344.6]
  assign io_out = count; // @[Counter.scala 25:10:@41347.4]
  assign io_next = count + 6'h1; // @[Counter.scala 26:11:@41348.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 6'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module SRAM_33( // @[:@41384.2]
  input         clock, // @[:@41385.4]
  input         reset, // @[:@41386.4]
  input  [5:0]  io_raddr, // @[:@41387.4]
  input         io_wen, // @[:@41387.4]
  input  [5:0]  io_waddr, // @[:@41387.4]
  input  [63:0] io_wdata_addr, // @[:@41387.4]
  input  [31:0] io_wdata_size, // @[:@41387.4]
  output [63:0] io_rdata_addr, // @[:@41387.4]
  output [31:0] io_rdata_size // @[:@41387.4]
);
  wire [95:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@41389.4]
  wire [95:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@41389.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@41389.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@41389.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@41389.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@41389.4]
  wire [5:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@41389.4]
  wire [5:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@41389.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@41389.4]
  wire [95:0] _T_17; // @[SRAM.scala 175:38:@41403.4]
  wire  _T_20; // @[SRAM.scala 182:49:@41408.4]
  wire  _T_21; // @[SRAM.scala 182:37:@41409.4]
  reg  _T_24; // @[SRAM.scala 182:29:@41410.4]
  reg [31:0] _RAND_0;
  reg [95:0] _T_28; // @[SRAM.scala 183:29:@41413.4]
  reg [95:0] _RAND_1;
  wire [95:0] _T_29; // @[SRAM.scala 184:22:@41415.4]
  SRAMVerilogAWS #(.DWIDTH(96), .WORDS(64), .AWIDTH(6)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@41389.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_17 = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:38:@41403.4]
  assign _T_20 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@41408.4]
  assign _T_21 = io_wen & _T_20; // @[SRAM.scala 182:37:@41409.4]
  assign _T_29 = _T_24 ? _T_28 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:22:@41415.4]
  assign io_rdata_addr = _T_29[95:32]; // @[SRAM.scala 184:16:@41424.4]
  assign io_rdata_size = _T_29[31:0]; // @[SRAM.scala 184:16:@41423.4]
  assign SRAMVerilogAWS_wdata = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:20:@41404.4]
  assign SRAMVerilogAWS_backpressure = 1'h1; // @[SRAM.scala 176:27:@41405.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@41401.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@41407.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@41406.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@41402.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@41400.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@41399.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_24 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  _T_28 = _RAND_1[95:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_24 <= 1'h0;
    end else begin
      _T_24 <= _T_21;
    end
    if (reset) begin
      _T_28 <= 96'h0;
    end else begin
      _T_28 <= _T_17;
    end
  end
endmodule
module FIFO( // @[:@41426.2]
  input         clock, // @[:@41427.4]
  input         reset, // @[:@41428.4]
  output        io_in_ready, // @[:@41429.4]
  input         io_in_valid, // @[:@41429.4]
  input  [63:0] io_in_bits_addr, // @[:@41429.4]
  input  [31:0] io_in_bits_size, // @[:@41429.4]
  input         io_out_ready, // @[:@41429.4]
  output        io_out_valid, // @[:@41429.4]
  output [63:0] io_out_bits_addr, // @[:@41429.4]
  output [31:0] io_out_bits_size // @[:@41429.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@41825.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@41825.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@41825.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@41825.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@41825.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@41835.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@41835.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@41835.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@41835.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@41835.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@41850.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@41850.4]
  wire [5:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@41850.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@41850.4]
  wire [5:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@41850.4]
  wire [63:0] SRAM_io_wdata_addr; // @[FIFO.scala 73:19:@41850.4]
  wire [31:0] SRAM_io_wdata_size; // @[FIFO.scala 73:19:@41850.4]
  wire [63:0] SRAM_io_rdata_addr; // @[FIFO.scala 73:19:@41850.4]
  wire [31:0] SRAM_io_rdata_size; // @[FIFO.scala 73:19:@41850.4]
  wire  writeEn; // @[FIFO.scala 30:29:@41823.4]
  wire  readEn; // @[FIFO.scala 31:29:@41824.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@41845.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@41846.4]
  wire  _T_824; // @[FIFO.scala 45:27:@41847.4]
  wire  empty; // @[FIFO.scala 45:24:@41848.4]
  wire  full; // @[FIFO.scala 46:23:@41849.4]
  wire  _T_827; // @[FIFO.scala 83:17:@41862.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@41863.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@41825.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@41835.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_33 SRAM ( // @[FIFO.scala 73:19:@41850.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata_addr(SRAM_io_wdata_addr),
    .io_wdata_size(SRAM_io_wdata_size),
    .io_rdata_addr(SRAM_io_rdata_addr),
    .io_rdata_size(SRAM_io_rdata_size)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@41823.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@41824.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@41846.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@41847.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@41848.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@41849.4]
  assign _T_827 = writeEn != readEn; // @[FIFO.scala 83:17:@41862.4]
  assign _GEN_0 = _T_827 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@41863.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@41869.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@41867.4]
  assign io_out_bits_addr = SRAM_io_rdata_addr; // @[FIFO.scala 79:17:@41860.4]
  assign io_out_bits_size = SRAM_io_rdata_size; // @[FIFO.scala 79:17:@41859.4]
  assign enqCounter_clock = clock; // @[:@41826.4]
  assign enqCounter_reset = reset; // @[:@41827.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@41833.4]
  assign deqCounter_clock = clock; // @[:@41836.4]
  assign deqCounter_reset = reset; // @[:@41837.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@41843.4]
  assign SRAM_clock = clock; // @[:@41851.4]
  assign SRAM_reset = reset; // @[:@41852.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@41854.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@41855.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@41856.4]
  assign SRAM_io_wdata_addr = io_in_bits_addr; // @[FIFO.scala 78:16:@41858.4]
  assign SRAM_io_wdata_size = io_in_bits_size; // @[FIFO.scala 78:16:@41857.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_827) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module Counter_2( // @[:@41871.2]
  input        clock, // @[:@41872.4]
  input        reset, // @[:@41873.4]
  input        io_enable, // @[:@41874.4]
  output [3:0] io_out // @[:@41874.4]
);
  reg [3:0] count; // @[Counter.scala 15:22:@41876.4]
  reg [31:0] _RAND_0;
  wire [4:0] _T_17; // @[Counter.scala 17:24:@41877.4]
  wire [3:0] newCount; // @[Counter.scala 17:24:@41878.4]
  wire [3:0] _GEN_0; // @[Counter.scala 21:26:@41883.6]
  assign _T_17 = count + 4'h1; // @[Counter.scala 17:24:@41877.4]
  assign newCount = count + 4'h1; // @[Counter.scala 17:24:@41878.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@41883.6]
  assign io_out = count; // @[Counter.scala 25:10:@41886.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 4'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module Counter_4( // @[:@41907.2]
  input        clock, // @[:@41908.4]
  input        reset, // @[:@41909.4]
  input        io_reset, // @[:@41910.4]
  input        io_enable, // @[:@41910.4]
  input  [1:0] io_stride, // @[:@41910.4]
  output [1:0] io_out, // @[:@41910.4]
  output [1:0] io_next // @[:@41910.4]
);
  reg [1:0] count; // @[Counter.scala 15:22:@41912.4]
  reg [31:0] _RAND_0;
  wire [2:0] _T_17; // @[Counter.scala 17:24:@41913.4]
  wire [1:0] newCount; // @[Counter.scala 17:24:@41914.4]
  wire [1:0] _GEN_0; // @[Counter.scala 21:26:@41919.6]
  wire [1:0] _GEN_1; // @[Counter.scala 19:18:@41915.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@41913.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@41914.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@41919.6]
  assign _GEN_1 = io_reset ? 2'h0 : _GEN_0; // @[Counter.scala 19:18:@41915.4]
  assign io_out = count; // @[Counter.scala 25:10:@41922.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@41923.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 2'h0;
    end else begin
      if (io_reset) begin
        count <= 2'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module SRAM_34( // @[:@41959.2]
  input         clock, // @[:@41960.4]
  input         reset, // @[:@41961.4]
  input  [1:0]  io_raddr, // @[:@41962.4]
  input         io_wen, // @[:@41962.4]
  input  [1:0]  io_waddr, // @[:@41962.4]
  input  [31:0] io_wdata, // @[:@41962.4]
  output [31:0] io_rdata, // @[:@41962.4]
  input         io_backpressure // @[:@41962.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@41964.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@41964.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@41964.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@41964.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@41964.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@41964.4]
  wire [1:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@41964.4]
  wire [1:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@41964.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@41964.4]
  wire  _T_19; // @[SRAM.scala 182:49:@41982.4]
  wire  _T_20; // @[SRAM.scala 182:37:@41983.4]
  reg  _T_23; // @[SRAM.scala 182:29:@41984.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@41986.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(4), .AWIDTH(2)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@41964.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@41982.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@41983.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@41991.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@41978.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@41979.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@41976.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@41981.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@41980.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@41977.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@41975.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@41974.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module FIFO_1( // @[:@41993.2]
  input         clock, // @[:@41994.4]
  input         reset, // @[:@41995.4]
  output        io_in_ready, // @[:@41996.4]
  input         io_in_valid, // @[:@41996.4]
  input  [31:0] io_in_bits, // @[:@41996.4]
  input         io_out_ready, // @[:@41996.4]
  output        io_out_valid, // @[:@41996.4]
  output [31:0] io_out_bits // @[:@41996.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@42022.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@42022.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@42022.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@42022.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@42022.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@42022.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@42022.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@42032.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@42032.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@42032.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@42032.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@42032.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@42032.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@42032.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@42047.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@42047.4]
  wire [1:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@42047.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@42047.4]
  wire [1:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@42047.4]
  wire [31:0] SRAM_io_wdata; // @[FIFO.scala 73:19:@42047.4]
  wire [31:0] SRAM_io_rdata; // @[FIFO.scala 73:19:@42047.4]
  wire  SRAM_io_backpressure; // @[FIFO.scala 73:19:@42047.4]
  wire  writeEn; // @[FIFO.scala 30:29:@42020.4]
  wire  readEn; // @[FIFO.scala 31:29:@42021.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@42042.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@42043.4]
  wire  _T_104; // @[FIFO.scala 45:27:@42044.4]
  wire  empty; // @[FIFO.scala 45:24:@42045.4]
  wire  full; // @[FIFO.scala 46:23:@42046.4]
  wire  _T_107; // @[FIFO.scala 83:17:@42057.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@42058.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@42022.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@42032.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_34 SRAM ( // @[FIFO.scala 73:19:@42047.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@42020.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@42021.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@42043.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@42044.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@42045.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@42046.4]
  assign _T_107 = writeEn != readEn; // @[FIFO.scala 83:17:@42057.4]
  assign _GEN_0 = _T_107 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@42058.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@42064.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@42062.4]
  assign io_out_bits = SRAM_io_rdata; // @[FIFO.scala 79:17:@42055.4]
  assign enqCounter_clock = clock; // @[:@42023.4]
  assign enqCounter_reset = reset; // @[:@42024.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@42030.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@42031.4]
  assign deqCounter_clock = clock; // @[:@42033.4]
  assign deqCounter_reset = reset; // @[:@42034.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@42040.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@42041.4]
  assign SRAM_clock = clock; // @[:@42048.4]
  assign SRAM_reset = reset; // @[:@42049.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@42051.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@42052.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@42053.4]
  assign SRAM_io_wdata = io_in_bits; // @[FIFO.scala 78:16:@42054.4]
  assign SRAM_io_backpressure = 1'h1; // @[FIFO.scala 80:23:@42056.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_107) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec( // @[:@44451.2]
  input         clock, // @[:@44452.4]
  input         reset, // @[:@44453.4]
  output        io_in_ready, // @[:@44454.4]
  input         io_in_valid, // @[:@44454.4]
  input  [31:0] io_in_bits_0, // @[:@44454.4]
  input         io_out_ready, // @[:@44454.4]
  output        io_out_valid, // @[:@44454.4]
  output [31:0] io_out_bits_0, // @[:@44454.4]
  output [31:0] io_out_bits_1, // @[:@44454.4]
  output [31:0] io_out_bits_2, // @[:@44454.4]
  output [31:0] io_out_bits_3, // @[:@44454.4]
  output [31:0] io_out_bits_4, // @[:@44454.4]
  output [31:0] io_out_bits_5, // @[:@44454.4]
  output [31:0] io_out_bits_6, // @[:@44454.4]
  output [31:0] io_out_bits_7, // @[:@44454.4]
  output [31:0] io_out_bits_8, // @[:@44454.4]
  output [31:0] io_out_bits_9, // @[:@44454.4]
  output [31:0] io_out_bits_10, // @[:@44454.4]
  output [31:0] io_out_bits_11, // @[:@44454.4]
  output [31:0] io_out_bits_12, // @[:@44454.4]
  output [31:0] io_out_bits_13, // @[:@44454.4]
  output [31:0] io_out_bits_14, // @[:@44454.4]
  output [31:0] io_out_bits_15 // @[:@44454.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@44458.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@44458.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@44458.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@44458.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@44469.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@44469.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@44469.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@44469.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@44482.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@44482.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@44482.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@44482.4]
  wire [31:0] fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@44482.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@44482.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@44482.4]
  wire [31:0] fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@44482.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@44517.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@44517.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@44517.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@44517.4]
  wire [31:0] fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@44517.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@44517.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@44517.4]
  wire [31:0] fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@44517.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@44552.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@44552.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@44552.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@44552.4]
  wire [31:0] fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@44552.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@44552.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@44552.4]
  wire [31:0] fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@44552.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@44587.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@44587.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@44587.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@44587.4]
  wire [31:0] fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@44587.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@44587.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@44587.4]
  wire [31:0] fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@44587.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@44622.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@44622.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@44622.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@44622.4]
  wire [31:0] fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@44622.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@44622.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@44622.4]
  wire [31:0] fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@44622.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@44657.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@44657.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@44657.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@44657.4]
  wire [31:0] fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@44657.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@44657.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@44657.4]
  wire [31:0] fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@44657.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@44692.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@44692.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@44692.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@44692.4]
  wire [31:0] fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@44692.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@44692.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@44692.4]
  wire [31:0] fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@44692.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@44727.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@44727.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@44727.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@44727.4]
  wire [31:0] fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@44727.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@44727.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@44727.4]
  wire [31:0] fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@44727.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@44762.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@44762.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@44762.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@44762.4]
  wire [31:0] fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@44762.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@44762.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@44762.4]
  wire [31:0] fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@44762.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@44797.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@44797.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@44797.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@44797.4]
  wire [31:0] fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@44797.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@44797.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@44797.4]
  wire [31:0] fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@44797.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@44832.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@44832.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@44832.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@44832.4]
  wire [31:0] fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@44832.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@44832.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@44832.4]
  wire [31:0] fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@44832.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@44867.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@44867.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@44867.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@44867.4]
  wire [31:0] fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@44867.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@44867.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@44867.4]
  wire [31:0] fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@44867.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@44902.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@44902.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@44902.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@44902.4]
  wire [31:0] fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@44902.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@44902.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@44902.4]
  wire [31:0] fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@44902.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@44937.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@44937.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@44937.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@44937.4]
  wire [31:0] fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@44937.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@44937.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@44937.4]
  wire [31:0] fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@44937.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@44972.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@44972.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@44972.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@44972.4]
  wire [31:0] fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@44972.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@44972.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@44972.4]
  wire [31:0] fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@44972.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@45007.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@45007.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@45007.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@45007.4]
  wire [31:0] fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@45007.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@45007.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@45007.4]
  wire [31:0] fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@45007.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@44457.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@44480.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@44507.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@44542.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@44577.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@44612.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@44647.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@44682.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@44717.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@44752.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@44787.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@44822.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@44857.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@44892.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@44927.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@44962.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@44997.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@45032.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45043.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45044.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@45074.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45045.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@45074.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45046.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@45074.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45047.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@45074.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45048.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@45074.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45049.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@45074.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45050.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@45074.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45051.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@45074.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45052.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@45074.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45053.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@45074.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45054.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@45074.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45055.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@45074.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45056.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@45074.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45057.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@45074.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45058.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@45093.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@45094.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@45095.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@45096.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@45097.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@45098.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@45099.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@45100.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@45101.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@45102.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@45103.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@45104.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@45105.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@45106.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@44458.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@44469.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_1 fifos_0 ( // @[FIFOVec.scala 40:19:@44482.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_1 fifos_1 ( // @[FIFOVec.scala 40:19:@44517.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_1 fifos_2 ( // @[FIFOVec.scala 40:19:@44552.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_1 fifos_3 ( // @[FIFOVec.scala 40:19:@44587.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_1 fifos_4 ( // @[FIFOVec.scala 40:19:@44622.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_1 fifos_5 ( // @[FIFOVec.scala 40:19:@44657.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_1 fifos_6 ( // @[FIFOVec.scala 40:19:@44692.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_1 fifos_7 ( // @[FIFOVec.scala 40:19:@44727.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_1 fifos_8 ( // @[FIFOVec.scala 40:19:@44762.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_1 fifos_9 ( // @[FIFOVec.scala 40:19:@44797.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_1 fifos_10 ( // @[FIFOVec.scala 40:19:@44832.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_1 fifos_11 ( // @[FIFOVec.scala 40:19:@44867.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_1 fifos_12 ( // @[FIFOVec.scala 40:19:@44902.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_1 fifos_13 ( // @[FIFOVec.scala 40:19:@44937.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_1 fifos_14 ( // @[FIFOVec.scala 40:19:@44972.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_1 fifos_15 ( // @[FIFOVec.scala 40:19:@45007.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@44457.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@44480.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@44507.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@44542.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@44577.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@44612.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@44647.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@44682.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@44717.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@44752.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@44787.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@44822.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@44857.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@44892.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@44927.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@44962.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@44997.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@45032.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45043.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45044.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@45074.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45045.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@45074.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45046.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@45074.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45047.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@45074.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45048.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@45074.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45049.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@45074.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45050.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@45074.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45051.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@45074.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45052.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@45074.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45053.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@45074.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45054.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@45074.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45055.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@45074.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45056.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@45074.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45057.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@45074.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@45042.4 FIFOVec.scala 49:42:@45058.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@45093.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@45094.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@45095.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@45096.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@45097.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@45098.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@45099.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@45100.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@45101.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@45102.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@45103.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@45104.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@45105.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@45106.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@45075.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@45109.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@45417.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@45418.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@45419.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@45420.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@45421.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@45422.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@45423.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@45424.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@45425.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@45426.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@45427.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@45428.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@45429.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@45430.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@45431.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@45432.4]
  assign enqCounter_clock = clock; // @[:@44459.4]
  assign enqCounter_reset = reset; // @[:@44460.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@44467.4]
  assign deqCounter_clock = clock; // @[:@44470.4]
  assign deqCounter_reset = reset; // @[:@44471.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@44478.4]
  assign fifos_0_clock = clock; // @[:@44483.4]
  assign fifos_0_reset = reset; // @[:@44484.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@44510.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44512.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44516.4]
  assign fifos_1_clock = clock; // @[:@44518.4]
  assign fifos_1_reset = reset; // @[:@44519.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@44545.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44547.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44551.4]
  assign fifos_2_clock = clock; // @[:@44553.4]
  assign fifos_2_reset = reset; // @[:@44554.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@44580.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44582.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44586.4]
  assign fifos_3_clock = clock; // @[:@44588.4]
  assign fifos_3_reset = reset; // @[:@44589.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@44615.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44617.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44621.4]
  assign fifos_4_clock = clock; // @[:@44623.4]
  assign fifos_4_reset = reset; // @[:@44624.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@44650.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44652.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44656.4]
  assign fifos_5_clock = clock; // @[:@44658.4]
  assign fifos_5_reset = reset; // @[:@44659.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@44685.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44687.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44691.4]
  assign fifos_6_clock = clock; // @[:@44693.4]
  assign fifos_6_reset = reset; // @[:@44694.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@44720.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44722.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44726.4]
  assign fifos_7_clock = clock; // @[:@44728.4]
  assign fifos_7_reset = reset; // @[:@44729.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@44755.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44757.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44761.4]
  assign fifos_8_clock = clock; // @[:@44763.4]
  assign fifos_8_reset = reset; // @[:@44764.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@44790.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44792.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44796.4]
  assign fifos_9_clock = clock; // @[:@44798.4]
  assign fifos_9_reset = reset; // @[:@44799.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@44825.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44827.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44831.4]
  assign fifos_10_clock = clock; // @[:@44833.4]
  assign fifos_10_reset = reset; // @[:@44834.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@44860.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44862.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44866.4]
  assign fifos_11_clock = clock; // @[:@44868.4]
  assign fifos_11_reset = reset; // @[:@44869.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@44895.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44897.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44901.4]
  assign fifos_12_clock = clock; // @[:@44903.4]
  assign fifos_12_reset = reset; // @[:@44904.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@44930.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44932.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44936.4]
  assign fifos_13_clock = clock; // @[:@44938.4]
  assign fifos_13_reset = reset; // @[:@44939.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@44965.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@44967.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@44971.4]
  assign fifos_14_clock = clock; // @[:@44973.4]
  assign fifos_14_reset = reset; // @[:@44974.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@45000.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@45002.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@45006.4]
  assign fifos_15_clock = clock; // @[:@45008.4]
  assign fifos_15_reset = reset; // @[:@45009.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@45035.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@45037.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@45041.4]
endmodule
module FFRAM( // @[:@45506.2]
  input        clock, // @[:@45507.4]
  input        reset, // @[:@45508.4]
  input  [1:0] io_raddr, // @[:@45509.4]
  input        io_wen, // @[:@45509.4]
  input  [1:0] io_waddr, // @[:@45509.4]
  input        io_wdata, // @[:@45509.4]
  output       io_rdata, // @[:@45509.4]
  input        io_banks_0_wdata_valid, // @[:@45509.4]
  input        io_banks_0_wdata_bits, // @[:@45509.4]
  input        io_banks_1_wdata_valid, // @[:@45509.4]
  input        io_banks_1_wdata_bits, // @[:@45509.4]
  input        io_banks_2_wdata_valid, // @[:@45509.4]
  input        io_banks_2_wdata_bits, // @[:@45509.4]
  input        io_banks_3_wdata_valid, // @[:@45509.4]
  input        io_banks_3_wdata_bits // @[:@45509.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@45513.4]
  reg [31:0] _RAND_0;
  wire  _T_88; // @[SRAM.scala 148:37:@45514.4]
  wire  _T_89; // @[SRAM.scala 148:25:@45515.4]
  wire  _T_90; // @[SRAM.scala 148:15:@45516.4]
  wire  _T_91; // @[SRAM.scala 149:15:@45518.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@45517.4]
  reg  regs_1; // @[SRAM.scala 145:20:@45524.4]
  reg [31:0] _RAND_1;
  wire  _T_97; // @[SRAM.scala 148:37:@45525.4]
  wire  _T_98; // @[SRAM.scala 148:25:@45526.4]
  wire  _T_99; // @[SRAM.scala 148:15:@45527.4]
  wire  _T_100; // @[SRAM.scala 149:15:@45529.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@45528.4]
  reg  regs_2; // @[SRAM.scala 145:20:@45535.4]
  reg [31:0] _RAND_2;
  wire  _T_106; // @[SRAM.scala 148:37:@45536.4]
  wire  _T_107; // @[SRAM.scala 148:25:@45537.4]
  wire  _T_108; // @[SRAM.scala 148:15:@45538.4]
  wire  _T_109; // @[SRAM.scala 149:15:@45540.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@45539.4]
  reg  regs_3; // @[SRAM.scala 145:20:@45546.4]
  reg [31:0] _RAND_3;
  wire  _T_115; // @[SRAM.scala 148:37:@45547.4]
  wire  _T_116; // @[SRAM.scala 148:25:@45548.4]
  wire  _T_117; // @[SRAM.scala 148:15:@45549.4]
  wire  _T_118; // @[SRAM.scala 149:15:@45551.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@45550.4]
  wire  _GEN_5; // @[SRAM.scala 155:12:@45560.4]
  wire  _GEN_6; // @[SRAM.scala 155:12:@45560.4]
  assign _T_88 = io_waddr == 2'h0; // @[SRAM.scala 148:37:@45514.4]
  assign _T_89 = io_wen & _T_88; // @[SRAM.scala 148:25:@45515.4]
  assign _T_90 = io_banks_0_wdata_valid | _T_89; // @[SRAM.scala 148:15:@45516.4]
  assign _T_91 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45518.6]
  assign _GEN_0 = _T_90 ? _T_91 : regs_0; // @[SRAM.scala 148:48:@45517.4]
  assign _T_97 = io_waddr == 2'h1; // @[SRAM.scala 148:37:@45525.4]
  assign _T_98 = io_wen & _T_97; // @[SRAM.scala 148:25:@45526.4]
  assign _T_99 = io_banks_1_wdata_valid | _T_98; // @[SRAM.scala 148:15:@45527.4]
  assign _T_100 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45529.6]
  assign _GEN_1 = _T_99 ? _T_100 : regs_1; // @[SRAM.scala 148:48:@45528.4]
  assign _T_106 = io_waddr == 2'h2; // @[SRAM.scala 148:37:@45536.4]
  assign _T_107 = io_wen & _T_106; // @[SRAM.scala 148:25:@45537.4]
  assign _T_108 = io_banks_2_wdata_valid | _T_107; // @[SRAM.scala 148:15:@45538.4]
  assign _T_109 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45540.6]
  assign _GEN_2 = _T_108 ? _T_109 : regs_2; // @[SRAM.scala 148:48:@45539.4]
  assign _T_115 = io_waddr == 2'h3; // @[SRAM.scala 148:37:@45547.4]
  assign _T_116 = io_wen & _T_115; // @[SRAM.scala 148:25:@45548.4]
  assign _T_117 = io_banks_3_wdata_valid | _T_116; // @[SRAM.scala 148:15:@45549.4]
  assign _T_118 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@45551.6]
  assign _GEN_3 = _T_117 ? _T_118 : regs_3; // @[SRAM.scala 148:48:@45550.4]
  assign _GEN_5 = 2'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@45560.4]
  assign _GEN_6 = 2'h2 == io_raddr ? regs_2 : _GEN_5; // @[SRAM.scala 155:12:@45560.4]
  assign io_rdata = 2'h3 == io_raddr ? regs_3 : _GEN_6; // @[SRAM.scala 155:12:@45560.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_90) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_99) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_108) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_117) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_17( // @[:@45562.2]
  input   clock, // @[:@45563.4]
  input   reset, // @[:@45564.4]
  output  io_in_ready, // @[:@45565.4]
  input   io_in_valid, // @[:@45565.4]
  input   io_in_bits, // @[:@45565.4]
  input   io_out_ready, // @[:@45565.4]
  output  io_out_valid, // @[:@45565.4]
  output  io_out_bits // @[:@45565.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@45591.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@45591.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@45591.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@45591.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@45591.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@45591.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@45591.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@45601.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@45601.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@45601.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@45601.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@45601.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@45601.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@45601.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@45616.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@45616.4]
  wire [1:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@45616.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@45616.4]
  wire [1:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@45616.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@45616.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@45616.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@45616.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@45616.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@45616.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@45616.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@45616.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@45616.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@45616.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@45616.4]
  wire  writeEn; // @[FIFO.scala 30:29:@45589.4]
  wire  readEn; // @[FIFO.scala 31:29:@45590.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@45611.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@45612.4]
  wire  _T_104; // @[FIFO.scala 45:27:@45613.4]
  wire  empty; // @[FIFO.scala 45:24:@45614.4]
  wire  full; // @[FIFO.scala 46:23:@45615.4]
  wire  _T_157; // @[FIFO.scala 83:17:@45702.4]
  wire  _GEN_4; // @[FIFO.scala 83:29:@45703.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@45591.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@45601.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM FFRAM ( // @[FIFO.scala 49:19:@45616.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@45589.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@45590.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@45612.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@45613.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@45614.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@45615.4]
  assign _T_157 = writeEn != readEn; // @[FIFO.scala 83:17:@45702.4]
  assign _GEN_4 = _T_157 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@45703.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@45709.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@45707.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@45641.4]
  assign enqCounter_clock = clock; // @[:@45592.4]
  assign enqCounter_reset = reset; // @[:@45593.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@45599.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@45600.4]
  assign deqCounter_clock = clock; // @[:@45602.4]
  assign deqCounter_reset = reset; // @[:@45603.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@45609.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@45610.4]
  assign FFRAM_clock = clock; // @[:@45617.4]
  assign FFRAM_reset = reset; // @[:@45618.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@45637.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@45638.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@45639.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@45640.4]
  assign FFRAM_io_banks_0_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@45643.4]
  assign FFRAM_io_banks_0_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@45642.4]
  assign FFRAM_io_banks_1_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@45646.4]
  assign FFRAM_io_banks_1_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@45645.4]
  assign FFRAM_io_banks_2_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@45649.4]
  assign FFRAM_io_banks_2_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@45648.4]
  assign FFRAM_io_banks_3_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@45652.4]
  assign FFRAM_io_banks_3_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@45651.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_157) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec_1( // @[:@49326.2]
  input   clock, // @[:@49327.4]
  input   reset, // @[:@49328.4]
  output  io_in_ready, // @[:@49329.4]
  input   io_in_valid, // @[:@49329.4]
  input   io_in_bits_0, // @[:@49329.4]
  input   io_out_ready, // @[:@49329.4]
  output  io_out_valid, // @[:@49329.4]
  output  io_out_bits_0, // @[:@49329.4]
  output  io_out_bits_1, // @[:@49329.4]
  output  io_out_bits_2, // @[:@49329.4]
  output  io_out_bits_3, // @[:@49329.4]
  output  io_out_bits_4, // @[:@49329.4]
  output  io_out_bits_5, // @[:@49329.4]
  output  io_out_bits_6, // @[:@49329.4]
  output  io_out_bits_7, // @[:@49329.4]
  output  io_out_bits_8, // @[:@49329.4]
  output  io_out_bits_9, // @[:@49329.4]
  output  io_out_bits_10, // @[:@49329.4]
  output  io_out_bits_11, // @[:@49329.4]
  output  io_out_bits_12, // @[:@49329.4]
  output  io_out_bits_13, // @[:@49329.4]
  output  io_out_bits_14, // @[:@49329.4]
  output  io_out_bits_15 // @[:@49329.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@49333.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@49333.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@49333.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@49333.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@49344.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@49344.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@49344.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@49344.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@49357.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@49357.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@49357.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@49357.4]
  wire  fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@49357.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@49357.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@49357.4]
  wire  fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@49357.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@49392.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@49392.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@49392.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@49392.4]
  wire  fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@49392.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@49392.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@49392.4]
  wire  fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@49392.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@49427.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@49427.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@49427.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@49427.4]
  wire  fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@49427.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@49427.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@49427.4]
  wire  fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@49427.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@49462.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@49462.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@49462.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@49462.4]
  wire  fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@49462.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@49462.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@49462.4]
  wire  fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@49462.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@49497.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@49497.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@49497.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@49497.4]
  wire  fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@49497.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@49497.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@49497.4]
  wire  fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@49497.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@49532.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@49532.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@49532.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@49532.4]
  wire  fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@49532.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@49532.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@49532.4]
  wire  fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@49532.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@49567.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@49567.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@49567.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@49567.4]
  wire  fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@49567.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@49567.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@49567.4]
  wire  fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@49567.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@49602.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@49602.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@49602.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@49602.4]
  wire  fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@49602.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@49602.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@49602.4]
  wire  fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@49602.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@49637.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@49637.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@49637.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@49637.4]
  wire  fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@49637.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@49637.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@49637.4]
  wire  fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@49637.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@49672.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@49672.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@49672.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@49672.4]
  wire  fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@49672.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@49672.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@49672.4]
  wire  fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@49672.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@49707.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@49707.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@49707.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@49707.4]
  wire  fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@49707.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@49707.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@49707.4]
  wire  fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@49707.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@49742.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@49742.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@49742.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@49742.4]
  wire  fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@49742.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@49742.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@49742.4]
  wire  fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@49742.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@49777.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@49777.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@49777.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@49777.4]
  wire  fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@49777.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@49777.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@49777.4]
  wire  fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@49777.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@49812.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@49812.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@49812.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@49812.4]
  wire  fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@49812.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@49812.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@49812.4]
  wire  fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@49812.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@49847.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@49847.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@49847.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@49847.4]
  wire  fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@49847.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@49847.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@49847.4]
  wire  fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@49847.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@49882.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@49882.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@49882.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@49882.4]
  wire  fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@49882.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@49882.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@49882.4]
  wire  fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@49882.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@49332.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@49355.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@49382.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@49417.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@49452.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@49487.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@49522.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@49557.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@49592.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@49627.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@49662.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@49697.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@49732.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@49767.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@49802.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@49837.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@49872.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@49907.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49918.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49919.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@49949.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49920.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@49949.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49921.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@49949.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49922.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@49949.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49923.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@49949.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49924.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@49949.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49925.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@49949.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49926.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@49949.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49927.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@49949.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49928.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@49949.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49929.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@49949.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49930.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@49949.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49931.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@49949.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49932.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@49949.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49933.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@49968.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@49969.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@49970.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@49971.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@49972.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@49973.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@49974.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@49975.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@49976.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@49977.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@49978.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@49979.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@49980.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@49981.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@49333.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@49344.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_17 fifos_0 ( // @[FIFOVec.scala 40:19:@49357.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_17 fifos_1 ( // @[FIFOVec.scala 40:19:@49392.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_17 fifos_2 ( // @[FIFOVec.scala 40:19:@49427.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_17 fifos_3 ( // @[FIFOVec.scala 40:19:@49462.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_17 fifos_4 ( // @[FIFOVec.scala 40:19:@49497.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_17 fifos_5 ( // @[FIFOVec.scala 40:19:@49532.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_17 fifos_6 ( // @[FIFOVec.scala 40:19:@49567.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_17 fifos_7 ( // @[FIFOVec.scala 40:19:@49602.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_17 fifos_8 ( // @[FIFOVec.scala 40:19:@49637.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_17 fifos_9 ( // @[FIFOVec.scala 40:19:@49672.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_17 fifos_10 ( // @[FIFOVec.scala 40:19:@49707.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_17 fifos_11 ( // @[FIFOVec.scala 40:19:@49742.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_17 fifos_12 ( // @[FIFOVec.scala 40:19:@49777.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_17 fifos_13 ( // @[FIFOVec.scala 40:19:@49812.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_17 fifos_14 ( // @[FIFOVec.scala 40:19:@49847.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_17 fifos_15 ( // @[FIFOVec.scala 40:19:@49882.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@49332.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@49355.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@49382.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@49417.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@49452.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@49487.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@49522.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@49557.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@49592.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@49627.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@49662.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@49697.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@49732.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@49767.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@49802.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@49837.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@49872.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@49907.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49918.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49919.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@49949.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49920.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@49949.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49921.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@49949.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49922.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@49949.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49923.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@49949.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49924.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@49949.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49925.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@49949.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49926.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@49949.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49927.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@49949.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49928.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@49949.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49929.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@49949.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49930.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@49949.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49931.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@49949.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49932.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@49949.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@49917.4 FIFOVec.scala 49:42:@49933.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@49968.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@49969.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@49970.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@49971.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@49972.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@49973.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@49974.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@49975.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@49976.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@49977.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@49978.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@49979.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@49980.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@49981.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@49950.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@49984.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@50292.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@50293.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@50294.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@50295.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@50296.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@50297.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@50298.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@50299.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@50300.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@50301.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@50302.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@50303.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@50304.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@50305.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@50306.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@50307.4]
  assign enqCounter_clock = clock; // @[:@49334.4]
  assign enqCounter_reset = reset; // @[:@49335.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@49342.4]
  assign deqCounter_clock = clock; // @[:@49345.4]
  assign deqCounter_reset = reset; // @[:@49346.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@49353.4]
  assign fifos_0_clock = clock; // @[:@49358.4]
  assign fifos_0_reset = reset; // @[:@49359.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@49385.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49387.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49391.4]
  assign fifos_1_clock = clock; // @[:@49393.4]
  assign fifos_1_reset = reset; // @[:@49394.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@49420.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49422.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49426.4]
  assign fifos_2_clock = clock; // @[:@49428.4]
  assign fifos_2_reset = reset; // @[:@49429.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@49455.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49457.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49461.4]
  assign fifos_3_clock = clock; // @[:@49463.4]
  assign fifos_3_reset = reset; // @[:@49464.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@49490.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49492.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49496.4]
  assign fifos_4_clock = clock; // @[:@49498.4]
  assign fifos_4_reset = reset; // @[:@49499.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@49525.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49527.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49531.4]
  assign fifos_5_clock = clock; // @[:@49533.4]
  assign fifos_5_reset = reset; // @[:@49534.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@49560.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49562.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49566.4]
  assign fifos_6_clock = clock; // @[:@49568.4]
  assign fifos_6_reset = reset; // @[:@49569.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@49595.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49597.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49601.4]
  assign fifos_7_clock = clock; // @[:@49603.4]
  assign fifos_7_reset = reset; // @[:@49604.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@49630.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49632.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49636.4]
  assign fifos_8_clock = clock; // @[:@49638.4]
  assign fifos_8_reset = reset; // @[:@49639.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@49665.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49667.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49671.4]
  assign fifos_9_clock = clock; // @[:@49673.4]
  assign fifos_9_reset = reset; // @[:@49674.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@49700.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49702.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49706.4]
  assign fifos_10_clock = clock; // @[:@49708.4]
  assign fifos_10_reset = reset; // @[:@49709.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@49735.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49737.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49741.4]
  assign fifos_11_clock = clock; // @[:@49743.4]
  assign fifos_11_reset = reset; // @[:@49744.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@49770.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49772.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49776.4]
  assign fifos_12_clock = clock; // @[:@49778.4]
  assign fifos_12_reset = reset; // @[:@49779.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@49805.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49807.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49811.4]
  assign fifos_13_clock = clock; // @[:@49813.4]
  assign fifos_13_reset = reset; // @[:@49814.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@49840.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49842.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49846.4]
  assign fifos_14_clock = clock; // @[:@49848.4]
  assign fifos_14_reset = reset; // @[:@49849.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@49875.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49877.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49881.4]
  assign fifos_15_clock = clock; // @[:@49883.4]
  assign fifos_15_reset = reset; // @[:@49884.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@49910.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@49912.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@49916.4]
endmodule
module FIFOWidthConvert( // @[:@50309.2]
  input         clock, // @[:@50310.4]
  input         reset, // @[:@50311.4]
  output        io_in_ready, // @[:@50312.4]
  input         io_in_valid, // @[:@50312.4]
  input  [31:0] io_in_bits_data_0, // @[:@50312.4]
  input         io_in_bits_strobe, // @[:@50312.4]
  input         io_out_ready, // @[:@50312.4]
  output        io_out_valid, // @[:@50312.4]
  output [31:0] io_out_bits_data_0, // @[:@50312.4]
  output [31:0] io_out_bits_data_1, // @[:@50312.4]
  output [31:0] io_out_bits_data_2, // @[:@50312.4]
  output [31:0] io_out_bits_data_3, // @[:@50312.4]
  output [31:0] io_out_bits_data_4, // @[:@50312.4]
  output [31:0] io_out_bits_data_5, // @[:@50312.4]
  output [31:0] io_out_bits_data_6, // @[:@50312.4]
  output [31:0] io_out_bits_data_7, // @[:@50312.4]
  output [31:0] io_out_bits_data_8, // @[:@50312.4]
  output [31:0] io_out_bits_data_9, // @[:@50312.4]
  output [31:0] io_out_bits_data_10, // @[:@50312.4]
  output [31:0] io_out_bits_data_11, // @[:@50312.4]
  output [31:0] io_out_bits_data_12, // @[:@50312.4]
  output [31:0] io_out_bits_data_13, // @[:@50312.4]
  output [31:0] io_out_bits_data_14, // @[:@50312.4]
  output [31:0] io_out_bits_data_15, // @[:@50312.4]
  output [63:0] io_out_bits_strobe // @[:@50312.4]
);
  wire  FIFOVec_clock; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire  FIFOVec_reset; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire  FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire  FIFOVec_io_in_valid; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire [31:0] FIFOVec_io_in_bits_0; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire  FIFOVec_io_out_ready; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire  FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire [31:0] FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire [31:0] FIFOVec_io_out_bits_1; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire [31:0] FIFOVec_io_out_bits_2; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire [31:0] FIFOVec_io_out_bits_3; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire [31:0] FIFOVec_io_out_bits_4; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire [31:0] FIFOVec_io_out_bits_5; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire [31:0] FIFOVec_io_out_bits_6; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire [31:0] FIFOVec_io_out_bits_7; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire [31:0] FIFOVec_io_out_bits_8; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire [31:0] FIFOVec_io_out_bits_9; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire [31:0] FIFOVec_io_out_bits_10; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire [31:0] FIFOVec_io_out_bits_11; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire [31:0] FIFOVec_io_out_bits_12; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire [31:0] FIFOVec_io_out_bits_13; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire [31:0] FIFOVec_io_out_bits_14; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire [31:0] FIFOVec_io_out_bits_15; // @[FIFOWidthConvert.scala 61:22:@50314.4]
  wire  FIFOVec_1_clock; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_reset; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_in_ready; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_in_valid; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_in_bits_0; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_out_ready; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_out_valid; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_out_bits_0; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_out_bits_1; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_out_bits_2; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_out_bits_3; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_out_bits_4; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_out_bits_5; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_out_bits_6; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_out_bits_7; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_out_bits_8; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_out_bits_9; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_out_bits_10; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_out_bits_11; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_out_bits_12; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_out_bits_13; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_out_bits_14; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire  FIFOVec_1_io_out_bits_15; // @[FIFOWidthConvert.scala 62:26:@50355.4]
  wire [319:0] _T_55; // @[Cat.scala 30:58:@50414.4]
  wire [511:0] _T_61; // @[Cat.scala 30:58:@50420.4]
  wire [9:0] _T_108; // @[Cat.scala 30:58:@50478.4]
  wire [15:0] _T_114; // @[Cat.scala 30:58:@50484.4]
  wire  _T_115; // @[FIFOWidthConvert.scala 36:14:@50485.4]
  wire  _T_119; // @[FIFOWidthConvert.scala 36:14:@50489.4]
  wire  _T_123; // @[FIFOWidthConvert.scala 36:14:@50493.4]
  wire  _T_127; // @[FIFOWidthConvert.scala 36:14:@50497.4]
  wire  _T_131; // @[FIFOWidthConvert.scala 36:14:@50501.4]
  wire  _T_135; // @[FIFOWidthConvert.scala 36:14:@50505.4]
  wire  _T_139; // @[FIFOWidthConvert.scala 36:14:@50509.4]
  wire  _T_143; // @[FIFOWidthConvert.scala 36:14:@50513.4]
  wire  _T_147; // @[FIFOWidthConvert.scala 36:14:@50517.4]
  wire  _T_151; // @[FIFOWidthConvert.scala 36:14:@50521.4]
  wire  _T_155; // @[FIFOWidthConvert.scala 36:14:@50525.4]
  wire  _T_159; // @[FIFOWidthConvert.scala 36:14:@50529.4]
  wire  _T_163; // @[FIFOWidthConvert.scala 36:14:@50533.4]
  wire  _T_167; // @[FIFOWidthConvert.scala 36:14:@50537.4]
  wire  _T_171; // @[FIFOWidthConvert.scala 36:14:@50541.4]
  wire  _T_175; // @[FIFOWidthConvert.scala 36:14:@50545.4]
  wire [9:0] _T_257; // @[Cat.scala 30:58:@50622.4]
  wire [18:0] _T_266; // @[Cat.scala 30:58:@50631.4]
  wire [27:0] _T_275; // @[Cat.scala 30:58:@50640.4]
  wire [36:0] _T_284; // @[Cat.scala 30:58:@50649.4]
  wire [45:0] _T_293; // @[Cat.scala 30:58:@50658.4]
  wire [54:0] _T_302; // @[Cat.scala 30:58:@50667.4]
  wire [62:0] _T_310; // @[Cat.scala 30:58:@50675.4]
  FIFOVec FIFOVec ( // @[FIFOWidthConvert.scala 61:22:@50314.4]
    .clock(FIFOVec_clock),
    .reset(FIFOVec_reset),
    .io_in_ready(FIFOVec_io_in_ready),
    .io_in_valid(FIFOVec_io_in_valid),
    .io_in_bits_0(FIFOVec_io_in_bits_0),
    .io_out_ready(FIFOVec_io_out_ready),
    .io_out_valid(FIFOVec_io_out_valid),
    .io_out_bits_0(FIFOVec_io_out_bits_0),
    .io_out_bits_1(FIFOVec_io_out_bits_1),
    .io_out_bits_2(FIFOVec_io_out_bits_2),
    .io_out_bits_3(FIFOVec_io_out_bits_3),
    .io_out_bits_4(FIFOVec_io_out_bits_4),
    .io_out_bits_5(FIFOVec_io_out_bits_5),
    .io_out_bits_6(FIFOVec_io_out_bits_6),
    .io_out_bits_7(FIFOVec_io_out_bits_7),
    .io_out_bits_8(FIFOVec_io_out_bits_8),
    .io_out_bits_9(FIFOVec_io_out_bits_9),
    .io_out_bits_10(FIFOVec_io_out_bits_10),
    .io_out_bits_11(FIFOVec_io_out_bits_11),
    .io_out_bits_12(FIFOVec_io_out_bits_12),
    .io_out_bits_13(FIFOVec_io_out_bits_13),
    .io_out_bits_14(FIFOVec_io_out_bits_14),
    .io_out_bits_15(FIFOVec_io_out_bits_15)
  );
  FIFOVec_1 FIFOVec_1 ( // @[FIFOWidthConvert.scala 62:26:@50355.4]
    .clock(FIFOVec_1_clock),
    .reset(FIFOVec_1_reset),
    .io_in_ready(FIFOVec_1_io_in_ready),
    .io_in_valid(FIFOVec_1_io_in_valid),
    .io_in_bits_0(FIFOVec_1_io_in_bits_0),
    .io_out_ready(FIFOVec_1_io_out_ready),
    .io_out_valid(FIFOVec_1_io_out_valid),
    .io_out_bits_0(FIFOVec_1_io_out_bits_0),
    .io_out_bits_1(FIFOVec_1_io_out_bits_1),
    .io_out_bits_2(FIFOVec_1_io_out_bits_2),
    .io_out_bits_3(FIFOVec_1_io_out_bits_3),
    .io_out_bits_4(FIFOVec_1_io_out_bits_4),
    .io_out_bits_5(FIFOVec_1_io_out_bits_5),
    .io_out_bits_6(FIFOVec_1_io_out_bits_6),
    .io_out_bits_7(FIFOVec_1_io_out_bits_7),
    .io_out_bits_8(FIFOVec_1_io_out_bits_8),
    .io_out_bits_9(FIFOVec_1_io_out_bits_9),
    .io_out_bits_10(FIFOVec_1_io_out_bits_10),
    .io_out_bits_11(FIFOVec_1_io_out_bits_11),
    .io_out_bits_12(FIFOVec_1_io_out_bits_12),
    .io_out_bits_13(FIFOVec_1_io_out_bits_13),
    .io_out_bits_14(FIFOVec_1_io_out_bits_14),
    .io_out_bits_15(FIFOVec_1_io_out_bits_15)
  );
  assign _T_55 = {FIFOVec_io_out_bits_15,FIFOVec_io_out_bits_14,FIFOVec_io_out_bits_13,FIFOVec_io_out_bits_12,FIFOVec_io_out_bits_11,FIFOVec_io_out_bits_10,FIFOVec_io_out_bits_9,FIFOVec_io_out_bits_8,FIFOVec_io_out_bits_7,FIFOVec_io_out_bits_6}; // @[Cat.scala 30:58:@50414.4]
  assign _T_61 = {_T_55,FIFOVec_io_out_bits_5,FIFOVec_io_out_bits_4,FIFOVec_io_out_bits_3,FIFOVec_io_out_bits_2,FIFOVec_io_out_bits_1,FIFOVec_io_out_bits_0}; // @[Cat.scala 30:58:@50420.4]
  assign _T_108 = {FIFOVec_1_io_out_bits_0,FIFOVec_1_io_out_bits_1,FIFOVec_1_io_out_bits_2,FIFOVec_1_io_out_bits_3,FIFOVec_1_io_out_bits_4,FIFOVec_1_io_out_bits_5,FIFOVec_1_io_out_bits_6,FIFOVec_1_io_out_bits_7,FIFOVec_1_io_out_bits_8,FIFOVec_1_io_out_bits_9}; // @[Cat.scala 30:58:@50478.4]
  assign _T_114 = {_T_108,FIFOVec_1_io_out_bits_10,FIFOVec_1_io_out_bits_11,FIFOVec_1_io_out_bits_12,FIFOVec_1_io_out_bits_13,FIFOVec_1_io_out_bits_14,FIFOVec_1_io_out_bits_15}; // @[Cat.scala 30:58:@50484.4]
  assign _T_115 = _T_114[0]; // @[FIFOWidthConvert.scala 36:14:@50485.4]
  assign _T_119 = _T_114[1]; // @[FIFOWidthConvert.scala 36:14:@50489.4]
  assign _T_123 = _T_114[2]; // @[FIFOWidthConvert.scala 36:14:@50493.4]
  assign _T_127 = _T_114[3]; // @[FIFOWidthConvert.scala 36:14:@50497.4]
  assign _T_131 = _T_114[4]; // @[FIFOWidthConvert.scala 36:14:@50501.4]
  assign _T_135 = _T_114[5]; // @[FIFOWidthConvert.scala 36:14:@50505.4]
  assign _T_139 = _T_114[6]; // @[FIFOWidthConvert.scala 36:14:@50509.4]
  assign _T_143 = _T_114[7]; // @[FIFOWidthConvert.scala 36:14:@50513.4]
  assign _T_147 = _T_114[8]; // @[FIFOWidthConvert.scala 36:14:@50517.4]
  assign _T_151 = _T_114[9]; // @[FIFOWidthConvert.scala 36:14:@50521.4]
  assign _T_155 = _T_114[10]; // @[FIFOWidthConvert.scala 36:14:@50525.4]
  assign _T_159 = _T_114[11]; // @[FIFOWidthConvert.scala 36:14:@50529.4]
  assign _T_163 = _T_114[12]; // @[FIFOWidthConvert.scala 36:14:@50533.4]
  assign _T_167 = _T_114[13]; // @[FIFOWidthConvert.scala 36:14:@50537.4]
  assign _T_171 = _T_114[14]; // @[FIFOWidthConvert.scala 36:14:@50541.4]
  assign _T_175 = _T_114[15]; // @[FIFOWidthConvert.scala 36:14:@50545.4]
  assign _T_257 = {_T_175,_T_175,_T_175,_T_175,_T_171,_T_171,_T_171,_T_171,_T_167,_T_167}; // @[Cat.scala 30:58:@50622.4]
  assign _T_266 = {_T_257,_T_167,_T_167,_T_163,_T_163,_T_163,_T_163,_T_159,_T_159,_T_159}; // @[Cat.scala 30:58:@50631.4]
  assign _T_275 = {_T_266,_T_159,_T_155,_T_155,_T_155,_T_155,_T_151,_T_151,_T_151,_T_151}; // @[Cat.scala 30:58:@50640.4]
  assign _T_284 = {_T_275,_T_147,_T_147,_T_147,_T_147,_T_143,_T_143,_T_143,_T_143,_T_139}; // @[Cat.scala 30:58:@50649.4]
  assign _T_293 = {_T_284,_T_139,_T_139,_T_139,_T_135,_T_135,_T_135,_T_135,_T_131,_T_131}; // @[Cat.scala 30:58:@50658.4]
  assign _T_302 = {_T_293,_T_131,_T_131,_T_127,_T_127,_T_127,_T_127,_T_123,_T_123,_T_123}; // @[Cat.scala 30:58:@50667.4]
  assign _T_310 = {_T_302,_T_123,_T_119,_T_119,_T_119,_T_119,_T_115,_T_115,_T_115}; // @[Cat.scala 30:58:@50675.4]
  assign io_in_ready = FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 71:17:@50404.4]
  assign io_out_valid = FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 72:18:@50405.4]
  assign io_out_bits_data_0 = _T_61[31:0]; // @[FIFOWidthConvert.scala 73:22:@50454.4]
  assign io_out_bits_data_1 = _T_61[63:32]; // @[FIFOWidthConvert.scala 73:22:@50455.4]
  assign io_out_bits_data_2 = _T_61[95:64]; // @[FIFOWidthConvert.scala 73:22:@50456.4]
  assign io_out_bits_data_3 = _T_61[127:96]; // @[FIFOWidthConvert.scala 73:22:@50457.4]
  assign io_out_bits_data_4 = _T_61[159:128]; // @[FIFOWidthConvert.scala 73:22:@50458.4]
  assign io_out_bits_data_5 = _T_61[191:160]; // @[FIFOWidthConvert.scala 73:22:@50459.4]
  assign io_out_bits_data_6 = _T_61[223:192]; // @[FIFOWidthConvert.scala 73:22:@50460.4]
  assign io_out_bits_data_7 = _T_61[255:224]; // @[FIFOWidthConvert.scala 73:22:@50461.4]
  assign io_out_bits_data_8 = _T_61[287:256]; // @[FIFOWidthConvert.scala 73:22:@50462.4]
  assign io_out_bits_data_9 = _T_61[319:288]; // @[FIFOWidthConvert.scala 73:22:@50463.4]
  assign io_out_bits_data_10 = _T_61[351:320]; // @[FIFOWidthConvert.scala 73:22:@50464.4]
  assign io_out_bits_data_11 = _T_61[383:352]; // @[FIFOWidthConvert.scala 73:22:@50465.4]
  assign io_out_bits_data_12 = _T_61[415:384]; // @[FIFOWidthConvert.scala 73:22:@50466.4]
  assign io_out_bits_data_13 = _T_61[447:416]; // @[FIFOWidthConvert.scala 73:22:@50467.4]
  assign io_out_bits_data_14 = _T_61[479:448]; // @[FIFOWidthConvert.scala 73:22:@50468.4]
  assign io_out_bits_data_15 = _T_61[511:480]; // @[FIFOWidthConvert.scala 73:22:@50469.4]
  assign io_out_bits_strobe = {_T_310,_T_115}; // @[FIFOWidthConvert.scala 74:24:@50677.4]
  assign FIFOVec_clock = clock; // @[:@50315.4]
  assign FIFOVec_reset = reset; // @[:@50316.4]
  assign FIFOVec_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 68:22:@50401.4]
  assign FIFOVec_io_in_bits_0 = io_in_bits_data_0; // @[FIFOWidthConvert.scala 67:24:@50400.4]
  assign FIFOVec_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 75:23:@50678.4]
  assign FIFOVec_1_clock = clock; // @[:@50356.4]
  assign FIFOVec_1_reset = reset; // @[:@50357.4]
  assign FIFOVec_1_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 70:26:@50403.4]
  assign FIFOVec_1_io_in_bits_0 = io_in_bits_strobe; // @[FIFOWidthConvert.scala 69:28:@50402.4]
  assign FIFOVec_1_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 76:27:@50679.4]
endmodule
module FFRAM_16( // @[:@50717.2]
  input        clock, // @[:@50718.4]
  input        reset, // @[:@50719.4]
  input  [5:0] io_raddr, // @[:@50720.4]
  input        io_wen, // @[:@50720.4]
  input  [5:0] io_waddr, // @[:@50720.4]
  input        io_wdata, // @[:@50720.4]
  output       io_rdata, // @[:@50720.4]
  input        io_banks_0_wdata_valid, // @[:@50720.4]
  input        io_banks_0_wdata_bits, // @[:@50720.4]
  input        io_banks_1_wdata_valid, // @[:@50720.4]
  input        io_banks_1_wdata_bits, // @[:@50720.4]
  input        io_banks_2_wdata_valid, // @[:@50720.4]
  input        io_banks_2_wdata_bits, // @[:@50720.4]
  input        io_banks_3_wdata_valid, // @[:@50720.4]
  input        io_banks_3_wdata_bits, // @[:@50720.4]
  input        io_banks_4_wdata_valid, // @[:@50720.4]
  input        io_banks_4_wdata_bits, // @[:@50720.4]
  input        io_banks_5_wdata_valid, // @[:@50720.4]
  input        io_banks_5_wdata_bits, // @[:@50720.4]
  input        io_banks_6_wdata_valid, // @[:@50720.4]
  input        io_banks_6_wdata_bits, // @[:@50720.4]
  input        io_banks_7_wdata_valid, // @[:@50720.4]
  input        io_banks_7_wdata_bits, // @[:@50720.4]
  input        io_banks_8_wdata_valid, // @[:@50720.4]
  input        io_banks_8_wdata_bits, // @[:@50720.4]
  input        io_banks_9_wdata_valid, // @[:@50720.4]
  input        io_banks_9_wdata_bits, // @[:@50720.4]
  input        io_banks_10_wdata_valid, // @[:@50720.4]
  input        io_banks_10_wdata_bits, // @[:@50720.4]
  input        io_banks_11_wdata_valid, // @[:@50720.4]
  input        io_banks_11_wdata_bits, // @[:@50720.4]
  input        io_banks_12_wdata_valid, // @[:@50720.4]
  input        io_banks_12_wdata_bits, // @[:@50720.4]
  input        io_banks_13_wdata_valid, // @[:@50720.4]
  input        io_banks_13_wdata_bits, // @[:@50720.4]
  input        io_banks_14_wdata_valid, // @[:@50720.4]
  input        io_banks_14_wdata_bits, // @[:@50720.4]
  input        io_banks_15_wdata_valid, // @[:@50720.4]
  input        io_banks_15_wdata_bits, // @[:@50720.4]
  input        io_banks_16_wdata_valid, // @[:@50720.4]
  input        io_banks_16_wdata_bits, // @[:@50720.4]
  input        io_banks_17_wdata_valid, // @[:@50720.4]
  input        io_banks_17_wdata_bits, // @[:@50720.4]
  input        io_banks_18_wdata_valid, // @[:@50720.4]
  input        io_banks_18_wdata_bits, // @[:@50720.4]
  input        io_banks_19_wdata_valid, // @[:@50720.4]
  input        io_banks_19_wdata_bits, // @[:@50720.4]
  input        io_banks_20_wdata_valid, // @[:@50720.4]
  input        io_banks_20_wdata_bits, // @[:@50720.4]
  input        io_banks_21_wdata_valid, // @[:@50720.4]
  input        io_banks_21_wdata_bits, // @[:@50720.4]
  input        io_banks_22_wdata_valid, // @[:@50720.4]
  input        io_banks_22_wdata_bits, // @[:@50720.4]
  input        io_banks_23_wdata_valid, // @[:@50720.4]
  input        io_banks_23_wdata_bits, // @[:@50720.4]
  input        io_banks_24_wdata_valid, // @[:@50720.4]
  input        io_banks_24_wdata_bits, // @[:@50720.4]
  input        io_banks_25_wdata_valid, // @[:@50720.4]
  input        io_banks_25_wdata_bits, // @[:@50720.4]
  input        io_banks_26_wdata_valid, // @[:@50720.4]
  input        io_banks_26_wdata_bits, // @[:@50720.4]
  input        io_banks_27_wdata_valid, // @[:@50720.4]
  input        io_banks_27_wdata_bits, // @[:@50720.4]
  input        io_banks_28_wdata_valid, // @[:@50720.4]
  input        io_banks_28_wdata_bits, // @[:@50720.4]
  input        io_banks_29_wdata_valid, // @[:@50720.4]
  input        io_banks_29_wdata_bits, // @[:@50720.4]
  input        io_banks_30_wdata_valid, // @[:@50720.4]
  input        io_banks_30_wdata_bits, // @[:@50720.4]
  input        io_banks_31_wdata_valid, // @[:@50720.4]
  input        io_banks_31_wdata_bits, // @[:@50720.4]
  input        io_banks_32_wdata_valid, // @[:@50720.4]
  input        io_banks_32_wdata_bits, // @[:@50720.4]
  input        io_banks_33_wdata_valid, // @[:@50720.4]
  input        io_banks_33_wdata_bits, // @[:@50720.4]
  input        io_banks_34_wdata_valid, // @[:@50720.4]
  input        io_banks_34_wdata_bits, // @[:@50720.4]
  input        io_banks_35_wdata_valid, // @[:@50720.4]
  input        io_banks_35_wdata_bits, // @[:@50720.4]
  input        io_banks_36_wdata_valid, // @[:@50720.4]
  input        io_banks_36_wdata_bits, // @[:@50720.4]
  input        io_banks_37_wdata_valid, // @[:@50720.4]
  input        io_banks_37_wdata_bits, // @[:@50720.4]
  input        io_banks_38_wdata_valid, // @[:@50720.4]
  input        io_banks_38_wdata_bits, // @[:@50720.4]
  input        io_banks_39_wdata_valid, // @[:@50720.4]
  input        io_banks_39_wdata_bits, // @[:@50720.4]
  input        io_banks_40_wdata_valid, // @[:@50720.4]
  input        io_banks_40_wdata_bits, // @[:@50720.4]
  input        io_banks_41_wdata_valid, // @[:@50720.4]
  input        io_banks_41_wdata_bits, // @[:@50720.4]
  input        io_banks_42_wdata_valid, // @[:@50720.4]
  input        io_banks_42_wdata_bits, // @[:@50720.4]
  input        io_banks_43_wdata_valid, // @[:@50720.4]
  input        io_banks_43_wdata_bits, // @[:@50720.4]
  input        io_banks_44_wdata_valid, // @[:@50720.4]
  input        io_banks_44_wdata_bits, // @[:@50720.4]
  input        io_banks_45_wdata_valid, // @[:@50720.4]
  input        io_banks_45_wdata_bits, // @[:@50720.4]
  input        io_banks_46_wdata_valid, // @[:@50720.4]
  input        io_banks_46_wdata_bits, // @[:@50720.4]
  input        io_banks_47_wdata_valid, // @[:@50720.4]
  input        io_banks_47_wdata_bits, // @[:@50720.4]
  input        io_banks_48_wdata_valid, // @[:@50720.4]
  input        io_banks_48_wdata_bits, // @[:@50720.4]
  input        io_banks_49_wdata_valid, // @[:@50720.4]
  input        io_banks_49_wdata_bits, // @[:@50720.4]
  input        io_banks_50_wdata_valid, // @[:@50720.4]
  input        io_banks_50_wdata_bits, // @[:@50720.4]
  input        io_banks_51_wdata_valid, // @[:@50720.4]
  input        io_banks_51_wdata_bits, // @[:@50720.4]
  input        io_banks_52_wdata_valid, // @[:@50720.4]
  input        io_banks_52_wdata_bits, // @[:@50720.4]
  input        io_banks_53_wdata_valid, // @[:@50720.4]
  input        io_banks_53_wdata_bits, // @[:@50720.4]
  input        io_banks_54_wdata_valid, // @[:@50720.4]
  input        io_banks_54_wdata_bits, // @[:@50720.4]
  input        io_banks_55_wdata_valid, // @[:@50720.4]
  input        io_banks_55_wdata_bits, // @[:@50720.4]
  input        io_banks_56_wdata_valid, // @[:@50720.4]
  input        io_banks_56_wdata_bits, // @[:@50720.4]
  input        io_banks_57_wdata_valid, // @[:@50720.4]
  input        io_banks_57_wdata_bits, // @[:@50720.4]
  input        io_banks_58_wdata_valid, // @[:@50720.4]
  input        io_banks_58_wdata_bits, // @[:@50720.4]
  input        io_banks_59_wdata_valid, // @[:@50720.4]
  input        io_banks_59_wdata_bits, // @[:@50720.4]
  input        io_banks_60_wdata_valid, // @[:@50720.4]
  input        io_banks_60_wdata_bits, // @[:@50720.4]
  input        io_banks_61_wdata_valid, // @[:@50720.4]
  input        io_banks_61_wdata_bits, // @[:@50720.4]
  input        io_banks_62_wdata_valid, // @[:@50720.4]
  input        io_banks_62_wdata_bits, // @[:@50720.4]
  input        io_banks_63_wdata_valid, // @[:@50720.4]
  input        io_banks_63_wdata_bits // @[:@50720.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@50724.4]
  reg [31:0] _RAND_0;
  wire  _T_688; // @[SRAM.scala 148:37:@50725.4]
  wire  _T_689; // @[SRAM.scala 148:25:@50726.4]
  wire  _T_690; // @[SRAM.scala 148:15:@50727.4]
  wire  _T_691; // @[SRAM.scala 149:15:@50729.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@50728.4]
  reg  regs_1; // @[SRAM.scala 145:20:@50735.4]
  reg [31:0] _RAND_1;
  wire  _T_697; // @[SRAM.scala 148:37:@50736.4]
  wire  _T_698; // @[SRAM.scala 148:25:@50737.4]
  wire  _T_699; // @[SRAM.scala 148:15:@50738.4]
  wire  _T_700; // @[SRAM.scala 149:15:@50740.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@50739.4]
  reg  regs_2; // @[SRAM.scala 145:20:@50746.4]
  reg [31:0] _RAND_2;
  wire  _T_706; // @[SRAM.scala 148:37:@50747.4]
  wire  _T_707; // @[SRAM.scala 148:25:@50748.4]
  wire  _T_708; // @[SRAM.scala 148:15:@50749.4]
  wire  _T_709; // @[SRAM.scala 149:15:@50751.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@50750.4]
  reg  regs_3; // @[SRAM.scala 145:20:@50757.4]
  reg [31:0] _RAND_3;
  wire  _T_715; // @[SRAM.scala 148:37:@50758.4]
  wire  _T_716; // @[SRAM.scala 148:25:@50759.4]
  wire  _T_717; // @[SRAM.scala 148:15:@50760.4]
  wire  _T_718; // @[SRAM.scala 149:15:@50762.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@50761.4]
  reg  regs_4; // @[SRAM.scala 145:20:@50768.4]
  reg [31:0] _RAND_4;
  wire  _T_724; // @[SRAM.scala 148:37:@50769.4]
  wire  _T_725; // @[SRAM.scala 148:25:@50770.4]
  wire  _T_726; // @[SRAM.scala 148:15:@50771.4]
  wire  _T_727; // @[SRAM.scala 149:15:@50773.6]
  wire  _GEN_4; // @[SRAM.scala 148:48:@50772.4]
  reg  regs_5; // @[SRAM.scala 145:20:@50779.4]
  reg [31:0] _RAND_5;
  wire  _T_733; // @[SRAM.scala 148:37:@50780.4]
  wire  _T_734; // @[SRAM.scala 148:25:@50781.4]
  wire  _T_735; // @[SRAM.scala 148:15:@50782.4]
  wire  _T_736; // @[SRAM.scala 149:15:@50784.6]
  wire  _GEN_5; // @[SRAM.scala 148:48:@50783.4]
  reg  regs_6; // @[SRAM.scala 145:20:@50790.4]
  reg [31:0] _RAND_6;
  wire  _T_742; // @[SRAM.scala 148:37:@50791.4]
  wire  _T_743; // @[SRAM.scala 148:25:@50792.4]
  wire  _T_744; // @[SRAM.scala 148:15:@50793.4]
  wire  _T_745; // @[SRAM.scala 149:15:@50795.6]
  wire  _GEN_6; // @[SRAM.scala 148:48:@50794.4]
  reg  regs_7; // @[SRAM.scala 145:20:@50801.4]
  reg [31:0] _RAND_7;
  wire  _T_751; // @[SRAM.scala 148:37:@50802.4]
  wire  _T_752; // @[SRAM.scala 148:25:@50803.4]
  wire  _T_753; // @[SRAM.scala 148:15:@50804.4]
  wire  _T_754; // @[SRAM.scala 149:15:@50806.6]
  wire  _GEN_7; // @[SRAM.scala 148:48:@50805.4]
  reg  regs_8; // @[SRAM.scala 145:20:@50812.4]
  reg [31:0] _RAND_8;
  wire  _T_760; // @[SRAM.scala 148:37:@50813.4]
  wire  _T_761; // @[SRAM.scala 148:25:@50814.4]
  wire  _T_762; // @[SRAM.scala 148:15:@50815.4]
  wire  _T_763; // @[SRAM.scala 149:15:@50817.6]
  wire  _GEN_8; // @[SRAM.scala 148:48:@50816.4]
  reg  regs_9; // @[SRAM.scala 145:20:@50823.4]
  reg [31:0] _RAND_9;
  wire  _T_769; // @[SRAM.scala 148:37:@50824.4]
  wire  _T_770; // @[SRAM.scala 148:25:@50825.4]
  wire  _T_771; // @[SRAM.scala 148:15:@50826.4]
  wire  _T_772; // @[SRAM.scala 149:15:@50828.6]
  wire  _GEN_9; // @[SRAM.scala 148:48:@50827.4]
  reg  regs_10; // @[SRAM.scala 145:20:@50834.4]
  reg [31:0] _RAND_10;
  wire  _T_778; // @[SRAM.scala 148:37:@50835.4]
  wire  _T_779; // @[SRAM.scala 148:25:@50836.4]
  wire  _T_780; // @[SRAM.scala 148:15:@50837.4]
  wire  _T_781; // @[SRAM.scala 149:15:@50839.6]
  wire  _GEN_10; // @[SRAM.scala 148:48:@50838.4]
  reg  regs_11; // @[SRAM.scala 145:20:@50845.4]
  reg [31:0] _RAND_11;
  wire  _T_787; // @[SRAM.scala 148:37:@50846.4]
  wire  _T_788; // @[SRAM.scala 148:25:@50847.4]
  wire  _T_789; // @[SRAM.scala 148:15:@50848.4]
  wire  _T_790; // @[SRAM.scala 149:15:@50850.6]
  wire  _GEN_11; // @[SRAM.scala 148:48:@50849.4]
  reg  regs_12; // @[SRAM.scala 145:20:@50856.4]
  reg [31:0] _RAND_12;
  wire  _T_796; // @[SRAM.scala 148:37:@50857.4]
  wire  _T_797; // @[SRAM.scala 148:25:@50858.4]
  wire  _T_798; // @[SRAM.scala 148:15:@50859.4]
  wire  _T_799; // @[SRAM.scala 149:15:@50861.6]
  wire  _GEN_12; // @[SRAM.scala 148:48:@50860.4]
  reg  regs_13; // @[SRAM.scala 145:20:@50867.4]
  reg [31:0] _RAND_13;
  wire  _T_805; // @[SRAM.scala 148:37:@50868.4]
  wire  _T_806; // @[SRAM.scala 148:25:@50869.4]
  wire  _T_807; // @[SRAM.scala 148:15:@50870.4]
  wire  _T_808; // @[SRAM.scala 149:15:@50872.6]
  wire  _GEN_13; // @[SRAM.scala 148:48:@50871.4]
  reg  regs_14; // @[SRAM.scala 145:20:@50878.4]
  reg [31:0] _RAND_14;
  wire  _T_814; // @[SRAM.scala 148:37:@50879.4]
  wire  _T_815; // @[SRAM.scala 148:25:@50880.4]
  wire  _T_816; // @[SRAM.scala 148:15:@50881.4]
  wire  _T_817; // @[SRAM.scala 149:15:@50883.6]
  wire  _GEN_14; // @[SRAM.scala 148:48:@50882.4]
  reg  regs_15; // @[SRAM.scala 145:20:@50889.4]
  reg [31:0] _RAND_15;
  wire  _T_823; // @[SRAM.scala 148:37:@50890.4]
  wire  _T_824; // @[SRAM.scala 148:25:@50891.4]
  wire  _T_825; // @[SRAM.scala 148:15:@50892.4]
  wire  _T_826; // @[SRAM.scala 149:15:@50894.6]
  wire  _GEN_15; // @[SRAM.scala 148:48:@50893.4]
  reg  regs_16; // @[SRAM.scala 145:20:@50900.4]
  reg [31:0] _RAND_16;
  wire  _T_832; // @[SRAM.scala 148:37:@50901.4]
  wire  _T_833; // @[SRAM.scala 148:25:@50902.4]
  wire  _T_834; // @[SRAM.scala 148:15:@50903.4]
  wire  _T_835; // @[SRAM.scala 149:15:@50905.6]
  wire  _GEN_16; // @[SRAM.scala 148:48:@50904.4]
  reg  regs_17; // @[SRAM.scala 145:20:@50911.4]
  reg [31:0] _RAND_17;
  wire  _T_841; // @[SRAM.scala 148:37:@50912.4]
  wire  _T_842; // @[SRAM.scala 148:25:@50913.4]
  wire  _T_843; // @[SRAM.scala 148:15:@50914.4]
  wire  _T_844; // @[SRAM.scala 149:15:@50916.6]
  wire  _GEN_17; // @[SRAM.scala 148:48:@50915.4]
  reg  regs_18; // @[SRAM.scala 145:20:@50922.4]
  reg [31:0] _RAND_18;
  wire  _T_850; // @[SRAM.scala 148:37:@50923.4]
  wire  _T_851; // @[SRAM.scala 148:25:@50924.4]
  wire  _T_852; // @[SRAM.scala 148:15:@50925.4]
  wire  _T_853; // @[SRAM.scala 149:15:@50927.6]
  wire  _GEN_18; // @[SRAM.scala 148:48:@50926.4]
  reg  regs_19; // @[SRAM.scala 145:20:@50933.4]
  reg [31:0] _RAND_19;
  wire  _T_859; // @[SRAM.scala 148:37:@50934.4]
  wire  _T_860; // @[SRAM.scala 148:25:@50935.4]
  wire  _T_861; // @[SRAM.scala 148:15:@50936.4]
  wire  _T_862; // @[SRAM.scala 149:15:@50938.6]
  wire  _GEN_19; // @[SRAM.scala 148:48:@50937.4]
  reg  regs_20; // @[SRAM.scala 145:20:@50944.4]
  reg [31:0] _RAND_20;
  wire  _T_868; // @[SRAM.scala 148:37:@50945.4]
  wire  _T_869; // @[SRAM.scala 148:25:@50946.4]
  wire  _T_870; // @[SRAM.scala 148:15:@50947.4]
  wire  _T_871; // @[SRAM.scala 149:15:@50949.6]
  wire  _GEN_20; // @[SRAM.scala 148:48:@50948.4]
  reg  regs_21; // @[SRAM.scala 145:20:@50955.4]
  reg [31:0] _RAND_21;
  wire  _T_877; // @[SRAM.scala 148:37:@50956.4]
  wire  _T_878; // @[SRAM.scala 148:25:@50957.4]
  wire  _T_879; // @[SRAM.scala 148:15:@50958.4]
  wire  _T_880; // @[SRAM.scala 149:15:@50960.6]
  wire  _GEN_21; // @[SRAM.scala 148:48:@50959.4]
  reg  regs_22; // @[SRAM.scala 145:20:@50966.4]
  reg [31:0] _RAND_22;
  wire  _T_886; // @[SRAM.scala 148:37:@50967.4]
  wire  _T_887; // @[SRAM.scala 148:25:@50968.4]
  wire  _T_888; // @[SRAM.scala 148:15:@50969.4]
  wire  _T_889; // @[SRAM.scala 149:15:@50971.6]
  wire  _GEN_22; // @[SRAM.scala 148:48:@50970.4]
  reg  regs_23; // @[SRAM.scala 145:20:@50977.4]
  reg [31:0] _RAND_23;
  wire  _T_895; // @[SRAM.scala 148:37:@50978.4]
  wire  _T_896; // @[SRAM.scala 148:25:@50979.4]
  wire  _T_897; // @[SRAM.scala 148:15:@50980.4]
  wire  _T_898; // @[SRAM.scala 149:15:@50982.6]
  wire  _GEN_23; // @[SRAM.scala 148:48:@50981.4]
  reg  regs_24; // @[SRAM.scala 145:20:@50988.4]
  reg [31:0] _RAND_24;
  wire  _T_904; // @[SRAM.scala 148:37:@50989.4]
  wire  _T_905; // @[SRAM.scala 148:25:@50990.4]
  wire  _T_906; // @[SRAM.scala 148:15:@50991.4]
  wire  _T_907; // @[SRAM.scala 149:15:@50993.6]
  wire  _GEN_24; // @[SRAM.scala 148:48:@50992.4]
  reg  regs_25; // @[SRAM.scala 145:20:@50999.4]
  reg [31:0] _RAND_25;
  wire  _T_913; // @[SRAM.scala 148:37:@51000.4]
  wire  _T_914; // @[SRAM.scala 148:25:@51001.4]
  wire  _T_915; // @[SRAM.scala 148:15:@51002.4]
  wire  _T_916; // @[SRAM.scala 149:15:@51004.6]
  wire  _GEN_25; // @[SRAM.scala 148:48:@51003.4]
  reg  regs_26; // @[SRAM.scala 145:20:@51010.4]
  reg [31:0] _RAND_26;
  wire  _T_922; // @[SRAM.scala 148:37:@51011.4]
  wire  _T_923; // @[SRAM.scala 148:25:@51012.4]
  wire  _T_924; // @[SRAM.scala 148:15:@51013.4]
  wire  _T_925; // @[SRAM.scala 149:15:@51015.6]
  wire  _GEN_26; // @[SRAM.scala 148:48:@51014.4]
  reg  regs_27; // @[SRAM.scala 145:20:@51021.4]
  reg [31:0] _RAND_27;
  wire  _T_931; // @[SRAM.scala 148:37:@51022.4]
  wire  _T_932; // @[SRAM.scala 148:25:@51023.4]
  wire  _T_933; // @[SRAM.scala 148:15:@51024.4]
  wire  _T_934; // @[SRAM.scala 149:15:@51026.6]
  wire  _GEN_27; // @[SRAM.scala 148:48:@51025.4]
  reg  regs_28; // @[SRAM.scala 145:20:@51032.4]
  reg [31:0] _RAND_28;
  wire  _T_940; // @[SRAM.scala 148:37:@51033.4]
  wire  _T_941; // @[SRAM.scala 148:25:@51034.4]
  wire  _T_942; // @[SRAM.scala 148:15:@51035.4]
  wire  _T_943; // @[SRAM.scala 149:15:@51037.6]
  wire  _GEN_28; // @[SRAM.scala 148:48:@51036.4]
  reg  regs_29; // @[SRAM.scala 145:20:@51043.4]
  reg [31:0] _RAND_29;
  wire  _T_949; // @[SRAM.scala 148:37:@51044.4]
  wire  _T_950; // @[SRAM.scala 148:25:@51045.4]
  wire  _T_951; // @[SRAM.scala 148:15:@51046.4]
  wire  _T_952; // @[SRAM.scala 149:15:@51048.6]
  wire  _GEN_29; // @[SRAM.scala 148:48:@51047.4]
  reg  regs_30; // @[SRAM.scala 145:20:@51054.4]
  reg [31:0] _RAND_30;
  wire  _T_958; // @[SRAM.scala 148:37:@51055.4]
  wire  _T_959; // @[SRAM.scala 148:25:@51056.4]
  wire  _T_960; // @[SRAM.scala 148:15:@51057.4]
  wire  _T_961; // @[SRAM.scala 149:15:@51059.6]
  wire  _GEN_30; // @[SRAM.scala 148:48:@51058.4]
  reg  regs_31; // @[SRAM.scala 145:20:@51065.4]
  reg [31:0] _RAND_31;
  wire  _T_967; // @[SRAM.scala 148:37:@51066.4]
  wire  _T_968; // @[SRAM.scala 148:25:@51067.4]
  wire  _T_969; // @[SRAM.scala 148:15:@51068.4]
  wire  _T_970; // @[SRAM.scala 149:15:@51070.6]
  wire  _GEN_31; // @[SRAM.scala 148:48:@51069.4]
  reg  regs_32; // @[SRAM.scala 145:20:@51076.4]
  reg [31:0] _RAND_32;
  wire  _T_976; // @[SRAM.scala 148:37:@51077.4]
  wire  _T_977; // @[SRAM.scala 148:25:@51078.4]
  wire  _T_978; // @[SRAM.scala 148:15:@51079.4]
  wire  _T_979; // @[SRAM.scala 149:15:@51081.6]
  wire  _GEN_32; // @[SRAM.scala 148:48:@51080.4]
  reg  regs_33; // @[SRAM.scala 145:20:@51087.4]
  reg [31:0] _RAND_33;
  wire  _T_985; // @[SRAM.scala 148:37:@51088.4]
  wire  _T_986; // @[SRAM.scala 148:25:@51089.4]
  wire  _T_987; // @[SRAM.scala 148:15:@51090.4]
  wire  _T_988; // @[SRAM.scala 149:15:@51092.6]
  wire  _GEN_33; // @[SRAM.scala 148:48:@51091.4]
  reg  regs_34; // @[SRAM.scala 145:20:@51098.4]
  reg [31:0] _RAND_34;
  wire  _T_994; // @[SRAM.scala 148:37:@51099.4]
  wire  _T_995; // @[SRAM.scala 148:25:@51100.4]
  wire  _T_996; // @[SRAM.scala 148:15:@51101.4]
  wire  _T_997; // @[SRAM.scala 149:15:@51103.6]
  wire  _GEN_34; // @[SRAM.scala 148:48:@51102.4]
  reg  regs_35; // @[SRAM.scala 145:20:@51109.4]
  reg [31:0] _RAND_35;
  wire  _T_1003; // @[SRAM.scala 148:37:@51110.4]
  wire  _T_1004; // @[SRAM.scala 148:25:@51111.4]
  wire  _T_1005; // @[SRAM.scala 148:15:@51112.4]
  wire  _T_1006; // @[SRAM.scala 149:15:@51114.6]
  wire  _GEN_35; // @[SRAM.scala 148:48:@51113.4]
  reg  regs_36; // @[SRAM.scala 145:20:@51120.4]
  reg [31:0] _RAND_36;
  wire  _T_1012; // @[SRAM.scala 148:37:@51121.4]
  wire  _T_1013; // @[SRAM.scala 148:25:@51122.4]
  wire  _T_1014; // @[SRAM.scala 148:15:@51123.4]
  wire  _T_1015; // @[SRAM.scala 149:15:@51125.6]
  wire  _GEN_36; // @[SRAM.scala 148:48:@51124.4]
  reg  regs_37; // @[SRAM.scala 145:20:@51131.4]
  reg [31:0] _RAND_37;
  wire  _T_1021; // @[SRAM.scala 148:37:@51132.4]
  wire  _T_1022; // @[SRAM.scala 148:25:@51133.4]
  wire  _T_1023; // @[SRAM.scala 148:15:@51134.4]
  wire  _T_1024; // @[SRAM.scala 149:15:@51136.6]
  wire  _GEN_37; // @[SRAM.scala 148:48:@51135.4]
  reg  regs_38; // @[SRAM.scala 145:20:@51142.4]
  reg [31:0] _RAND_38;
  wire  _T_1030; // @[SRAM.scala 148:37:@51143.4]
  wire  _T_1031; // @[SRAM.scala 148:25:@51144.4]
  wire  _T_1032; // @[SRAM.scala 148:15:@51145.4]
  wire  _T_1033; // @[SRAM.scala 149:15:@51147.6]
  wire  _GEN_38; // @[SRAM.scala 148:48:@51146.4]
  reg  regs_39; // @[SRAM.scala 145:20:@51153.4]
  reg [31:0] _RAND_39;
  wire  _T_1039; // @[SRAM.scala 148:37:@51154.4]
  wire  _T_1040; // @[SRAM.scala 148:25:@51155.4]
  wire  _T_1041; // @[SRAM.scala 148:15:@51156.4]
  wire  _T_1042; // @[SRAM.scala 149:15:@51158.6]
  wire  _GEN_39; // @[SRAM.scala 148:48:@51157.4]
  reg  regs_40; // @[SRAM.scala 145:20:@51164.4]
  reg [31:0] _RAND_40;
  wire  _T_1048; // @[SRAM.scala 148:37:@51165.4]
  wire  _T_1049; // @[SRAM.scala 148:25:@51166.4]
  wire  _T_1050; // @[SRAM.scala 148:15:@51167.4]
  wire  _T_1051; // @[SRAM.scala 149:15:@51169.6]
  wire  _GEN_40; // @[SRAM.scala 148:48:@51168.4]
  reg  regs_41; // @[SRAM.scala 145:20:@51175.4]
  reg [31:0] _RAND_41;
  wire  _T_1057; // @[SRAM.scala 148:37:@51176.4]
  wire  _T_1058; // @[SRAM.scala 148:25:@51177.4]
  wire  _T_1059; // @[SRAM.scala 148:15:@51178.4]
  wire  _T_1060; // @[SRAM.scala 149:15:@51180.6]
  wire  _GEN_41; // @[SRAM.scala 148:48:@51179.4]
  reg  regs_42; // @[SRAM.scala 145:20:@51186.4]
  reg [31:0] _RAND_42;
  wire  _T_1066; // @[SRAM.scala 148:37:@51187.4]
  wire  _T_1067; // @[SRAM.scala 148:25:@51188.4]
  wire  _T_1068; // @[SRAM.scala 148:15:@51189.4]
  wire  _T_1069; // @[SRAM.scala 149:15:@51191.6]
  wire  _GEN_42; // @[SRAM.scala 148:48:@51190.4]
  reg  regs_43; // @[SRAM.scala 145:20:@51197.4]
  reg [31:0] _RAND_43;
  wire  _T_1075; // @[SRAM.scala 148:37:@51198.4]
  wire  _T_1076; // @[SRAM.scala 148:25:@51199.4]
  wire  _T_1077; // @[SRAM.scala 148:15:@51200.4]
  wire  _T_1078; // @[SRAM.scala 149:15:@51202.6]
  wire  _GEN_43; // @[SRAM.scala 148:48:@51201.4]
  reg  regs_44; // @[SRAM.scala 145:20:@51208.4]
  reg [31:0] _RAND_44;
  wire  _T_1084; // @[SRAM.scala 148:37:@51209.4]
  wire  _T_1085; // @[SRAM.scala 148:25:@51210.4]
  wire  _T_1086; // @[SRAM.scala 148:15:@51211.4]
  wire  _T_1087; // @[SRAM.scala 149:15:@51213.6]
  wire  _GEN_44; // @[SRAM.scala 148:48:@51212.4]
  reg  regs_45; // @[SRAM.scala 145:20:@51219.4]
  reg [31:0] _RAND_45;
  wire  _T_1093; // @[SRAM.scala 148:37:@51220.4]
  wire  _T_1094; // @[SRAM.scala 148:25:@51221.4]
  wire  _T_1095; // @[SRAM.scala 148:15:@51222.4]
  wire  _T_1096; // @[SRAM.scala 149:15:@51224.6]
  wire  _GEN_45; // @[SRAM.scala 148:48:@51223.4]
  reg  regs_46; // @[SRAM.scala 145:20:@51230.4]
  reg [31:0] _RAND_46;
  wire  _T_1102; // @[SRAM.scala 148:37:@51231.4]
  wire  _T_1103; // @[SRAM.scala 148:25:@51232.4]
  wire  _T_1104; // @[SRAM.scala 148:15:@51233.4]
  wire  _T_1105; // @[SRAM.scala 149:15:@51235.6]
  wire  _GEN_46; // @[SRAM.scala 148:48:@51234.4]
  reg  regs_47; // @[SRAM.scala 145:20:@51241.4]
  reg [31:0] _RAND_47;
  wire  _T_1111; // @[SRAM.scala 148:37:@51242.4]
  wire  _T_1112; // @[SRAM.scala 148:25:@51243.4]
  wire  _T_1113; // @[SRAM.scala 148:15:@51244.4]
  wire  _T_1114; // @[SRAM.scala 149:15:@51246.6]
  wire  _GEN_47; // @[SRAM.scala 148:48:@51245.4]
  reg  regs_48; // @[SRAM.scala 145:20:@51252.4]
  reg [31:0] _RAND_48;
  wire  _T_1120; // @[SRAM.scala 148:37:@51253.4]
  wire  _T_1121; // @[SRAM.scala 148:25:@51254.4]
  wire  _T_1122; // @[SRAM.scala 148:15:@51255.4]
  wire  _T_1123; // @[SRAM.scala 149:15:@51257.6]
  wire  _GEN_48; // @[SRAM.scala 148:48:@51256.4]
  reg  regs_49; // @[SRAM.scala 145:20:@51263.4]
  reg [31:0] _RAND_49;
  wire  _T_1129; // @[SRAM.scala 148:37:@51264.4]
  wire  _T_1130; // @[SRAM.scala 148:25:@51265.4]
  wire  _T_1131; // @[SRAM.scala 148:15:@51266.4]
  wire  _T_1132; // @[SRAM.scala 149:15:@51268.6]
  wire  _GEN_49; // @[SRAM.scala 148:48:@51267.4]
  reg  regs_50; // @[SRAM.scala 145:20:@51274.4]
  reg [31:0] _RAND_50;
  wire  _T_1138; // @[SRAM.scala 148:37:@51275.4]
  wire  _T_1139; // @[SRAM.scala 148:25:@51276.4]
  wire  _T_1140; // @[SRAM.scala 148:15:@51277.4]
  wire  _T_1141; // @[SRAM.scala 149:15:@51279.6]
  wire  _GEN_50; // @[SRAM.scala 148:48:@51278.4]
  reg  regs_51; // @[SRAM.scala 145:20:@51285.4]
  reg [31:0] _RAND_51;
  wire  _T_1147; // @[SRAM.scala 148:37:@51286.4]
  wire  _T_1148; // @[SRAM.scala 148:25:@51287.4]
  wire  _T_1149; // @[SRAM.scala 148:15:@51288.4]
  wire  _T_1150; // @[SRAM.scala 149:15:@51290.6]
  wire  _GEN_51; // @[SRAM.scala 148:48:@51289.4]
  reg  regs_52; // @[SRAM.scala 145:20:@51296.4]
  reg [31:0] _RAND_52;
  wire  _T_1156; // @[SRAM.scala 148:37:@51297.4]
  wire  _T_1157; // @[SRAM.scala 148:25:@51298.4]
  wire  _T_1158; // @[SRAM.scala 148:15:@51299.4]
  wire  _T_1159; // @[SRAM.scala 149:15:@51301.6]
  wire  _GEN_52; // @[SRAM.scala 148:48:@51300.4]
  reg  regs_53; // @[SRAM.scala 145:20:@51307.4]
  reg [31:0] _RAND_53;
  wire  _T_1165; // @[SRAM.scala 148:37:@51308.4]
  wire  _T_1166; // @[SRAM.scala 148:25:@51309.4]
  wire  _T_1167; // @[SRAM.scala 148:15:@51310.4]
  wire  _T_1168; // @[SRAM.scala 149:15:@51312.6]
  wire  _GEN_53; // @[SRAM.scala 148:48:@51311.4]
  reg  regs_54; // @[SRAM.scala 145:20:@51318.4]
  reg [31:0] _RAND_54;
  wire  _T_1174; // @[SRAM.scala 148:37:@51319.4]
  wire  _T_1175; // @[SRAM.scala 148:25:@51320.4]
  wire  _T_1176; // @[SRAM.scala 148:15:@51321.4]
  wire  _T_1177; // @[SRAM.scala 149:15:@51323.6]
  wire  _GEN_54; // @[SRAM.scala 148:48:@51322.4]
  reg  regs_55; // @[SRAM.scala 145:20:@51329.4]
  reg [31:0] _RAND_55;
  wire  _T_1183; // @[SRAM.scala 148:37:@51330.4]
  wire  _T_1184; // @[SRAM.scala 148:25:@51331.4]
  wire  _T_1185; // @[SRAM.scala 148:15:@51332.4]
  wire  _T_1186; // @[SRAM.scala 149:15:@51334.6]
  wire  _GEN_55; // @[SRAM.scala 148:48:@51333.4]
  reg  regs_56; // @[SRAM.scala 145:20:@51340.4]
  reg [31:0] _RAND_56;
  wire  _T_1192; // @[SRAM.scala 148:37:@51341.4]
  wire  _T_1193; // @[SRAM.scala 148:25:@51342.4]
  wire  _T_1194; // @[SRAM.scala 148:15:@51343.4]
  wire  _T_1195; // @[SRAM.scala 149:15:@51345.6]
  wire  _GEN_56; // @[SRAM.scala 148:48:@51344.4]
  reg  regs_57; // @[SRAM.scala 145:20:@51351.4]
  reg [31:0] _RAND_57;
  wire  _T_1201; // @[SRAM.scala 148:37:@51352.4]
  wire  _T_1202; // @[SRAM.scala 148:25:@51353.4]
  wire  _T_1203; // @[SRAM.scala 148:15:@51354.4]
  wire  _T_1204; // @[SRAM.scala 149:15:@51356.6]
  wire  _GEN_57; // @[SRAM.scala 148:48:@51355.4]
  reg  regs_58; // @[SRAM.scala 145:20:@51362.4]
  reg [31:0] _RAND_58;
  wire  _T_1210; // @[SRAM.scala 148:37:@51363.4]
  wire  _T_1211; // @[SRAM.scala 148:25:@51364.4]
  wire  _T_1212; // @[SRAM.scala 148:15:@51365.4]
  wire  _T_1213; // @[SRAM.scala 149:15:@51367.6]
  wire  _GEN_58; // @[SRAM.scala 148:48:@51366.4]
  reg  regs_59; // @[SRAM.scala 145:20:@51373.4]
  reg [31:0] _RAND_59;
  wire  _T_1219; // @[SRAM.scala 148:37:@51374.4]
  wire  _T_1220; // @[SRAM.scala 148:25:@51375.4]
  wire  _T_1221; // @[SRAM.scala 148:15:@51376.4]
  wire  _T_1222; // @[SRAM.scala 149:15:@51378.6]
  wire  _GEN_59; // @[SRAM.scala 148:48:@51377.4]
  reg  regs_60; // @[SRAM.scala 145:20:@51384.4]
  reg [31:0] _RAND_60;
  wire  _T_1228; // @[SRAM.scala 148:37:@51385.4]
  wire  _T_1229; // @[SRAM.scala 148:25:@51386.4]
  wire  _T_1230; // @[SRAM.scala 148:15:@51387.4]
  wire  _T_1231; // @[SRAM.scala 149:15:@51389.6]
  wire  _GEN_60; // @[SRAM.scala 148:48:@51388.4]
  reg  regs_61; // @[SRAM.scala 145:20:@51395.4]
  reg [31:0] _RAND_61;
  wire  _T_1237; // @[SRAM.scala 148:37:@51396.4]
  wire  _T_1238; // @[SRAM.scala 148:25:@51397.4]
  wire  _T_1239; // @[SRAM.scala 148:15:@51398.4]
  wire  _T_1240; // @[SRAM.scala 149:15:@51400.6]
  wire  _GEN_61; // @[SRAM.scala 148:48:@51399.4]
  reg  regs_62; // @[SRAM.scala 145:20:@51406.4]
  reg [31:0] _RAND_62;
  wire  _T_1246; // @[SRAM.scala 148:37:@51407.4]
  wire  _T_1247; // @[SRAM.scala 148:25:@51408.4]
  wire  _T_1248; // @[SRAM.scala 148:15:@51409.4]
  wire  _T_1249; // @[SRAM.scala 149:15:@51411.6]
  wire  _GEN_62; // @[SRAM.scala 148:48:@51410.4]
  reg  regs_63; // @[SRAM.scala 145:20:@51417.4]
  reg [31:0] _RAND_63;
  wire  _T_1255; // @[SRAM.scala 148:37:@51418.4]
  wire  _T_1256; // @[SRAM.scala 148:25:@51419.4]
  wire  _T_1257; // @[SRAM.scala 148:15:@51420.4]
  wire  _T_1258; // @[SRAM.scala 149:15:@51422.6]
  wire  _GEN_63; // @[SRAM.scala 148:48:@51421.4]
  wire  _GEN_65; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_66; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_67; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_68; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_69; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_70; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_71; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_72; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_73; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_74; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_75; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_76; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_77; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_78; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_79; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_80; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_81; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_82; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_83; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_84; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_85; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_86; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_87; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_88; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_89; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_90; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_91; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_92; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_93; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_94; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_95; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_96; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_97; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_98; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_99; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_100; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_101; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_102; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_103; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_104; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_105; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_106; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_107; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_108; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_109; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_110; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_111; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_112; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_113; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_114; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_115; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_116; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_117; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_118; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_119; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_120; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_121; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_122; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_123; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_124; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_125; // @[SRAM.scala 155:12:@51491.4]
  wire  _GEN_126; // @[SRAM.scala 155:12:@51491.4]
  assign _T_688 = io_waddr == 6'h0; // @[SRAM.scala 148:37:@50725.4]
  assign _T_689 = io_wen & _T_688; // @[SRAM.scala 148:25:@50726.4]
  assign _T_690 = io_banks_0_wdata_valid | _T_689; // @[SRAM.scala 148:15:@50727.4]
  assign _T_691 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50729.6]
  assign _GEN_0 = _T_690 ? _T_691 : regs_0; // @[SRAM.scala 148:48:@50728.4]
  assign _T_697 = io_waddr == 6'h1; // @[SRAM.scala 148:37:@50736.4]
  assign _T_698 = io_wen & _T_697; // @[SRAM.scala 148:25:@50737.4]
  assign _T_699 = io_banks_1_wdata_valid | _T_698; // @[SRAM.scala 148:15:@50738.4]
  assign _T_700 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50740.6]
  assign _GEN_1 = _T_699 ? _T_700 : regs_1; // @[SRAM.scala 148:48:@50739.4]
  assign _T_706 = io_waddr == 6'h2; // @[SRAM.scala 148:37:@50747.4]
  assign _T_707 = io_wen & _T_706; // @[SRAM.scala 148:25:@50748.4]
  assign _T_708 = io_banks_2_wdata_valid | _T_707; // @[SRAM.scala 148:15:@50749.4]
  assign _T_709 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50751.6]
  assign _GEN_2 = _T_708 ? _T_709 : regs_2; // @[SRAM.scala 148:48:@50750.4]
  assign _T_715 = io_waddr == 6'h3; // @[SRAM.scala 148:37:@50758.4]
  assign _T_716 = io_wen & _T_715; // @[SRAM.scala 148:25:@50759.4]
  assign _T_717 = io_banks_3_wdata_valid | _T_716; // @[SRAM.scala 148:15:@50760.4]
  assign _T_718 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50762.6]
  assign _GEN_3 = _T_717 ? _T_718 : regs_3; // @[SRAM.scala 148:48:@50761.4]
  assign _T_724 = io_waddr == 6'h4; // @[SRAM.scala 148:37:@50769.4]
  assign _T_725 = io_wen & _T_724; // @[SRAM.scala 148:25:@50770.4]
  assign _T_726 = io_banks_4_wdata_valid | _T_725; // @[SRAM.scala 148:15:@50771.4]
  assign _T_727 = io_banks_4_wdata_valid ? io_banks_4_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50773.6]
  assign _GEN_4 = _T_726 ? _T_727 : regs_4; // @[SRAM.scala 148:48:@50772.4]
  assign _T_733 = io_waddr == 6'h5; // @[SRAM.scala 148:37:@50780.4]
  assign _T_734 = io_wen & _T_733; // @[SRAM.scala 148:25:@50781.4]
  assign _T_735 = io_banks_5_wdata_valid | _T_734; // @[SRAM.scala 148:15:@50782.4]
  assign _T_736 = io_banks_5_wdata_valid ? io_banks_5_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50784.6]
  assign _GEN_5 = _T_735 ? _T_736 : regs_5; // @[SRAM.scala 148:48:@50783.4]
  assign _T_742 = io_waddr == 6'h6; // @[SRAM.scala 148:37:@50791.4]
  assign _T_743 = io_wen & _T_742; // @[SRAM.scala 148:25:@50792.4]
  assign _T_744 = io_banks_6_wdata_valid | _T_743; // @[SRAM.scala 148:15:@50793.4]
  assign _T_745 = io_banks_6_wdata_valid ? io_banks_6_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50795.6]
  assign _GEN_6 = _T_744 ? _T_745 : regs_6; // @[SRAM.scala 148:48:@50794.4]
  assign _T_751 = io_waddr == 6'h7; // @[SRAM.scala 148:37:@50802.4]
  assign _T_752 = io_wen & _T_751; // @[SRAM.scala 148:25:@50803.4]
  assign _T_753 = io_banks_7_wdata_valid | _T_752; // @[SRAM.scala 148:15:@50804.4]
  assign _T_754 = io_banks_7_wdata_valid ? io_banks_7_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50806.6]
  assign _GEN_7 = _T_753 ? _T_754 : regs_7; // @[SRAM.scala 148:48:@50805.4]
  assign _T_760 = io_waddr == 6'h8; // @[SRAM.scala 148:37:@50813.4]
  assign _T_761 = io_wen & _T_760; // @[SRAM.scala 148:25:@50814.4]
  assign _T_762 = io_banks_8_wdata_valid | _T_761; // @[SRAM.scala 148:15:@50815.4]
  assign _T_763 = io_banks_8_wdata_valid ? io_banks_8_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50817.6]
  assign _GEN_8 = _T_762 ? _T_763 : regs_8; // @[SRAM.scala 148:48:@50816.4]
  assign _T_769 = io_waddr == 6'h9; // @[SRAM.scala 148:37:@50824.4]
  assign _T_770 = io_wen & _T_769; // @[SRAM.scala 148:25:@50825.4]
  assign _T_771 = io_banks_9_wdata_valid | _T_770; // @[SRAM.scala 148:15:@50826.4]
  assign _T_772 = io_banks_9_wdata_valid ? io_banks_9_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50828.6]
  assign _GEN_9 = _T_771 ? _T_772 : regs_9; // @[SRAM.scala 148:48:@50827.4]
  assign _T_778 = io_waddr == 6'ha; // @[SRAM.scala 148:37:@50835.4]
  assign _T_779 = io_wen & _T_778; // @[SRAM.scala 148:25:@50836.4]
  assign _T_780 = io_banks_10_wdata_valid | _T_779; // @[SRAM.scala 148:15:@50837.4]
  assign _T_781 = io_banks_10_wdata_valid ? io_banks_10_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50839.6]
  assign _GEN_10 = _T_780 ? _T_781 : regs_10; // @[SRAM.scala 148:48:@50838.4]
  assign _T_787 = io_waddr == 6'hb; // @[SRAM.scala 148:37:@50846.4]
  assign _T_788 = io_wen & _T_787; // @[SRAM.scala 148:25:@50847.4]
  assign _T_789 = io_banks_11_wdata_valid | _T_788; // @[SRAM.scala 148:15:@50848.4]
  assign _T_790 = io_banks_11_wdata_valid ? io_banks_11_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50850.6]
  assign _GEN_11 = _T_789 ? _T_790 : regs_11; // @[SRAM.scala 148:48:@50849.4]
  assign _T_796 = io_waddr == 6'hc; // @[SRAM.scala 148:37:@50857.4]
  assign _T_797 = io_wen & _T_796; // @[SRAM.scala 148:25:@50858.4]
  assign _T_798 = io_banks_12_wdata_valid | _T_797; // @[SRAM.scala 148:15:@50859.4]
  assign _T_799 = io_banks_12_wdata_valid ? io_banks_12_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50861.6]
  assign _GEN_12 = _T_798 ? _T_799 : regs_12; // @[SRAM.scala 148:48:@50860.4]
  assign _T_805 = io_waddr == 6'hd; // @[SRAM.scala 148:37:@50868.4]
  assign _T_806 = io_wen & _T_805; // @[SRAM.scala 148:25:@50869.4]
  assign _T_807 = io_banks_13_wdata_valid | _T_806; // @[SRAM.scala 148:15:@50870.4]
  assign _T_808 = io_banks_13_wdata_valid ? io_banks_13_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50872.6]
  assign _GEN_13 = _T_807 ? _T_808 : regs_13; // @[SRAM.scala 148:48:@50871.4]
  assign _T_814 = io_waddr == 6'he; // @[SRAM.scala 148:37:@50879.4]
  assign _T_815 = io_wen & _T_814; // @[SRAM.scala 148:25:@50880.4]
  assign _T_816 = io_banks_14_wdata_valid | _T_815; // @[SRAM.scala 148:15:@50881.4]
  assign _T_817 = io_banks_14_wdata_valid ? io_banks_14_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50883.6]
  assign _GEN_14 = _T_816 ? _T_817 : regs_14; // @[SRAM.scala 148:48:@50882.4]
  assign _T_823 = io_waddr == 6'hf; // @[SRAM.scala 148:37:@50890.4]
  assign _T_824 = io_wen & _T_823; // @[SRAM.scala 148:25:@50891.4]
  assign _T_825 = io_banks_15_wdata_valid | _T_824; // @[SRAM.scala 148:15:@50892.4]
  assign _T_826 = io_banks_15_wdata_valid ? io_banks_15_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50894.6]
  assign _GEN_15 = _T_825 ? _T_826 : regs_15; // @[SRAM.scala 148:48:@50893.4]
  assign _T_832 = io_waddr == 6'h10; // @[SRAM.scala 148:37:@50901.4]
  assign _T_833 = io_wen & _T_832; // @[SRAM.scala 148:25:@50902.4]
  assign _T_834 = io_banks_16_wdata_valid | _T_833; // @[SRAM.scala 148:15:@50903.4]
  assign _T_835 = io_banks_16_wdata_valid ? io_banks_16_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50905.6]
  assign _GEN_16 = _T_834 ? _T_835 : regs_16; // @[SRAM.scala 148:48:@50904.4]
  assign _T_841 = io_waddr == 6'h11; // @[SRAM.scala 148:37:@50912.4]
  assign _T_842 = io_wen & _T_841; // @[SRAM.scala 148:25:@50913.4]
  assign _T_843 = io_banks_17_wdata_valid | _T_842; // @[SRAM.scala 148:15:@50914.4]
  assign _T_844 = io_banks_17_wdata_valid ? io_banks_17_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50916.6]
  assign _GEN_17 = _T_843 ? _T_844 : regs_17; // @[SRAM.scala 148:48:@50915.4]
  assign _T_850 = io_waddr == 6'h12; // @[SRAM.scala 148:37:@50923.4]
  assign _T_851 = io_wen & _T_850; // @[SRAM.scala 148:25:@50924.4]
  assign _T_852 = io_banks_18_wdata_valid | _T_851; // @[SRAM.scala 148:15:@50925.4]
  assign _T_853 = io_banks_18_wdata_valid ? io_banks_18_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50927.6]
  assign _GEN_18 = _T_852 ? _T_853 : regs_18; // @[SRAM.scala 148:48:@50926.4]
  assign _T_859 = io_waddr == 6'h13; // @[SRAM.scala 148:37:@50934.4]
  assign _T_860 = io_wen & _T_859; // @[SRAM.scala 148:25:@50935.4]
  assign _T_861 = io_banks_19_wdata_valid | _T_860; // @[SRAM.scala 148:15:@50936.4]
  assign _T_862 = io_banks_19_wdata_valid ? io_banks_19_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50938.6]
  assign _GEN_19 = _T_861 ? _T_862 : regs_19; // @[SRAM.scala 148:48:@50937.4]
  assign _T_868 = io_waddr == 6'h14; // @[SRAM.scala 148:37:@50945.4]
  assign _T_869 = io_wen & _T_868; // @[SRAM.scala 148:25:@50946.4]
  assign _T_870 = io_banks_20_wdata_valid | _T_869; // @[SRAM.scala 148:15:@50947.4]
  assign _T_871 = io_banks_20_wdata_valid ? io_banks_20_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50949.6]
  assign _GEN_20 = _T_870 ? _T_871 : regs_20; // @[SRAM.scala 148:48:@50948.4]
  assign _T_877 = io_waddr == 6'h15; // @[SRAM.scala 148:37:@50956.4]
  assign _T_878 = io_wen & _T_877; // @[SRAM.scala 148:25:@50957.4]
  assign _T_879 = io_banks_21_wdata_valid | _T_878; // @[SRAM.scala 148:15:@50958.4]
  assign _T_880 = io_banks_21_wdata_valid ? io_banks_21_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50960.6]
  assign _GEN_21 = _T_879 ? _T_880 : regs_21; // @[SRAM.scala 148:48:@50959.4]
  assign _T_886 = io_waddr == 6'h16; // @[SRAM.scala 148:37:@50967.4]
  assign _T_887 = io_wen & _T_886; // @[SRAM.scala 148:25:@50968.4]
  assign _T_888 = io_banks_22_wdata_valid | _T_887; // @[SRAM.scala 148:15:@50969.4]
  assign _T_889 = io_banks_22_wdata_valid ? io_banks_22_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50971.6]
  assign _GEN_22 = _T_888 ? _T_889 : regs_22; // @[SRAM.scala 148:48:@50970.4]
  assign _T_895 = io_waddr == 6'h17; // @[SRAM.scala 148:37:@50978.4]
  assign _T_896 = io_wen & _T_895; // @[SRAM.scala 148:25:@50979.4]
  assign _T_897 = io_banks_23_wdata_valid | _T_896; // @[SRAM.scala 148:15:@50980.4]
  assign _T_898 = io_banks_23_wdata_valid ? io_banks_23_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50982.6]
  assign _GEN_23 = _T_897 ? _T_898 : regs_23; // @[SRAM.scala 148:48:@50981.4]
  assign _T_904 = io_waddr == 6'h18; // @[SRAM.scala 148:37:@50989.4]
  assign _T_905 = io_wen & _T_904; // @[SRAM.scala 148:25:@50990.4]
  assign _T_906 = io_banks_24_wdata_valid | _T_905; // @[SRAM.scala 148:15:@50991.4]
  assign _T_907 = io_banks_24_wdata_valid ? io_banks_24_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@50993.6]
  assign _GEN_24 = _T_906 ? _T_907 : regs_24; // @[SRAM.scala 148:48:@50992.4]
  assign _T_913 = io_waddr == 6'h19; // @[SRAM.scala 148:37:@51000.4]
  assign _T_914 = io_wen & _T_913; // @[SRAM.scala 148:25:@51001.4]
  assign _T_915 = io_banks_25_wdata_valid | _T_914; // @[SRAM.scala 148:15:@51002.4]
  assign _T_916 = io_banks_25_wdata_valid ? io_banks_25_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51004.6]
  assign _GEN_25 = _T_915 ? _T_916 : regs_25; // @[SRAM.scala 148:48:@51003.4]
  assign _T_922 = io_waddr == 6'h1a; // @[SRAM.scala 148:37:@51011.4]
  assign _T_923 = io_wen & _T_922; // @[SRAM.scala 148:25:@51012.4]
  assign _T_924 = io_banks_26_wdata_valid | _T_923; // @[SRAM.scala 148:15:@51013.4]
  assign _T_925 = io_banks_26_wdata_valid ? io_banks_26_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51015.6]
  assign _GEN_26 = _T_924 ? _T_925 : regs_26; // @[SRAM.scala 148:48:@51014.4]
  assign _T_931 = io_waddr == 6'h1b; // @[SRAM.scala 148:37:@51022.4]
  assign _T_932 = io_wen & _T_931; // @[SRAM.scala 148:25:@51023.4]
  assign _T_933 = io_banks_27_wdata_valid | _T_932; // @[SRAM.scala 148:15:@51024.4]
  assign _T_934 = io_banks_27_wdata_valid ? io_banks_27_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51026.6]
  assign _GEN_27 = _T_933 ? _T_934 : regs_27; // @[SRAM.scala 148:48:@51025.4]
  assign _T_940 = io_waddr == 6'h1c; // @[SRAM.scala 148:37:@51033.4]
  assign _T_941 = io_wen & _T_940; // @[SRAM.scala 148:25:@51034.4]
  assign _T_942 = io_banks_28_wdata_valid | _T_941; // @[SRAM.scala 148:15:@51035.4]
  assign _T_943 = io_banks_28_wdata_valid ? io_banks_28_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51037.6]
  assign _GEN_28 = _T_942 ? _T_943 : regs_28; // @[SRAM.scala 148:48:@51036.4]
  assign _T_949 = io_waddr == 6'h1d; // @[SRAM.scala 148:37:@51044.4]
  assign _T_950 = io_wen & _T_949; // @[SRAM.scala 148:25:@51045.4]
  assign _T_951 = io_banks_29_wdata_valid | _T_950; // @[SRAM.scala 148:15:@51046.4]
  assign _T_952 = io_banks_29_wdata_valid ? io_banks_29_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51048.6]
  assign _GEN_29 = _T_951 ? _T_952 : regs_29; // @[SRAM.scala 148:48:@51047.4]
  assign _T_958 = io_waddr == 6'h1e; // @[SRAM.scala 148:37:@51055.4]
  assign _T_959 = io_wen & _T_958; // @[SRAM.scala 148:25:@51056.4]
  assign _T_960 = io_banks_30_wdata_valid | _T_959; // @[SRAM.scala 148:15:@51057.4]
  assign _T_961 = io_banks_30_wdata_valid ? io_banks_30_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51059.6]
  assign _GEN_30 = _T_960 ? _T_961 : regs_30; // @[SRAM.scala 148:48:@51058.4]
  assign _T_967 = io_waddr == 6'h1f; // @[SRAM.scala 148:37:@51066.4]
  assign _T_968 = io_wen & _T_967; // @[SRAM.scala 148:25:@51067.4]
  assign _T_969 = io_banks_31_wdata_valid | _T_968; // @[SRAM.scala 148:15:@51068.4]
  assign _T_970 = io_banks_31_wdata_valid ? io_banks_31_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51070.6]
  assign _GEN_31 = _T_969 ? _T_970 : regs_31; // @[SRAM.scala 148:48:@51069.4]
  assign _T_976 = io_waddr == 6'h20; // @[SRAM.scala 148:37:@51077.4]
  assign _T_977 = io_wen & _T_976; // @[SRAM.scala 148:25:@51078.4]
  assign _T_978 = io_banks_32_wdata_valid | _T_977; // @[SRAM.scala 148:15:@51079.4]
  assign _T_979 = io_banks_32_wdata_valid ? io_banks_32_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51081.6]
  assign _GEN_32 = _T_978 ? _T_979 : regs_32; // @[SRAM.scala 148:48:@51080.4]
  assign _T_985 = io_waddr == 6'h21; // @[SRAM.scala 148:37:@51088.4]
  assign _T_986 = io_wen & _T_985; // @[SRAM.scala 148:25:@51089.4]
  assign _T_987 = io_banks_33_wdata_valid | _T_986; // @[SRAM.scala 148:15:@51090.4]
  assign _T_988 = io_banks_33_wdata_valid ? io_banks_33_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51092.6]
  assign _GEN_33 = _T_987 ? _T_988 : regs_33; // @[SRAM.scala 148:48:@51091.4]
  assign _T_994 = io_waddr == 6'h22; // @[SRAM.scala 148:37:@51099.4]
  assign _T_995 = io_wen & _T_994; // @[SRAM.scala 148:25:@51100.4]
  assign _T_996 = io_banks_34_wdata_valid | _T_995; // @[SRAM.scala 148:15:@51101.4]
  assign _T_997 = io_banks_34_wdata_valid ? io_banks_34_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51103.6]
  assign _GEN_34 = _T_996 ? _T_997 : regs_34; // @[SRAM.scala 148:48:@51102.4]
  assign _T_1003 = io_waddr == 6'h23; // @[SRAM.scala 148:37:@51110.4]
  assign _T_1004 = io_wen & _T_1003; // @[SRAM.scala 148:25:@51111.4]
  assign _T_1005 = io_banks_35_wdata_valid | _T_1004; // @[SRAM.scala 148:15:@51112.4]
  assign _T_1006 = io_banks_35_wdata_valid ? io_banks_35_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51114.6]
  assign _GEN_35 = _T_1005 ? _T_1006 : regs_35; // @[SRAM.scala 148:48:@51113.4]
  assign _T_1012 = io_waddr == 6'h24; // @[SRAM.scala 148:37:@51121.4]
  assign _T_1013 = io_wen & _T_1012; // @[SRAM.scala 148:25:@51122.4]
  assign _T_1014 = io_banks_36_wdata_valid | _T_1013; // @[SRAM.scala 148:15:@51123.4]
  assign _T_1015 = io_banks_36_wdata_valid ? io_banks_36_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51125.6]
  assign _GEN_36 = _T_1014 ? _T_1015 : regs_36; // @[SRAM.scala 148:48:@51124.4]
  assign _T_1021 = io_waddr == 6'h25; // @[SRAM.scala 148:37:@51132.4]
  assign _T_1022 = io_wen & _T_1021; // @[SRAM.scala 148:25:@51133.4]
  assign _T_1023 = io_banks_37_wdata_valid | _T_1022; // @[SRAM.scala 148:15:@51134.4]
  assign _T_1024 = io_banks_37_wdata_valid ? io_banks_37_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51136.6]
  assign _GEN_37 = _T_1023 ? _T_1024 : regs_37; // @[SRAM.scala 148:48:@51135.4]
  assign _T_1030 = io_waddr == 6'h26; // @[SRAM.scala 148:37:@51143.4]
  assign _T_1031 = io_wen & _T_1030; // @[SRAM.scala 148:25:@51144.4]
  assign _T_1032 = io_banks_38_wdata_valid | _T_1031; // @[SRAM.scala 148:15:@51145.4]
  assign _T_1033 = io_banks_38_wdata_valid ? io_banks_38_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51147.6]
  assign _GEN_38 = _T_1032 ? _T_1033 : regs_38; // @[SRAM.scala 148:48:@51146.4]
  assign _T_1039 = io_waddr == 6'h27; // @[SRAM.scala 148:37:@51154.4]
  assign _T_1040 = io_wen & _T_1039; // @[SRAM.scala 148:25:@51155.4]
  assign _T_1041 = io_banks_39_wdata_valid | _T_1040; // @[SRAM.scala 148:15:@51156.4]
  assign _T_1042 = io_banks_39_wdata_valid ? io_banks_39_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51158.6]
  assign _GEN_39 = _T_1041 ? _T_1042 : regs_39; // @[SRAM.scala 148:48:@51157.4]
  assign _T_1048 = io_waddr == 6'h28; // @[SRAM.scala 148:37:@51165.4]
  assign _T_1049 = io_wen & _T_1048; // @[SRAM.scala 148:25:@51166.4]
  assign _T_1050 = io_banks_40_wdata_valid | _T_1049; // @[SRAM.scala 148:15:@51167.4]
  assign _T_1051 = io_banks_40_wdata_valid ? io_banks_40_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51169.6]
  assign _GEN_40 = _T_1050 ? _T_1051 : regs_40; // @[SRAM.scala 148:48:@51168.4]
  assign _T_1057 = io_waddr == 6'h29; // @[SRAM.scala 148:37:@51176.4]
  assign _T_1058 = io_wen & _T_1057; // @[SRAM.scala 148:25:@51177.4]
  assign _T_1059 = io_banks_41_wdata_valid | _T_1058; // @[SRAM.scala 148:15:@51178.4]
  assign _T_1060 = io_banks_41_wdata_valid ? io_banks_41_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51180.6]
  assign _GEN_41 = _T_1059 ? _T_1060 : regs_41; // @[SRAM.scala 148:48:@51179.4]
  assign _T_1066 = io_waddr == 6'h2a; // @[SRAM.scala 148:37:@51187.4]
  assign _T_1067 = io_wen & _T_1066; // @[SRAM.scala 148:25:@51188.4]
  assign _T_1068 = io_banks_42_wdata_valid | _T_1067; // @[SRAM.scala 148:15:@51189.4]
  assign _T_1069 = io_banks_42_wdata_valid ? io_banks_42_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51191.6]
  assign _GEN_42 = _T_1068 ? _T_1069 : regs_42; // @[SRAM.scala 148:48:@51190.4]
  assign _T_1075 = io_waddr == 6'h2b; // @[SRAM.scala 148:37:@51198.4]
  assign _T_1076 = io_wen & _T_1075; // @[SRAM.scala 148:25:@51199.4]
  assign _T_1077 = io_banks_43_wdata_valid | _T_1076; // @[SRAM.scala 148:15:@51200.4]
  assign _T_1078 = io_banks_43_wdata_valid ? io_banks_43_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51202.6]
  assign _GEN_43 = _T_1077 ? _T_1078 : regs_43; // @[SRAM.scala 148:48:@51201.4]
  assign _T_1084 = io_waddr == 6'h2c; // @[SRAM.scala 148:37:@51209.4]
  assign _T_1085 = io_wen & _T_1084; // @[SRAM.scala 148:25:@51210.4]
  assign _T_1086 = io_banks_44_wdata_valid | _T_1085; // @[SRAM.scala 148:15:@51211.4]
  assign _T_1087 = io_banks_44_wdata_valid ? io_banks_44_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51213.6]
  assign _GEN_44 = _T_1086 ? _T_1087 : regs_44; // @[SRAM.scala 148:48:@51212.4]
  assign _T_1093 = io_waddr == 6'h2d; // @[SRAM.scala 148:37:@51220.4]
  assign _T_1094 = io_wen & _T_1093; // @[SRAM.scala 148:25:@51221.4]
  assign _T_1095 = io_banks_45_wdata_valid | _T_1094; // @[SRAM.scala 148:15:@51222.4]
  assign _T_1096 = io_banks_45_wdata_valid ? io_banks_45_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51224.6]
  assign _GEN_45 = _T_1095 ? _T_1096 : regs_45; // @[SRAM.scala 148:48:@51223.4]
  assign _T_1102 = io_waddr == 6'h2e; // @[SRAM.scala 148:37:@51231.4]
  assign _T_1103 = io_wen & _T_1102; // @[SRAM.scala 148:25:@51232.4]
  assign _T_1104 = io_banks_46_wdata_valid | _T_1103; // @[SRAM.scala 148:15:@51233.4]
  assign _T_1105 = io_banks_46_wdata_valid ? io_banks_46_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51235.6]
  assign _GEN_46 = _T_1104 ? _T_1105 : regs_46; // @[SRAM.scala 148:48:@51234.4]
  assign _T_1111 = io_waddr == 6'h2f; // @[SRAM.scala 148:37:@51242.4]
  assign _T_1112 = io_wen & _T_1111; // @[SRAM.scala 148:25:@51243.4]
  assign _T_1113 = io_banks_47_wdata_valid | _T_1112; // @[SRAM.scala 148:15:@51244.4]
  assign _T_1114 = io_banks_47_wdata_valid ? io_banks_47_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51246.6]
  assign _GEN_47 = _T_1113 ? _T_1114 : regs_47; // @[SRAM.scala 148:48:@51245.4]
  assign _T_1120 = io_waddr == 6'h30; // @[SRAM.scala 148:37:@51253.4]
  assign _T_1121 = io_wen & _T_1120; // @[SRAM.scala 148:25:@51254.4]
  assign _T_1122 = io_banks_48_wdata_valid | _T_1121; // @[SRAM.scala 148:15:@51255.4]
  assign _T_1123 = io_banks_48_wdata_valid ? io_banks_48_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51257.6]
  assign _GEN_48 = _T_1122 ? _T_1123 : regs_48; // @[SRAM.scala 148:48:@51256.4]
  assign _T_1129 = io_waddr == 6'h31; // @[SRAM.scala 148:37:@51264.4]
  assign _T_1130 = io_wen & _T_1129; // @[SRAM.scala 148:25:@51265.4]
  assign _T_1131 = io_banks_49_wdata_valid | _T_1130; // @[SRAM.scala 148:15:@51266.4]
  assign _T_1132 = io_banks_49_wdata_valid ? io_banks_49_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51268.6]
  assign _GEN_49 = _T_1131 ? _T_1132 : regs_49; // @[SRAM.scala 148:48:@51267.4]
  assign _T_1138 = io_waddr == 6'h32; // @[SRAM.scala 148:37:@51275.4]
  assign _T_1139 = io_wen & _T_1138; // @[SRAM.scala 148:25:@51276.4]
  assign _T_1140 = io_banks_50_wdata_valid | _T_1139; // @[SRAM.scala 148:15:@51277.4]
  assign _T_1141 = io_banks_50_wdata_valid ? io_banks_50_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51279.6]
  assign _GEN_50 = _T_1140 ? _T_1141 : regs_50; // @[SRAM.scala 148:48:@51278.4]
  assign _T_1147 = io_waddr == 6'h33; // @[SRAM.scala 148:37:@51286.4]
  assign _T_1148 = io_wen & _T_1147; // @[SRAM.scala 148:25:@51287.4]
  assign _T_1149 = io_banks_51_wdata_valid | _T_1148; // @[SRAM.scala 148:15:@51288.4]
  assign _T_1150 = io_banks_51_wdata_valid ? io_banks_51_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51290.6]
  assign _GEN_51 = _T_1149 ? _T_1150 : regs_51; // @[SRAM.scala 148:48:@51289.4]
  assign _T_1156 = io_waddr == 6'h34; // @[SRAM.scala 148:37:@51297.4]
  assign _T_1157 = io_wen & _T_1156; // @[SRAM.scala 148:25:@51298.4]
  assign _T_1158 = io_banks_52_wdata_valid | _T_1157; // @[SRAM.scala 148:15:@51299.4]
  assign _T_1159 = io_banks_52_wdata_valid ? io_banks_52_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51301.6]
  assign _GEN_52 = _T_1158 ? _T_1159 : regs_52; // @[SRAM.scala 148:48:@51300.4]
  assign _T_1165 = io_waddr == 6'h35; // @[SRAM.scala 148:37:@51308.4]
  assign _T_1166 = io_wen & _T_1165; // @[SRAM.scala 148:25:@51309.4]
  assign _T_1167 = io_banks_53_wdata_valid | _T_1166; // @[SRAM.scala 148:15:@51310.4]
  assign _T_1168 = io_banks_53_wdata_valid ? io_banks_53_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51312.6]
  assign _GEN_53 = _T_1167 ? _T_1168 : regs_53; // @[SRAM.scala 148:48:@51311.4]
  assign _T_1174 = io_waddr == 6'h36; // @[SRAM.scala 148:37:@51319.4]
  assign _T_1175 = io_wen & _T_1174; // @[SRAM.scala 148:25:@51320.4]
  assign _T_1176 = io_banks_54_wdata_valid | _T_1175; // @[SRAM.scala 148:15:@51321.4]
  assign _T_1177 = io_banks_54_wdata_valid ? io_banks_54_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51323.6]
  assign _GEN_54 = _T_1176 ? _T_1177 : regs_54; // @[SRAM.scala 148:48:@51322.4]
  assign _T_1183 = io_waddr == 6'h37; // @[SRAM.scala 148:37:@51330.4]
  assign _T_1184 = io_wen & _T_1183; // @[SRAM.scala 148:25:@51331.4]
  assign _T_1185 = io_banks_55_wdata_valid | _T_1184; // @[SRAM.scala 148:15:@51332.4]
  assign _T_1186 = io_banks_55_wdata_valid ? io_banks_55_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51334.6]
  assign _GEN_55 = _T_1185 ? _T_1186 : regs_55; // @[SRAM.scala 148:48:@51333.4]
  assign _T_1192 = io_waddr == 6'h38; // @[SRAM.scala 148:37:@51341.4]
  assign _T_1193 = io_wen & _T_1192; // @[SRAM.scala 148:25:@51342.4]
  assign _T_1194 = io_banks_56_wdata_valid | _T_1193; // @[SRAM.scala 148:15:@51343.4]
  assign _T_1195 = io_banks_56_wdata_valid ? io_banks_56_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51345.6]
  assign _GEN_56 = _T_1194 ? _T_1195 : regs_56; // @[SRAM.scala 148:48:@51344.4]
  assign _T_1201 = io_waddr == 6'h39; // @[SRAM.scala 148:37:@51352.4]
  assign _T_1202 = io_wen & _T_1201; // @[SRAM.scala 148:25:@51353.4]
  assign _T_1203 = io_banks_57_wdata_valid | _T_1202; // @[SRAM.scala 148:15:@51354.4]
  assign _T_1204 = io_banks_57_wdata_valid ? io_banks_57_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51356.6]
  assign _GEN_57 = _T_1203 ? _T_1204 : regs_57; // @[SRAM.scala 148:48:@51355.4]
  assign _T_1210 = io_waddr == 6'h3a; // @[SRAM.scala 148:37:@51363.4]
  assign _T_1211 = io_wen & _T_1210; // @[SRAM.scala 148:25:@51364.4]
  assign _T_1212 = io_banks_58_wdata_valid | _T_1211; // @[SRAM.scala 148:15:@51365.4]
  assign _T_1213 = io_banks_58_wdata_valid ? io_banks_58_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51367.6]
  assign _GEN_58 = _T_1212 ? _T_1213 : regs_58; // @[SRAM.scala 148:48:@51366.4]
  assign _T_1219 = io_waddr == 6'h3b; // @[SRAM.scala 148:37:@51374.4]
  assign _T_1220 = io_wen & _T_1219; // @[SRAM.scala 148:25:@51375.4]
  assign _T_1221 = io_banks_59_wdata_valid | _T_1220; // @[SRAM.scala 148:15:@51376.4]
  assign _T_1222 = io_banks_59_wdata_valid ? io_banks_59_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51378.6]
  assign _GEN_59 = _T_1221 ? _T_1222 : regs_59; // @[SRAM.scala 148:48:@51377.4]
  assign _T_1228 = io_waddr == 6'h3c; // @[SRAM.scala 148:37:@51385.4]
  assign _T_1229 = io_wen & _T_1228; // @[SRAM.scala 148:25:@51386.4]
  assign _T_1230 = io_banks_60_wdata_valid | _T_1229; // @[SRAM.scala 148:15:@51387.4]
  assign _T_1231 = io_banks_60_wdata_valid ? io_banks_60_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51389.6]
  assign _GEN_60 = _T_1230 ? _T_1231 : regs_60; // @[SRAM.scala 148:48:@51388.4]
  assign _T_1237 = io_waddr == 6'h3d; // @[SRAM.scala 148:37:@51396.4]
  assign _T_1238 = io_wen & _T_1237; // @[SRAM.scala 148:25:@51397.4]
  assign _T_1239 = io_banks_61_wdata_valid | _T_1238; // @[SRAM.scala 148:15:@51398.4]
  assign _T_1240 = io_banks_61_wdata_valid ? io_banks_61_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51400.6]
  assign _GEN_61 = _T_1239 ? _T_1240 : regs_61; // @[SRAM.scala 148:48:@51399.4]
  assign _T_1246 = io_waddr == 6'h3e; // @[SRAM.scala 148:37:@51407.4]
  assign _T_1247 = io_wen & _T_1246; // @[SRAM.scala 148:25:@51408.4]
  assign _T_1248 = io_banks_62_wdata_valid | _T_1247; // @[SRAM.scala 148:15:@51409.4]
  assign _T_1249 = io_banks_62_wdata_valid ? io_banks_62_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51411.6]
  assign _GEN_62 = _T_1248 ? _T_1249 : regs_62; // @[SRAM.scala 148:48:@51410.4]
  assign _T_1255 = io_waddr == 6'h3f; // @[SRAM.scala 148:37:@51418.4]
  assign _T_1256 = io_wen & _T_1255; // @[SRAM.scala 148:25:@51419.4]
  assign _T_1257 = io_banks_63_wdata_valid | _T_1256; // @[SRAM.scala 148:15:@51420.4]
  assign _T_1258 = io_banks_63_wdata_valid ? io_banks_63_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@51422.6]
  assign _GEN_63 = _T_1257 ? _T_1258 : regs_63; // @[SRAM.scala 148:48:@51421.4]
  assign _GEN_65 = 6'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_66 = 6'h2 == io_raddr ? regs_2 : _GEN_65; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_67 = 6'h3 == io_raddr ? regs_3 : _GEN_66; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_68 = 6'h4 == io_raddr ? regs_4 : _GEN_67; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_69 = 6'h5 == io_raddr ? regs_5 : _GEN_68; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_70 = 6'h6 == io_raddr ? regs_6 : _GEN_69; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_71 = 6'h7 == io_raddr ? regs_7 : _GEN_70; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_72 = 6'h8 == io_raddr ? regs_8 : _GEN_71; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_73 = 6'h9 == io_raddr ? regs_9 : _GEN_72; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_74 = 6'ha == io_raddr ? regs_10 : _GEN_73; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_75 = 6'hb == io_raddr ? regs_11 : _GEN_74; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_76 = 6'hc == io_raddr ? regs_12 : _GEN_75; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_77 = 6'hd == io_raddr ? regs_13 : _GEN_76; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_78 = 6'he == io_raddr ? regs_14 : _GEN_77; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_79 = 6'hf == io_raddr ? regs_15 : _GEN_78; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_80 = 6'h10 == io_raddr ? regs_16 : _GEN_79; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_81 = 6'h11 == io_raddr ? regs_17 : _GEN_80; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_82 = 6'h12 == io_raddr ? regs_18 : _GEN_81; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_83 = 6'h13 == io_raddr ? regs_19 : _GEN_82; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_84 = 6'h14 == io_raddr ? regs_20 : _GEN_83; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_85 = 6'h15 == io_raddr ? regs_21 : _GEN_84; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_86 = 6'h16 == io_raddr ? regs_22 : _GEN_85; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_87 = 6'h17 == io_raddr ? regs_23 : _GEN_86; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_88 = 6'h18 == io_raddr ? regs_24 : _GEN_87; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_89 = 6'h19 == io_raddr ? regs_25 : _GEN_88; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_90 = 6'h1a == io_raddr ? regs_26 : _GEN_89; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_91 = 6'h1b == io_raddr ? regs_27 : _GEN_90; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_92 = 6'h1c == io_raddr ? regs_28 : _GEN_91; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_93 = 6'h1d == io_raddr ? regs_29 : _GEN_92; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_94 = 6'h1e == io_raddr ? regs_30 : _GEN_93; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_95 = 6'h1f == io_raddr ? regs_31 : _GEN_94; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_96 = 6'h20 == io_raddr ? regs_32 : _GEN_95; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_97 = 6'h21 == io_raddr ? regs_33 : _GEN_96; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_98 = 6'h22 == io_raddr ? regs_34 : _GEN_97; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_99 = 6'h23 == io_raddr ? regs_35 : _GEN_98; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_100 = 6'h24 == io_raddr ? regs_36 : _GEN_99; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_101 = 6'h25 == io_raddr ? regs_37 : _GEN_100; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_102 = 6'h26 == io_raddr ? regs_38 : _GEN_101; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_103 = 6'h27 == io_raddr ? regs_39 : _GEN_102; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_104 = 6'h28 == io_raddr ? regs_40 : _GEN_103; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_105 = 6'h29 == io_raddr ? regs_41 : _GEN_104; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_106 = 6'h2a == io_raddr ? regs_42 : _GEN_105; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_107 = 6'h2b == io_raddr ? regs_43 : _GEN_106; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_108 = 6'h2c == io_raddr ? regs_44 : _GEN_107; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_109 = 6'h2d == io_raddr ? regs_45 : _GEN_108; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_110 = 6'h2e == io_raddr ? regs_46 : _GEN_109; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_111 = 6'h2f == io_raddr ? regs_47 : _GEN_110; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_112 = 6'h30 == io_raddr ? regs_48 : _GEN_111; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_113 = 6'h31 == io_raddr ? regs_49 : _GEN_112; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_114 = 6'h32 == io_raddr ? regs_50 : _GEN_113; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_115 = 6'h33 == io_raddr ? regs_51 : _GEN_114; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_116 = 6'h34 == io_raddr ? regs_52 : _GEN_115; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_117 = 6'h35 == io_raddr ? regs_53 : _GEN_116; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_118 = 6'h36 == io_raddr ? regs_54 : _GEN_117; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_119 = 6'h37 == io_raddr ? regs_55 : _GEN_118; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_120 = 6'h38 == io_raddr ? regs_56 : _GEN_119; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_121 = 6'h39 == io_raddr ? regs_57 : _GEN_120; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_122 = 6'h3a == io_raddr ? regs_58 : _GEN_121; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_123 = 6'h3b == io_raddr ? regs_59 : _GEN_122; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_124 = 6'h3c == io_raddr ? regs_60 : _GEN_123; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_125 = 6'h3d == io_raddr ? regs_61 : _GEN_124; // @[SRAM.scala 155:12:@51491.4]
  assign _GEN_126 = 6'h3e == io_raddr ? regs_62 : _GEN_125; // @[SRAM.scala 155:12:@51491.4]
  assign io_rdata = 6'h3f == io_raddr ? regs_63 : _GEN_126; // @[SRAM.scala 155:12:@51491.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_690) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_699) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_708) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_717) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_4 <= 1'h0;
    end else begin
      if (_T_726) begin
        if (io_banks_4_wdata_valid) begin
          regs_4 <= io_banks_4_wdata_bits;
        end else begin
          regs_4 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_5 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (io_banks_5_wdata_valid) begin
          regs_5 <= io_banks_5_wdata_bits;
        end else begin
          regs_5 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_6 <= 1'h0;
    end else begin
      if (_T_744) begin
        if (io_banks_6_wdata_valid) begin
          regs_6 <= io_banks_6_wdata_bits;
        end else begin
          regs_6 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_7 <= 1'h0;
    end else begin
      if (_T_753) begin
        if (io_banks_7_wdata_valid) begin
          regs_7 <= io_banks_7_wdata_bits;
        end else begin
          regs_7 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_8 <= 1'h0;
    end else begin
      if (_T_762) begin
        if (io_banks_8_wdata_valid) begin
          regs_8 <= io_banks_8_wdata_bits;
        end else begin
          regs_8 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_9 <= 1'h0;
    end else begin
      if (_T_771) begin
        if (io_banks_9_wdata_valid) begin
          regs_9 <= io_banks_9_wdata_bits;
        end else begin
          regs_9 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_10 <= 1'h0;
    end else begin
      if (_T_780) begin
        if (io_banks_10_wdata_valid) begin
          regs_10 <= io_banks_10_wdata_bits;
        end else begin
          regs_10 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_11 <= 1'h0;
    end else begin
      if (_T_789) begin
        if (io_banks_11_wdata_valid) begin
          regs_11 <= io_banks_11_wdata_bits;
        end else begin
          regs_11 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_12 <= 1'h0;
    end else begin
      if (_T_798) begin
        if (io_banks_12_wdata_valid) begin
          regs_12 <= io_banks_12_wdata_bits;
        end else begin
          regs_12 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_13 <= 1'h0;
    end else begin
      if (_T_807) begin
        if (io_banks_13_wdata_valid) begin
          regs_13 <= io_banks_13_wdata_bits;
        end else begin
          regs_13 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_14 <= 1'h0;
    end else begin
      if (_T_816) begin
        if (io_banks_14_wdata_valid) begin
          regs_14 <= io_banks_14_wdata_bits;
        end else begin
          regs_14 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_15 <= 1'h0;
    end else begin
      if (_T_825) begin
        if (io_banks_15_wdata_valid) begin
          regs_15 <= io_banks_15_wdata_bits;
        end else begin
          regs_15 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_16 <= 1'h0;
    end else begin
      if (_T_834) begin
        if (io_banks_16_wdata_valid) begin
          regs_16 <= io_banks_16_wdata_bits;
        end else begin
          regs_16 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_17 <= 1'h0;
    end else begin
      if (_T_843) begin
        if (io_banks_17_wdata_valid) begin
          regs_17 <= io_banks_17_wdata_bits;
        end else begin
          regs_17 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_18 <= 1'h0;
    end else begin
      if (_T_852) begin
        if (io_banks_18_wdata_valid) begin
          regs_18 <= io_banks_18_wdata_bits;
        end else begin
          regs_18 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_19 <= 1'h0;
    end else begin
      if (_T_861) begin
        if (io_banks_19_wdata_valid) begin
          regs_19 <= io_banks_19_wdata_bits;
        end else begin
          regs_19 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_20 <= 1'h0;
    end else begin
      if (_T_870) begin
        if (io_banks_20_wdata_valid) begin
          regs_20 <= io_banks_20_wdata_bits;
        end else begin
          regs_20 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_21 <= 1'h0;
    end else begin
      if (_T_879) begin
        if (io_banks_21_wdata_valid) begin
          regs_21 <= io_banks_21_wdata_bits;
        end else begin
          regs_21 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_22 <= 1'h0;
    end else begin
      if (_T_888) begin
        if (io_banks_22_wdata_valid) begin
          regs_22 <= io_banks_22_wdata_bits;
        end else begin
          regs_22 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_23 <= 1'h0;
    end else begin
      if (_T_897) begin
        if (io_banks_23_wdata_valid) begin
          regs_23 <= io_banks_23_wdata_bits;
        end else begin
          regs_23 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_24 <= 1'h0;
    end else begin
      if (_T_906) begin
        if (io_banks_24_wdata_valid) begin
          regs_24 <= io_banks_24_wdata_bits;
        end else begin
          regs_24 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_25 <= 1'h0;
    end else begin
      if (_T_915) begin
        if (io_banks_25_wdata_valid) begin
          regs_25 <= io_banks_25_wdata_bits;
        end else begin
          regs_25 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_26 <= 1'h0;
    end else begin
      if (_T_924) begin
        if (io_banks_26_wdata_valid) begin
          regs_26 <= io_banks_26_wdata_bits;
        end else begin
          regs_26 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_27 <= 1'h0;
    end else begin
      if (_T_933) begin
        if (io_banks_27_wdata_valid) begin
          regs_27 <= io_banks_27_wdata_bits;
        end else begin
          regs_27 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_28 <= 1'h0;
    end else begin
      if (_T_942) begin
        if (io_banks_28_wdata_valid) begin
          regs_28 <= io_banks_28_wdata_bits;
        end else begin
          regs_28 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_29 <= 1'h0;
    end else begin
      if (_T_951) begin
        if (io_banks_29_wdata_valid) begin
          regs_29 <= io_banks_29_wdata_bits;
        end else begin
          regs_29 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_30 <= 1'h0;
    end else begin
      if (_T_960) begin
        if (io_banks_30_wdata_valid) begin
          regs_30 <= io_banks_30_wdata_bits;
        end else begin
          regs_30 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_31 <= 1'h0;
    end else begin
      if (_T_969) begin
        if (io_banks_31_wdata_valid) begin
          regs_31 <= io_banks_31_wdata_bits;
        end else begin
          regs_31 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_32 <= 1'h0;
    end else begin
      if (_T_978) begin
        if (io_banks_32_wdata_valid) begin
          regs_32 <= io_banks_32_wdata_bits;
        end else begin
          regs_32 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_33 <= 1'h0;
    end else begin
      if (_T_987) begin
        if (io_banks_33_wdata_valid) begin
          regs_33 <= io_banks_33_wdata_bits;
        end else begin
          regs_33 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_34 <= 1'h0;
    end else begin
      if (_T_996) begin
        if (io_banks_34_wdata_valid) begin
          regs_34 <= io_banks_34_wdata_bits;
        end else begin
          regs_34 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_35 <= 1'h0;
    end else begin
      if (_T_1005) begin
        if (io_banks_35_wdata_valid) begin
          regs_35 <= io_banks_35_wdata_bits;
        end else begin
          regs_35 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_36 <= 1'h0;
    end else begin
      if (_T_1014) begin
        if (io_banks_36_wdata_valid) begin
          regs_36 <= io_banks_36_wdata_bits;
        end else begin
          regs_36 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_37 <= 1'h0;
    end else begin
      if (_T_1023) begin
        if (io_banks_37_wdata_valid) begin
          regs_37 <= io_banks_37_wdata_bits;
        end else begin
          regs_37 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_38 <= 1'h0;
    end else begin
      if (_T_1032) begin
        if (io_banks_38_wdata_valid) begin
          regs_38 <= io_banks_38_wdata_bits;
        end else begin
          regs_38 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_39 <= 1'h0;
    end else begin
      if (_T_1041) begin
        if (io_banks_39_wdata_valid) begin
          regs_39 <= io_banks_39_wdata_bits;
        end else begin
          regs_39 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_40 <= 1'h0;
    end else begin
      if (_T_1050) begin
        if (io_banks_40_wdata_valid) begin
          regs_40 <= io_banks_40_wdata_bits;
        end else begin
          regs_40 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_41 <= 1'h0;
    end else begin
      if (_T_1059) begin
        if (io_banks_41_wdata_valid) begin
          regs_41 <= io_banks_41_wdata_bits;
        end else begin
          regs_41 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_42 <= 1'h0;
    end else begin
      if (_T_1068) begin
        if (io_banks_42_wdata_valid) begin
          regs_42 <= io_banks_42_wdata_bits;
        end else begin
          regs_42 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_43 <= 1'h0;
    end else begin
      if (_T_1077) begin
        if (io_banks_43_wdata_valid) begin
          regs_43 <= io_banks_43_wdata_bits;
        end else begin
          regs_43 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_44 <= 1'h0;
    end else begin
      if (_T_1086) begin
        if (io_banks_44_wdata_valid) begin
          regs_44 <= io_banks_44_wdata_bits;
        end else begin
          regs_44 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_45 <= 1'h0;
    end else begin
      if (_T_1095) begin
        if (io_banks_45_wdata_valid) begin
          regs_45 <= io_banks_45_wdata_bits;
        end else begin
          regs_45 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_46 <= 1'h0;
    end else begin
      if (_T_1104) begin
        if (io_banks_46_wdata_valid) begin
          regs_46 <= io_banks_46_wdata_bits;
        end else begin
          regs_46 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_47 <= 1'h0;
    end else begin
      if (_T_1113) begin
        if (io_banks_47_wdata_valid) begin
          regs_47 <= io_banks_47_wdata_bits;
        end else begin
          regs_47 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_48 <= 1'h0;
    end else begin
      if (_T_1122) begin
        if (io_banks_48_wdata_valid) begin
          regs_48 <= io_banks_48_wdata_bits;
        end else begin
          regs_48 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_49 <= 1'h0;
    end else begin
      if (_T_1131) begin
        if (io_banks_49_wdata_valid) begin
          regs_49 <= io_banks_49_wdata_bits;
        end else begin
          regs_49 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_50 <= 1'h0;
    end else begin
      if (_T_1140) begin
        if (io_banks_50_wdata_valid) begin
          regs_50 <= io_banks_50_wdata_bits;
        end else begin
          regs_50 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_51 <= 1'h0;
    end else begin
      if (_T_1149) begin
        if (io_banks_51_wdata_valid) begin
          regs_51 <= io_banks_51_wdata_bits;
        end else begin
          regs_51 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_52 <= 1'h0;
    end else begin
      if (_T_1158) begin
        if (io_banks_52_wdata_valid) begin
          regs_52 <= io_banks_52_wdata_bits;
        end else begin
          regs_52 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_53 <= 1'h0;
    end else begin
      if (_T_1167) begin
        if (io_banks_53_wdata_valid) begin
          regs_53 <= io_banks_53_wdata_bits;
        end else begin
          regs_53 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_54 <= 1'h0;
    end else begin
      if (_T_1176) begin
        if (io_banks_54_wdata_valid) begin
          regs_54 <= io_banks_54_wdata_bits;
        end else begin
          regs_54 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_55 <= 1'h0;
    end else begin
      if (_T_1185) begin
        if (io_banks_55_wdata_valid) begin
          regs_55 <= io_banks_55_wdata_bits;
        end else begin
          regs_55 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_56 <= 1'h0;
    end else begin
      if (_T_1194) begin
        if (io_banks_56_wdata_valid) begin
          regs_56 <= io_banks_56_wdata_bits;
        end else begin
          regs_56 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_57 <= 1'h0;
    end else begin
      if (_T_1203) begin
        if (io_banks_57_wdata_valid) begin
          regs_57 <= io_banks_57_wdata_bits;
        end else begin
          regs_57 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_58 <= 1'h0;
    end else begin
      if (_T_1212) begin
        if (io_banks_58_wdata_valid) begin
          regs_58 <= io_banks_58_wdata_bits;
        end else begin
          regs_58 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_59 <= 1'h0;
    end else begin
      if (_T_1221) begin
        if (io_banks_59_wdata_valid) begin
          regs_59 <= io_banks_59_wdata_bits;
        end else begin
          regs_59 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_60 <= 1'h0;
    end else begin
      if (_T_1230) begin
        if (io_banks_60_wdata_valid) begin
          regs_60 <= io_banks_60_wdata_bits;
        end else begin
          regs_60 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_61 <= 1'h0;
    end else begin
      if (_T_1239) begin
        if (io_banks_61_wdata_valid) begin
          regs_61 <= io_banks_61_wdata_bits;
        end else begin
          regs_61 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_62 <= 1'h0;
    end else begin
      if (_T_1248) begin
        if (io_banks_62_wdata_valid) begin
          regs_62 <= io_banks_62_wdata_bits;
        end else begin
          regs_62 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_63 <= 1'h0;
    end else begin
      if (_T_1257) begin
        if (io_banks_63_wdata_valid) begin
          regs_63 <= io_banks_63_wdata_bits;
        end else begin
          regs_63 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_33( // @[:@51493.2]
  input   clock, // @[:@51494.4]
  input   reset, // @[:@51495.4]
  output  io_in_ready, // @[:@51496.4]
  input   io_in_valid, // @[:@51496.4]
  input   io_in_bits, // @[:@51496.4]
  input   io_out_ready, // @[:@51496.4]
  output  io_out_valid, // @[:@51496.4]
  output  io_out_bits, // @[:@51496.4]
  input   io_banks_0_wdata_valid, // @[:@51496.4]
  input   io_banks_0_wdata_bits, // @[:@51496.4]
  input   io_banks_1_wdata_valid, // @[:@51496.4]
  input   io_banks_1_wdata_bits, // @[:@51496.4]
  input   io_banks_2_wdata_valid, // @[:@51496.4]
  input   io_banks_2_wdata_bits, // @[:@51496.4]
  input   io_banks_3_wdata_valid, // @[:@51496.4]
  input   io_banks_3_wdata_bits, // @[:@51496.4]
  input   io_banks_4_wdata_valid, // @[:@51496.4]
  input   io_banks_4_wdata_bits, // @[:@51496.4]
  input   io_banks_5_wdata_valid, // @[:@51496.4]
  input   io_banks_5_wdata_bits, // @[:@51496.4]
  input   io_banks_6_wdata_valid, // @[:@51496.4]
  input   io_banks_6_wdata_bits, // @[:@51496.4]
  input   io_banks_7_wdata_valid, // @[:@51496.4]
  input   io_banks_7_wdata_bits, // @[:@51496.4]
  input   io_banks_8_wdata_valid, // @[:@51496.4]
  input   io_banks_8_wdata_bits, // @[:@51496.4]
  input   io_banks_9_wdata_valid, // @[:@51496.4]
  input   io_banks_9_wdata_bits, // @[:@51496.4]
  input   io_banks_10_wdata_valid, // @[:@51496.4]
  input   io_banks_10_wdata_bits, // @[:@51496.4]
  input   io_banks_11_wdata_valid, // @[:@51496.4]
  input   io_banks_11_wdata_bits, // @[:@51496.4]
  input   io_banks_12_wdata_valid, // @[:@51496.4]
  input   io_banks_12_wdata_bits, // @[:@51496.4]
  input   io_banks_13_wdata_valid, // @[:@51496.4]
  input   io_banks_13_wdata_bits, // @[:@51496.4]
  input   io_banks_14_wdata_valid, // @[:@51496.4]
  input   io_banks_14_wdata_bits, // @[:@51496.4]
  input   io_banks_15_wdata_valid, // @[:@51496.4]
  input   io_banks_15_wdata_bits, // @[:@51496.4]
  input   io_banks_16_wdata_valid, // @[:@51496.4]
  input   io_banks_16_wdata_bits, // @[:@51496.4]
  input   io_banks_17_wdata_valid, // @[:@51496.4]
  input   io_banks_17_wdata_bits, // @[:@51496.4]
  input   io_banks_18_wdata_valid, // @[:@51496.4]
  input   io_banks_18_wdata_bits, // @[:@51496.4]
  input   io_banks_19_wdata_valid, // @[:@51496.4]
  input   io_banks_19_wdata_bits, // @[:@51496.4]
  input   io_banks_20_wdata_valid, // @[:@51496.4]
  input   io_banks_20_wdata_bits, // @[:@51496.4]
  input   io_banks_21_wdata_valid, // @[:@51496.4]
  input   io_banks_21_wdata_bits, // @[:@51496.4]
  input   io_banks_22_wdata_valid, // @[:@51496.4]
  input   io_banks_22_wdata_bits, // @[:@51496.4]
  input   io_banks_23_wdata_valid, // @[:@51496.4]
  input   io_banks_23_wdata_bits, // @[:@51496.4]
  input   io_banks_24_wdata_valid, // @[:@51496.4]
  input   io_banks_24_wdata_bits, // @[:@51496.4]
  input   io_banks_25_wdata_valid, // @[:@51496.4]
  input   io_banks_25_wdata_bits, // @[:@51496.4]
  input   io_banks_26_wdata_valid, // @[:@51496.4]
  input   io_banks_26_wdata_bits, // @[:@51496.4]
  input   io_banks_27_wdata_valid, // @[:@51496.4]
  input   io_banks_27_wdata_bits, // @[:@51496.4]
  input   io_banks_28_wdata_valid, // @[:@51496.4]
  input   io_banks_28_wdata_bits, // @[:@51496.4]
  input   io_banks_29_wdata_valid, // @[:@51496.4]
  input   io_banks_29_wdata_bits, // @[:@51496.4]
  input   io_banks_30_wdata_valid, // @[:@51496.4]
  input   io_banks_30_wdata_bits, // @[:@51496.4]
  input   io_banks_31_wdata_valid, // @[:@51496.4]
  input   io_banks_31_wdata_bits, // @[:@51496.4]
  input   io_banks_32_wdata_valid, // @[:@51496.4]
  input   io_banks_32_wdata_bits, // @[:@51496.4]
  input   io_banks_33_wdata_valid, // @[:@51496.4]
  input   io_banks_33_wdata_bits, // @[:@51496.4]
  input   io_banks_34_wdata_valid, // @[:@51496.4]
  input   io_banks_34_wdata_bits, // @[:@51496.4]
  input   io_banks_35_wdata_valid, // @[:@51496.4]
  input   io_banks_35_wdata_bits, // @[:@51496.4]
  input   io_banks_36_wdata_valid, // @[:@51496.4]
  input   io_banks_36_wdata_bits, // @[:@51496.4]
  input   io_banks_37_wdata_valid, // @[:@51496.4]
  input   io_banks_37_wdata_bits, // @[:@51496.4]
  input   io_banks_38_wdata_valid, // @[:@51496.4]
  input   io_banks_38_wdata_bits, // @[:@51496.4]
  input   io_banks_39_wdata_valid, // @[:@51496.4]
  input   io_banks_39_wdata_bits, // @[:@51496.4]
  input   io_banks_40_wdata_valid, // @[:@51496.4]
  input   io_banks_40_wdata_bits, // @[:@51496.4]
  input   io_banks_41_wdata_valid, // @[:@51496.4]
  input   io_banks_41_wdata_bits, // @[:@51496.4]
  input   io_banks_42_wdata_valid, // @[:@51496.4]
  input   io_banks_42_wdata_bits, // @[:@51496.4]
  input   io_banks_43_wdata_valid, // @[:@51496.4]
  input   io_banks_43_wdata_bits, // @[:@51496.4]
  input   io_banks_44_wdata_valid, // @[:@51496.4]
  input   io_banks_44_wdata_bits, // @[:@51496.4]
  input   io_banks_45_wdata_valid, // @[:@51496.4]
  input   io_banks_45_wdata_bits, // @[:@51496.4]
  input   io_banks_46_wdata_valid, // @[:@51496.4]
  input   io_banks_46_wdata_bits, // @[:@51496.4]
  input   io_banks_47_wdata_valid, // @[:@51496.4]
  input   io_banks_47_wdata_bits, // @[:@51496.4]
  input   io_banks_48_wdata_valid, // @[:@51496.4]
  input   io_banks_48_wdata_bits, // @[:@51496.4]
  input   io_banks_49_wdata_valid, // @[:@51496.4]
  input   io_banks_49_wdata_bits, // @[:@51496.4]
  input   io_banks_50_wdata_valid, // @[:@51496.4]
  input   io_banks_50_wdata_bits, // @[:@51496.4]
  input   io_banks_51_wdata_valid, // @[:@51496.4]
  input   io_banks_51_wdata_bits, // @[:@51496.4]
  input   io_banks_52_wdata_valid, // @[:@51496.4]
  input   io_banks_52_wdata_bits, // @[:@51496.4]
  input   io_banks_53_wdata_valid, // @[:@51496.4]
  input   io_banks_53_wdata_bits, // @[:@51496.4]
  input   io_banks_54_wdata_valid, // @[:@51496.4]
  input   io_banks_54_wdata_bits, // @[:@51496.4]
  input   io_banks_55_wdata_valid, // @[:@51496.4]
  input   io_banks_55_wdata_bits, // @[:@51496.4]
  input   io_banks_56_wdata_valid, // @[:@51496.4]
  input   io_banks_56_wdata_bits, // @[:@51496.4]
  input   io_banks_57_wdata_valid, // @[:@51496.4]
  input   io_banks_57_wdata_bits, // @[:@51496.4]
  input   io_banks_58_wdata_valid, // @[:@51496.4]
  input   io_banks_58_wdata_bits, // @[:@51496.4]
  input   io_banks_59_wdata_valid, // @[:@51496.4]
  input   io_banks_59_wdata_bits, // @[:@51496.4]
  input   io_banks_60_wdata_valid, // @[:@51496.4]
  input   io_banks_60_wdata_bits, // @[:@51496.4]
  input   io_banks_61_wdata_valid, // @[:@51496.4]
  input   io_banks_61_wdata_bits, // @[:@51496.4]
  input   io_banks_62_wdata_valid, // @[:@51496.4]
  input   io_banks_62_wdata_bits, // @[:@51496.4]
  input   io_banks_63_wdata_valid, // @[:@51496.4]
  input   io_banks_63_wdata_bits // @[:@51496.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@51762.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@51762.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@51762.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@51762.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@51762.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@51772.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@51772.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@51772.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@51772.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@51772.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@51787.4]
  wire [5:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@51787.4]
  wire [5:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_4_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_4_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_5_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_5_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_6_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_6_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_7_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_7_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_8_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_8_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_9_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_9_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_10_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_10_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_11_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_11_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_12_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_12_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_13_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_13_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_14_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_14_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_15_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_15_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_16_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_16_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_17_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_17_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_18_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_18_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_19_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_19_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_20_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_20_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_21_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_21_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_22_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_22_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_23_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_23_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_24_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_24_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_25_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_25_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_26_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_26_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_27_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_27_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_28_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_28_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_29_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_29_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_30_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_30_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_31_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_31_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_32_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_32_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_33_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_33_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_34_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_34_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_35_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_35_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_36_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_36_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_37_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_37_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_38_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_38_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_39_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_39_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_40_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_40_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_41_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_41_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_42_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_42_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_43_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_43_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_44_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_44_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_45_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_45_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_46_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_46_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_47_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_47_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_48_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_48_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_49_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_49_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_50_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_50_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_51_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_51_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_52_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_52_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_53_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_53_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_54_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_54_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_55_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_55_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_56_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_56_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_57_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_57_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_58_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_58_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_59_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_59_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_60_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_60_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_61_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_61_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_62_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_62_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_63_wdata_valid; // @[FIFO.scala 49:19:@51787.4]
  wire  FFRAM_io_banks_63_wdata_bits; // @[FIFO.scala 49:19:@51787.4]
  wire  writeEn; // @[FIFO.scala 30:29:@51760.4]
  wire  readEn; // @[FIFO.scala 31:29:@51761.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@51782.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@51783.4]
  wire  _T_824; // @[FIFO.scala 45:27:@51784.4]
  wire  empty; // @[FIFO.scala 45:24:@51785.4]
  wire  full; // @[FIFO.scala 46:23:@51786.4]
  wire  _T_1657; // @[FIFO.scala 83:17:@52953.4]
  wire  _GEN_64; // @[FIFO.scala 83:29:@52954.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@51762.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@51772.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM_16 FFRAM ( // @[FIFO.scala 49:19:@51787.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(FFRAM_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(FFRAM_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(FFRAM_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(FFRAM_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(FFRAM_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(FFRAM_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(FFRAM_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(FFRAM_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(FFRAM_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(FFRAM_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(FFRAM_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(FFRAM_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(FFRAM_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(FFRAM_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(FFRAM_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(FFRAM_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(FFRAM_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(FFRAM_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(FFRAM_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(FFRAM_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(FFRAM_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(FFRAM_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(FFRAM_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(FFRAM_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(FFRAM_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(FFRAM_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(FFRAM_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(FFRAM_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(FFRAM_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(FFRAM_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(FFRAM_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(FFRAM_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(FFRAM_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(FFRAM_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(FFRAM_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(FFRAM_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(FFRAM_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(FFRAM_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(FFRAM_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(FFRAM_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(FFRAM_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(FFRAM_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(FFRAM_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(FFRAM_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(FFRAM_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(FFRAM_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(FFRAM_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(FFRAM_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(FFRAM_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(FFRAM_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(FFRAM_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(FFRAM_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(FFRAM_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(FFRAM_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(FFRAM_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(FFRAM_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(FFRAM_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(FFRAM_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(FFRAM_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(FFRAM_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(FFRAM_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(FFRAM_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(FFRAM_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(FFRAM_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(FFRAM_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(FFRAM_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(FFRAM_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(FFRAM_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(FFRAM_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(FFRAM_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(FFRAM_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(FFRAM_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(FFRAM_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(FFRAM_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(FFRAM_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(FFRAM_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(FFRAM_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(FFRAM_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(FFRAM_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(FFRAM_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(FFRAM_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(FFRAM_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(FFRAM_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(FFRAM_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(FFRAM_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(FFRAM_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(FFRAM_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(FFRAM_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(FFRAM_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(FFRAM_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(FFRAM_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(FFRAM_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(FFRAM_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(FFRAM_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(FFRAM_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(FFRAM_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(FFRAM_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(FFRAM_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(FFRAM_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(FFRAM_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(FFRAM_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(FFRAM_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(FFRAM_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(FFRAM_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(FFRAM_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(FFRAM_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(FFRAM_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(FFRAM_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(FFRAM_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(FFRAM_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(FFRAM_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(FFRAM_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(FFRAM_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(FFRAM_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(FFRAM_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(FFRAM_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(FFRAM_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(FFRAM_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(FFRAM_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(FFRAM_io_banks_63_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@51760.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@51761.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@51783.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@51784.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@51785.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@51786.4]
  assign _T_1657 = writeEn != readEn; // @[FIFO.scala 83:17:@52953.4]
  assign _GEN_64 = _T_1657 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@52954.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@52960.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@52958.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@51992.4]
  assign enqCounter_clock = clock; // @[:@51763.4]
  assign enqCounter_reset = reset; // @[:@51764.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@51770.4]
  assign deqCounter_clock = clock; // @[:@51773.4]
  assign deqCounter_reset = reset; // @[:@51774.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@51780.4]
  assign FFRAM_clock = clock; // @[:@51788.4]
  assign FFRAM_reset = reset; // @[:@51789.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@51988.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@51989.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@51990.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@51991.4]
  assign FFRAM_io_banks_0_wdata_valid = io_banks_0_wdata_valid; // @[FIFO.scala 59:15:@51994.4]
  assign FFRAM_io_banks_0_wdata_bits = io_banks_0_wdata_bits; // @[FIFO.scala 59:15:@51993.4]
  assign FFRAM_io_banks_1_wdata_valid = io_banks_1_wdata_valid; // @[FIFO.scala 59:15:@51997.4]
  assign FFRAM_io_banks_1_wdata_bits = io_banks_1_wdata_bits; // @[FIFO.scala 59:15:@51996.4]
  assign FFRAM_io_banks_2_wdata_valid = io_banks_2_wdata_valid; // @[FIFO.scala 59:15:@52000.4]
  assign FFRAM_io_banks_2_wdata_bits = io_banks_2_wdata_bits; // @[FIFO.scala 59:15:@51999.4]
  assign FFRAM_io_banks_3_wdata_valid = io_banks_3_wdata_valid; // @[FIFO.scala 59:15:@52003.4]
  assign FFRAM_io_banks_3_wdata_bits = io_banks_3_wdata_bits; // @[FIFO.scala 59:15:@52002.4]
  assign FFRAM_io_banks_4_wdata_valid = io_banks_4_wdata_valid; // @[FIFO.scala 59:15:@52006.4]
  assign FFRAM_io_banks_4_wdata_bits = io_banks_4_wdata_bits; // @[FIFO.scala 59:15:@52005.4]
  assign FFRAM_io_banks_5_wdata_valid = io_banks_5_wdata_valid; // @[FIFO.scala 59:15:@52009.4]
  assign FFRAM_io_banks_5_wdata_bits = io_banks_5_wdata_bits; // @[FIFO.scala 59:15:@52008.4]
  assign FFRAM_io_banks_6_wdata_valid = io_banks_6_wdata_valid; // @[FIFO.scala 59:15:@52012.4]
  assign FFRAM_io_banks_6_wdata_bits = io_banks_6_wdata_bits; // @[FIFO.scala 59:15:@52011.4]
  assign FFRAM_io_banks_7_wdata_valid = io_banks_7_wdata_valid; // @[FIFO.scala 59:15:@52015.4]
  assign FFRAM_io_banks_7_wdata_bits = io_banks_7_wdata_bits; // @[FIFO.scala 59:15:@52014.4]
  assign FFRAM_io_banks_8_wdata_valid = io_banks_8_wdata_valid; // @[FIFO.scala 59:15:@52018.4]
  assign FFRAM_io_banks_8_wdata_bits = io_banks_8_wdata_bits; // @[FIFO.scala 59:15:@52017.4]
  assign FFRAM_io_banks_9_wdata_valid = io_banks_9_wdata_valid; // @[FIFO.scala 59:15:@52021.4]
  assign FFRAM_io_banks_9_wdata_bits = io_banks_9_wdata_bits; // @[FIFO.scala 59:15:@52020.4]
  assign FFRAM_io_banks_10_wdata_valid = io_banks_10_wdata_valid; // @[FIFO.scala 59:15:@52024.4]
  assign FFRAM_io_banks_10_wdata_bits = io_banks_10_wdata_bits; // @[FIFO.scala 59:15:@52023.4]
  assign FFRAM_io_banks_11_wdata_valid = io_banks_11_wdata_valid; // @[FIFO.scala 59:15:@52027.4]
  assign FFRAM_io_banks_11_wdata_bits = io_banks_11_wdata_bits; // @[FIFO.scala 59:15:@52026.4]
  assign FFRAM_io_banks_12_wdata_valid = io_banks_12_wdata_valid; // @[FIFO.scala 59:15:@52030.4]
  assign FFRAM_io_banks_12_wdata_bits = io_banks_12_wdata_bits; // @[FIFO.scala 59:15:@52029.4]
  assign FFRAM_io_banks_13_wdata_valid = io_banks_13_wdata_valid; // @[FIFO.scala 59:15:@52033.4]
  assign FFRAM_io_banks_13_wdata_bits = io_banks_13_wdata_bits; // @[FIFO.scala 59:15:@52032.4]
  assign FFRAM_io_banks_14_wdata_valid = io_banks_14_wdata_valid; // @[FIFO.scala 59:15:@52036.4]
  assign FFRAM_io_banks_14_wdata_bits = io_banks_14_wdata_bits; // @[FIFO.scala 59:15:@52035.4]
  assign FFRAM_io_banks_15_wdata_valid = io_banks_15_wdata_valid; // @[FIFO.scala 59:15:@52039.4]
  assign FFRAM_io_banks_15_wdata_bits = io_banks_15_wdata_bits; // @[FIFO.scala 59:15:@52038.4]
  assign FFRAM_io_banks_16_wdata_valid = io_banks_16_wdata_valid; // @[FIFO.scala 59:15:@52042.4]
  assign FFRAM_io_banks_16_wdata_bits = io_banks_16_wdata_bits; // @[FIFO.scala 59:15:@52041.4]
  assign FFRAM_io_banks_17_wdata_valid = io_banks_17_wdata_valid; // @[FIFO.scala 59:15:@52045.4]
  assign FFRAM_io_banks_17_wdata_bits = io_banks_17_wdata_bits; // @[FIFO.scala 59:15:@52044.4]
  assign FFRAM_io_banks_18_wdata_valid = io_banks_18_wdata_valid; // @[FIFO.scala 59:15:@52048.4]
  assign FFRAM_io_banks_18_wdata_bits = io_banks_18_wdata_bits; // @[FIFO.scala 59:15:@52047.4]
  assign FFRAM_io_banks_19_wdata_valid = io_banks_19_wdata_valid; // @[FIFO.scala 59:15:@52051.4]
  assign FFRAM_io_banks_19_wdata_bits = io_banks_19_wdata_bits; // @[FIFO.scala 59:15:@52050.4]
  assign FFRAM_io_banks_20_wdata_valid = io_banks_20_wdata_valid; // @[FIFO.scala 59:15:@52054.4]
  assign FFRAM_io_banks_20_wdata_bits = io_banks_20_wdata_bits; // @[FIFO.scala 59:15:@52053.4]
  assign FFRAM_io_banks_21_wdata_valid = io_banks_21_wdata_valid; // @[FIFO.scala 59:15:@52057.4]
  assign FFRAM_io_banks_21_wdata_bits = io_banks_21_wdata_bits; // @[FIFO.scala 59:15:@52056.4]
  assign FFRAM_io_banks_22_wdata_valid = io_banks_22_wdata_valid; // @[FIFO.scala 59:15:@52060.4]
  assign FFRAM_io_banks_22_wdata_bits = io_banks_22_wdata_bits; // @[FIFO.scala 59:15:@52059.4]
  assign FFRAM_io_banks_23_wdata_valid = io_banks_23_wdata_valid; // @[FIFO.scala 59:15:@52063.4]
  assign FFRAM_io_banks_23_wdata_bits = io_banks_23_wdata_bits; // @[FIFO.scala 59:15:@52062.4]
  assign FFRAM_io_banks_24_wdata_valid = io_banks_24_wdata_valid; // @[FIFO.scala 59:15:@52066.4]
  assign FFRAM_io_banks_24_wdata_bits = io_banks_24_wdata_bits; // @[FIFO.scala 59:15:@52065.4]
  assign FFRAM_io_banks_25_wdata_valid = io_banks_25_wdata_valid; // @[FIFO.scala 59:15:@52069.4]
  assign FFRAM_io_banks_25_wdata_bits = io_banks_25_wdata_bits; // @[FIFO.scala 59:15:@52068.4]
  assign FFRAM_io_banks_26_wdata_valid = io_banks_26_wdata_valid; // @[FIFO.scala 59:15:@52072.4]
  assign FFRAM_io_banks_26_wdata_bits = io_banks_26_wdata_bits; // @[FIFO.scala 59:15:@52071.4]
  assign FFRAM_io_banks_27_wdata_valid = io_banks_27_wdata_valid; // @[FIFO.scala 59:15:@52075.4]
  assign FFRAM_io_banks_27_wdata_bits = io_banks_27_wdata_bits; // @[FIFO.scala 59:15:@52074.4]
  assign FFRAM_io_banks_28_wdata_valid = io_banks_28_wdata_valid; // @[FIFO.scala 59:15:@52078.4]
  assign FFRAM_io_banks_28_wdata_bits = io_banks_28_wdata_bits; // @[FIFO.scala 59:15:@52077.4]
  assign FFRAM_io_banks_29_wdata_valid = io_banks_29_wdata_valid; // @[FIFO.scala 59:15:@52081.4]
  assign FFRAM_io_banks_29_wdata_bits = io_banks_29_wdata_bits; // @[FIFO.scala 59:15:@52080.4]
  assign FFRAM_io_banks_30_wdata_valid = io_banks_30_wdata_valid; // @[FIFO.scala 59:15:@52084.4]
  assign FFRAM_io_banks_30_wdata_bits = io_banks_30_wdata_bits; // @[FIFO.scala 59:15:@52083.4]
  assign FFRAM_io_banks_31_wdata_valid = io_banks_31_wdata_valid; // @[FIFO.scala 59:15:@52087.4]
  assign FFRAM_io_banks_31_wdata_bits = io_banks_31_wdata_bits; // @[FIFO.scala 59:15:@52086.4]
  assign FFRAM_io_banks_32_wdata_valid = io_banks_32_wdata_valid; // @[FIFO.scala 59:15:@52090.4]
  assign FFRAM_io_banks_32_wdata_bits = io_banks_32_wdata_bits; // @[FIFO.scala 59:15:@52089.4]
  assign FFRAM_io_banks_33_wdata_valid = io_banks_33_wdata_valid; // @[FIFO.scala 59:15:@52093.4]
  assign FFRAM_io_banks_33_wdata_bits = io_banks_33_wdata_bits; // @[FIFO.scala 59:15:@52092.4]
  assign FFRAM_io_banks_34_wdata_valid = io_banks_34_wdata_valid; // @[FIFO.scala 59:15:@52096.4]
  assign FFRAM_io_banks_34_wdata_bits = io_banks_34_wdata_bits; // @[FIFO.scala 59:15:@52095.4]
  assign FFRAM_io_banks_35_wdata_valid = io_banks_35_wdata_valid; // @[FIFO.scala 59:15:@52099.4]
  assign FFRAM_io_banks_35_wdata_bits = io_banks_35_wdata_bits; // @[FIFO.scala 59:15:@52098.4]
  assign FFRAM_io_banks_36_wdata_valid = io_banks_36_wdata_valid; // @[FIFO.scala 59:15:@52102.4]
  assign FFRAM_io_banks_36_wdata_bits = io_banks_36_wdata_bits; // @[FIFO.scala 59:15:@52101.4]
  assign FFRAM_io_banks_37_wdata_valid = io_banks_37_wdata_valid; // @[FIFO.scala 59:15:@52105.4]
  assign FFRAM_io_banks_37_wdata_bits = io_banks_37_wdata_bits; // @[FIFO.scala 59:15:@52104.4]
  assign FFRAM_io_banks_38_wdata_valid = io_banks_38_wdata_valid; // @[FIFO.scala 59:15:@52108.4]
  assign FFRAM_io_banks_38_wdata_bits = io_banks_38_wdata_bits; // @[FIFO.scala 59:15:@52107.4]
  assign FFRAM_io_banks_39_wdata_valid = io_banks_39_wdata_valid; // @[FIFO.scala 59:15:@52111.4]
  assign FFRAM_io_banks_39_wdata_bits = io_banks_39_wdata_bits; // @[FIFO.scala 59:15:@52110.4]
  assign FFRAM_io_banks_40_wdata_valid = io_banks_40_wdata_valid; // @[FIFO.scala 59:15:@52114.4]
  assign FFRAM_io_banks_40_wdata_bits = io_banks_40_wdata_bits; // @[FIFO.scala 59:15:@52113.4]
  assign FFRAM_io_banks_41_wdata_valid = io_banks_41_wdata_valid; // @[FIFO.scala 59:15:@52117.4]
  assign FFRAM_io_banks_41_wdata_bits = io_banks_41_wdata_bits; // @[FIFO.scala 59:15:@52116.4]
  assign FFRAM_io_banks_42_wdata_valid = io_banks_42_wdata_valid; // @[FIFO.scala 59:15:@52120.4]
  assign FFRAM_io_banks_42_wdata_bits = io_banks_42_wdata_bits; // @[FIFO.scala 59:15:@52119.4]
  assign FFRAM_io_banks_43_wdata_valid = io_banks_43_wdata_valid; // @[FIFO.scala 59:15:@52123.4]
  assign FFRAM_io_banks_43_wdata_bits = io_banks_43_wdata_bits; // @[FIFO.scala 59:15:@52122.4]
  assign FFRAM_io_banks_44_wdata_valid = io_banks_44_wdata_valid; // @[FIFO.scala 59:15:@52126.4]
  assign FFRAM_io_banks_44_wdata_bits = io_banks_44_wdata_bits; // @[FIFO.scala 59:15:@52125.4]
  assign FFRAM_io_banks_45_wdata_valid = io_banks_45_wdata_valid; // @[FIFO.scala 59:15:@52129.4]
  assign FFRAM_io_banks_45_wdata_bits = io_banks_45_wdata_bits; // @[FIFO.scala 59:15:@52128.4]
  assign FFRAM_io_banks_46_wdata_valid = io_banks_46_wdata_valid; // @[FIFO.scala 59:15:@52132.4]
  assign FFRAM_io_banks_46_wdata_bits = io_banks_46_wdata_bits; // @[FIFO.scala 59:15:@52131.4]
  assign FFRAM_io_banks_47_wdata_valid = io_banks_47_wdata_valid; // @[FIFO.scala 59:15:@52135.4]
  assign FFRAM_io_banks_47_wdata_bits = io_banks_47_wdata_bits; // @[FIFO.scala 59:15:@52134.4]
  assign FFRAM_io_banks_48_wdata_valid = io_banks_48_wdata_valid; // @[FIFO.scala 59:15:@52138.4]
  assign FFRAM_io_banks_48_wdata_bits = io_banks_48_wdata_bits; // @[FIFO.scala 59:15:@52137.4]
  assign FFRAM_io_banks_49_wdata_valid = io_banks_49_wdata_valid; // @[FIFO.scala 59:15:@52141.4]
  assign FFRAM_io_banks_49_wdata_bits = io_banks_49_wdata_bits; // @[FIFO.scala 59:15:@52140.4]
  assign FFRAM_io_banks_50_wdata_valid = io_banks_50_wdata_valid; // @[FIFO.scala 59:15:@52144.4]
  assign FFRAM_io_banks_50_wdata_bits = io_banks_50_wdata_bits; // @[FIFO.scala 59:15:@52143.4]
  assign FFRAM_io_banks_51_wdata_valid = io_banks_51_wdata_valid; // @[FIFO.scala 59:15:@52147.4]
  assign FFRAM_io_banks_51_wdata_bits = io_banks_51_wdata_bits; // @[FIFO.scala 59:15:@52146.4]
  assign FFRAM_io_banks_52_wdata_valid = io_banks_52_wdata_valid; // @[FIFO.scala 59:15:@52150.4]
  assign FFRAM_io_banks_52_wdata_bits = io_banks_52_wdata_bits; // @[FIFO.scala 59:15:@52149.4]
  assign FFRAM_io_banks_53_wdata_valid = io_banks_53_wdata_valid; // @[FIFO.scala 59:15:@52153.4]
  assign FFRAM_io_banks_53_wdata_bits = io_banks_53_wdata_bits; // @[FIFO.scala 59:15:@52152.4]
  assign FFRAM_io_banks_54_wdata_valid = io_banks_54_wdata_valid; // @[FIFO.scala 59:15:@52156.4]
  assign FFRAM_io_banks_54_wdata_bits = io_banks_54_wdata_bits; // @[FIFO.scala 59:15:@52155.4]
  assign FFRAM_io_banks_55_wdata_valid = io_banks_55_wdata_valid; // @[FIFO.scala 59:15:@52159.4]
  assign FFRAM_io_banks_55_wdata_bits = io_banks_55_wdata_bits; // @[FIFO.scala 59:15:@52158.4]
  assign FFRAM_io_banks_56_wdata_valid = io_banks_56_wdata_valid; // @[FIFO.scala 59:15:@52162.4]
  assign FFRAM_io_banks_56_wdata_bits = io_banks_56_wdata_bits; // @[FIFO.scala 59:15:@52161.4]
  assign FFRAM_io_banks_57_wdata_valid = io_banks_57_wdata_valid; // @[FIFO.scala 59:15:@52165.4]
  assign FFRAM_io_banks_57_wdata_bits = io_banks_57_wdata_bits; // @[FIFO.scala 59:15:@52164.4]
  assign FFRAM_io_banks_58_wdata_valid = io_banks_58_wdata_valid; // @[FIFO.scala 59:15:@52168.4]
  assign FFRAM_io_banks_58_wdata_bits = io_banks_58_wdata_bits; // @[FIFO.scala 59:15:@52167.4]
  assign FFRAM_io_banks_59_wdata_valid = io_banks_59_wdata_valid; // @[FIFO.scala 59:15:@52171.4]
  assign FFRAM_io_banks_59_wdata_bits = io_banks_59_wdata_bits; // @[FIFO.scala 59:15:@52170.4]
  assign FFRAM_io_banks_60_wdata_valid = io_banks_60_wdata_valid; // @[FIFO.scala 59:15:@52174.4]
  assign FFRAM_io_banks_60_wdata_bits = io_banks_60_wdata_bits; // @[FIFO.scala 59:15:@52173.4]
  assign FFRAM_io_banks_61_wdata_valid = io_banks_61_wdata_valid; // @[FIFO.scala 59:15:@52177.4]
  assign FFRAM_io_banks_61_wdata_bits = io_banks_61_wdata_bits; // @[FIFO.scala 59:15:@52176.4]
  assign FFRAM_io_banks_62_wdata_valid = io_banks_62_wdata_valid; // @[FIFO.scala 59:15:@52180.4]
  assign FFRAM_io_banks_62_wdata_bits = io_banks_62_wdata_bits; // @[FIFO.scala 59:15:@52179.4]
  assign FFRAM_io_banks_63_wdata_valid = io_banks_63_wdata_valid; // @[FIFO.scala 59:15:@52183.4]
  assign FFRAM_io_banks_63_wdata_bits = io_banks_63_wdata_bits; // @[FIFO.scala 59:15:@52182.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_1657) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module StreamControllerStore( // @[:@52962.2]
  input         clock, // @[:@52963.4]
  input         reset, // @[:@52964.4]
  input         io_dram_cmd_ready, // @[:@52965.4]
  output        io_dram_cmd_valid, // @[:@52965.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@52965.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@52965.4]
  input         io_dram_wdata_ready, // @[:@52965.4]
  output        io_dram_wdata_valid, // @[:@52965.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@52965.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@52965.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@52965.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@52965.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@52965.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@52965.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@52965.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@52965.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@52965.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@52965.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@52965.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@52965.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@52965.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@52965.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@52965.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@52965.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@52965.4]
  output        io_dram_wresp_ready, // @[:@52965.4]
  input         io_dram_wresp_valid, // @[:@52965.4]
  output        io_store_cmd_ready, // @[:@52965.4]
  input         io_store_cmd_valid, // @[:@52965.4]
  input  [63:0] io_store_cmd_bits_addr, // @[:@52965.4]
  input  [31:0] io_store_cmd_bits_size, // @[:@52965.4]
  output        io_store_data_ready, // @[:@52965.4]
  input         io_store_data_valid, // @[:@52965.4]
  input  [31:0] io_store_data_bits_wdata_0, // @[:@52965.4]
  input         io_store_data_bits_wstrb, // @[:@52965.4]
  input         io_store_wresp_ready, // @[:@52965.4]
  output        io_store_wresp_valid, // @[:@52965.4]
  output        io_store_wresp_bits // @[:@52965.4]
);
  wire  cmd_clock; // @[StreamController.scala 75:19:@53090.4]
  wire  cmd_reset; // @[StreamController.scala 75:19:@53090.4]
  wire  cmd_io_in_ready; // @[StreamController.scala 75:19:@53090.4]
  wire  cmd_io_in_valid; // @[StreamController.scala 75:19:@53090.4]
  wire [63:0] cmd_io_in_bits_addr; // @[StreamController.scala 75:19:@53090.4]
  wire [31:0] cmd_io_in_bits_size; // @[StreamController.scala 75:19:@53090.4]
  wire  cmd_io_out_ready; // @[StreamController.scala 75:19:@53090.4]
  wire  cmd_io_out_valid; // @[StreamController.scala 75:19:@53090.4]
  wire [63:0] cmd_io_out_bits_addr; // @[StreamController.scala 75:19:@53090.4]
  wire [31:0] cmd_io_out_bits_size; // @[StreamController.scala 75:19:@53090.4]
  wire  wdata_clock; // @[StreamController.scala 88:21:@53496.4]
  wire  wdata_reset; // @[StreamController.scala 88:21:@53496.4]
  wire  wdata_io_in_ready; // @[StreamController.scala 88:21:@53496.4]
  wire  wdata_io_in_valid; // @[StreamController.scala 88:21:@53496.4]
  wire [31:0] wdata_io_in_bits_data_0; // @[StreamController.scala 88:21:@53496.4]
  wire  wdata_io_in_bits_strobe; // @[StreamController.scala 88:21:@53496.4]
  wire  wdata_io_out_ready; // @[StreamController.scala 88:21:@53496.4]
  wire  wdata_io_out_valid; // @[StreamController.scala 88:21:@53496.4]
  wire [31:0] wdata_io_out_bits_data_0; // @[StreamController.scala 88:21:@53496.4]
  wire [31:0] wdata_io_out_bits_data_1; // @[StreamController.scala 88:21:@53496.4]
  wire [31:0] wdata_io_out_bits_data_2; // @[StreamController.scala 88:21:@53496.4]
  wire [31:0] wdata_io_out_bits_data_3; // @[StreamController.scala 88:21:@53496.4]
  wire [31:0] wdata_io_out_bits_data_4; // @[StreamController.scala 88:21:@53496.4]
  wire [31:0] wdata_io_out_bits_data_5; // @[StreamController.scala 88:21:@53496.4]
  wire [31:0] wdata_io_out_bits_data_6; // @[StreamController.scala 88:21:@53496.4]
  wire [31:0] wdata_io_out_bits_data_7; // @[StreamController.scala 88:21:@53496.4]
  wire [31:0] wdata_io_out_bits_data_8; // @[StreamController.scala 88:21:@53496.4]
  wire [31:0] wdata_io_out_bits_data_9; // @[StreamController.scala 88:21:@53496.4]
  wire [31:0] wdata_io_out_bits_data_10; // @[StreamController.scala 88:21:@53496.4]
  wire [31:0] wdata_io_out_bits_data_11; // @[StreamController.scala 88:21:@53496.4]
  wire [31:0] wdata_io_out_bits_data_12; // @[StreamController.scala 88:21:@53496.4]
  wire [31:0] wdata_io_out_bits_data_13; // @[StreamController.scala 88:21:@53496.4]
  wire [31:0] wdata_io_out_bits_data_14; // @[StreamController.scala 88:21:@53496.4]
  wire [31:0] wdata_io_out_bits_data_15; // @[StreamController.scala 88:21:@53496.4]
  wire [63:0] wdata_io_out_bits_strobe; // @[StreamController.scala 88:21:@53496.4]
  wire  wresp_clock; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_reset; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_in_ready; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_in_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_in_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_out_ready; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_out_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_out_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_0_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_0_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_1_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_1_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_2_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_2_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_3_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_3_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_4_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_4_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_5_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_5_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_6_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_6_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_7_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_7_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_8_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_8_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_9_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_9_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_10_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_10_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_11_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_11_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_12_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_12_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_13_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_13_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_14_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_14_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_15_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_15_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_16_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_16_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_17_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_17_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_18_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_18_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_19_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_19_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_20_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_20_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_21_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_21_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_22_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_22_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_23_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_23_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_24_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_24_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_25_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_25_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_26_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_26_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_27_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_27_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_28_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_28_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_29_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_29_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_30_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_30_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_31_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_31_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_32_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_32_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_33_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_33_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_34_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_34_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_35_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_35_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_36_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_36_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_37_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_37_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_38_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_38_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_39_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_39_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_40_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_40_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_41_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_41_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_42_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_42_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_43_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_43_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_44_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_44_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_45_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_45_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_46_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_46_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_47_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_47_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_48_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_48_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_49_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_49_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_50_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_50_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_51_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_51_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_52_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_52_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_53_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_53_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_54_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_54_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_55_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_55_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_56_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_56_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_57_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_57_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_58_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_58_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_59_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_59_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_60_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_60_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_61_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_61_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_62_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_62_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_63_wdata_valid; // @[StreamController.scala 100:21:@53737.4]
  wire  wresp_io_banks_63_wdata_bits; // @[StreamController.scala 100:21:@53737.4]
  wire [25:0] _T_111; // @[StreamController.scala 21:10:@53493.4]
  FIFO cmd ( // @[StreamController.scala 75:19:@53090.4]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_in_ready(cmd_io_in_ready),
    .io_in_valid(cmd_io_in_valid),
    .io_in_bits_addr(cmd_io_in_bits_addr),
    .io_in_bits_size(cmd_io_in_bits_size),
    .io_out_ready(cmd_io_out_ready),
    .io_out_valid(cmd_io_out_valid),
    .io_out_bits_addr(cmd_io_out_bits_addr),
    .io_out_bits_size(cmd_io_out_bits_size)
  );
  FIFOWidthConvert wdata ( // @[StreamController.scala 88:21:@53496.4]
    .clock(wdata_clock),
    .reset(wdata_reset),
    .io_in_ready(wdata_io_in_ready),
    .io_in_valid(wdata_io_in_valid),
    .io_in_bits_data_0(wdata_io_in_bits_data_0),
    .io_in_bits_strobe(wdata_io_in_bits_strobe),
    .io_out_ready(wdata_io_out_ready),
    .io_out_valid(wdata_io_out_valid),
    .io_out_bits_data_0(wdata_io_out_bits_data_0),
    .io_out_bits_data_1(wdata_io_out_bits_data_1),
    .io_out_bits_data_2(wdata_io_out_bits_data_2),
    .io_out_bits_data_3(wdata_io_out_bits_data_3),
    .io_out_bits_data_4(wdata_io_out_bits_data_4),
    .io_out_bits_data_5(wdata_io_out_bits_data_5),
    .io_out_bits_data_6(wdata_io_out_bits_data_6),
    .io_out_bits_data_7(wdata_io_out_bits_data_7),
    .io_out_bits_data_8(wdata_io_out_bits_data_8),
    .io_out_bits_data_9(wdata_io_out_bits_data_9),
    .io_out_bits_data_10(wdata_io_out_bits_data_10),
    .io_out_bits_data_11(wdata_io_out_bits_data_11),
    .io_out_bits_data_12(wdata_io_out_bits_data_12),
    .io_out_bits_data_13(wdata_io_out_bits_data_13),
    .io_out_bits_data_14(wdata_io_out_bits_data_14),
    .io_out_bits_data_15(wdata_io_out_bits_data_15),
    .io_out_bits_strobe(wdata_io_out_bits_strobe)
  );
  FIFO_33 wresp ( // @[StreamController.scala 100:21:@53737.4]
    .clock(wresp_clock),
    .reset(wresp_reset),
    .io_in_ready(wresp_io_in_ready),
    .io_in_valid(wresp_io_in_valid),
    .io_in_bits(wresp_io_in_bits),
    .io_out_ready(wresp_io_out_ready),
    .io_out_valid(wresp_io_out_valid),
    .io_out_bits(wresp_io_out_bits),
    .io_banks_0_wdata_valid(wresp_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(wresp_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(wresp_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(wresp_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(wresp_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(wresp_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(wresp_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(wresp_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(wresp_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(wresp_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(wresp_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(wresp_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(wresp_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(wresp_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(wresp_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(wresp_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(wresp_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(wresp_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(wresp_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(wresp_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(wresp_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(wresp_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(wresp_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(wresp_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(wresp_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(wresp_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(wresp_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(wresp_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(wresp_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(wresp_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(wresp_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(wresp_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(wresp_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(wresp_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(wresp_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(wresp_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(wresp_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(wresp_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(wresp_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(wresp_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(wresp_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(wresp_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(wresp_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(wresp_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(wresp_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(wresp_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(wresp_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(wresp_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(wresp_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(wresp_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(wresp_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(wresp_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(wresp_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(wresp_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(wresp_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(wresp_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(wresp_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(wresp_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(wresp_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(wresp_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(wresp_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(wresp_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(wresp_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(wresp_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(wresp_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(wresp_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(wresp_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(wresp_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(wresp_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(wresp_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(wresp_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(wresp_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(wresp_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(wresp_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(wresp_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(wresp_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(wresp_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(wresp_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(wresp_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(wresp_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(wresp_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(wresp_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(wresp_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(wresp_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(wresp_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(wresp_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(wresp_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(wresp_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(wresp_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(wresp_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(wresp_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(wresp_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(wresp_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(wresp_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(wresp_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(wresp_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(wresp_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(wresp_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(wresp_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(wresp_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(wresp_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(wresp_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(wresp_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(wresp_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(wresp_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(wresp_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(wresp_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(wresp_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(wresp_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(wresp_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(wresp_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(wresp_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(wresp_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(wresp_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(wresp_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(wresp_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(wresp_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(wresp_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(wresp_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(wresp_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(wresp_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(wresp_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(wresp_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(wresp_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(wresp_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(wresp_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(wresp_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(wresp_io_banks_63_wdata_bits)
  );
  assign _T_111 = cmd_io_out_bits_size[31:6]; // @[StreamController.scala 21:10:@53493.4]
  assign io_dram_cmd_valid = cmd_io_out_valid; // @[StreamController.scala 81:21:@53490.4]
  assign io_dram_cmd_bits_addr = cmd_io_out_bits_addr; // @[StreamController.scala 83:25:@53491.4]
  assign io_dram_cmd_bits_size = {{6'd0}, _T_111}; // @[StreamController.scala 85:25:@53494.4]
  assign io_dram_wdata_valid = wdata_io_out_valid; // @[StreamController.scala 95:23:@53526.4]
  assign io_dram_wdata_bits_wdata_0 = wdata_io_out_bits_data_0; // @[StreamController.scala 96:28:@53527.4]
  assign io_dram_wdata_bits_wdata_1 = wdata_io_out_bits_data_1; // @[StreamController.scala 96:28:@53528.4]
  assign io_dram_wdata_bits_wdata_2 = wdata_io_out_bits_data_2; // @[StreamController.scala 96:28:@53529.4]
  assign io_dram_wdata_bits_wdata_3 = wdata_io_out_bits_data_3; // @[StreamController.scala 96:28:@53530.4]
  assign io_dram_wdata_bits_wdata_4 = wdata_io_out_bits_data_4; // @[StreamController.scala 96:28:@53531.4]
  assign io_dram_wdata_bits_wdata_5 = wdata_io_out_bits_data_5; // @[StreamController.scala 96:28:@53532.4]
  assign io_dram_wdata_bits_wdata_6 = wdata_io_out_bits_data_6; // @[StreamController.scala 96:28:@53533.4]
  assign io_dram_wdata_bits_wdata_7 = wdata_io_out_bits_data_7; // @[StreamController.scala 96:28:@53534.4]
  assign io_dram_wdata_bits_wdata_8 = wdata_io_out_bits_data_8; // @[StreamController.scala 96:28:@53535.4]
  assign io_dram_wdata_bits_wdata_9 = wdata_io_out_bits_data_9; // @[StreamController.scala 96:28:@53536.4]
  assign io_dram_wdata_bits_wdata_10 = wdata_io_out_bits_data_10; // @[StreamController.scala 96:28:@53537.4]
  assign io_dram_wdata_bits_wdata_11 = wdata_io_out_bits_data_11; // @[StreamController.scala 96:28:@53538.4]
  assign io_dram_wdata_bits_wdata_12 = wdata_io_out_bits_data_12; // @[StreamController.scala 96:28:@53539.4]
  assign io_dram_wdata_bits_wdata_13 = wdata_io_out_bits_data_13; // @[StreamController.scala 96:28:@53540.4]
  assign io_dram_wdata_bits_wdata_14 = wdata_io_out_bits_data_14; // @[StreamController.scala 96:28:@53541.4]
  assign io_dram_wdata_bits_wdata_15 = wdata_io_out_bits_data_15; // @[StreamController.scala 96:28:@53542.4]
  assign io_dram_wdata_bits_wstrb_0 = wdata_io_out_bits_strobe[63]; // @[StreamController.scala 97:28:@53672.4]
  assign io_dram_wdata_bits_wstrb_1 = wdata_io_out_bits_strobe[62]; // @[StreamController.scala 97:28:@53673.4]
  assign io_dram_wdata_bits_wstrb_2 = wdata_io_out_bits_strobe[61]; // @[StreamController.scala 97:28:@53674.4]
  assign io_dram_wdata_bits_wstrb_3 = wdata_io_out_bits_strobe[60]; // @[StreamController.scala 97:28:@53675.4]
  assign io_dram_wdata_bits_wstrb_4 = wdata_io_out_bits_strobe[59]; // @[StreamController.scala 97:28:@53676.4]
  assign io_dram_wdata_bits_wstrb_5 = wdata_io_out_bits_strobe[58]; // @[StreamController.scala 97:28:@53677.4]
  assign io_dram_wdata_bits_wstrb_6 = wdata_io_out_bits_strobe[57]; // @[StreamController.scala 97:28:@53678.4]
  assign io_dram_wdata_bits_wstrb_7 = wdata_io_out_bits_strobe[56]; // @[StreamController.scala 97:28:@53679.4]
  assign io_dram_wdata_bits_wstrb_8 = wdata_io_out_bits_strobe[55]; // @[StreamController.scala 97:28:@53680.4]
  assign io_dram_wdata_bits_wstrb_9 = wdata_io_out_bits_strobe[54]; // @[StreamController.scala 97:28:@53681.4]
  assign io_dram_wdata_bits_wstrb_10 = wdata_io_out_bits_strobe[53]; // @[StreamController.scala 97:28:@53682.4]
  assign io_dram_wdata_bits_wstrb_11 = wdata_io_out_bits_strobe[52]; // @[StreamController.scala 97:28:@53683.4]
  assign io_dram_wdata_bits_wstrb_12 = wdata_io_out_bits_strobe[51]; // @[StreamController.scala 97:28:@53684.4]
  assign io_dram_wdata_bits_wstrb_13 = wdata_io_out_bits_strobe[50]; // @[StreamController.scala 97:28:@53685.4]
  assign io_dram_wdata_bits_wstrb_14 = wdata_io_out_bits_strobe[49]; // @[StreamController.scala 97:28:@53686.4]
  assign io_dram_wdata_bits_wstrb_15 = wdata_io_out_bits_strobe[48]; // @[StreamController.scala 97:28:@53687.4]
  assign io_dram_wdata_bits_wstrb_16 = wdata_io_out_bits_strobe[47]; // @[StreamController.scala 97:28:@53688.4]
  assign io_dram_wdata_bits_wstrb_17 = wdata_io_out_bits_strobe[46]; // @[StreamController.scala 97:28:@53689.4]
  assign io_dram_wdata_bits_wstrb_18 = wdata_io_out_bits_strobe[45]; // @[StreamController.scala 97:28:@53690.4]
  assign io_dram_wdata_bits_wstrb_19 = wdata_io_out_bits_strobe[44]; // @[StreamController.scala 97:28:@53691.4]
  assign io_dram_wdata_bits_wstrb_20 = wdata_io_out_bits_strobe[43]; // @[StreamController.scala 97:28:@53692.4]
  assign io_dram_wdata_bits_wstrb_21 = wdata_io_out_bits_strobe[42]; // @[StreamController.scala 97:28:@53693.4]
  assign io_dram_wdata_bits_wstrb_22 = wdata_io_out_bits_strobe[41]; // @[StreamController.scala 97:28:@53694.4]
  assign io_dram_wdata_bits_wstrb_23 = wdata_io_out_bits_strobe[40]; // @[StreamController.scala 97:28:@53695.4]
  assign io_dram_wdata_bits_wstrb_24 = wdata_io_out_bits_strobe[39]; // @[StreamController.scala 97:28:@53696.4]
  assign io_dram_wdata_bits_wstrb_25 = wdata_io_out_bits_strobe[38]; // @[StreamController.scala 97:28:@53697.4]
  assign io_dram_wdata_bits_wstrb_26 = wdata_io_out_bits_strobe[37]; // @[StreamController.scala 97:28:@53698.4]
  assign io_dram_wdata_bits_wstrb_27 = wdata_io_out_bits_strobe[36]; // @[StreamController.scala 97:28:@53699.4]
  assign io_dram_wdata_bits_wstrb_28 = wdata_io_out_bits_strobe[35]; // @[StreamController.scala 97:28:@53700.4]
  assign io_dram_wdata_bits_wstrb_29 = wdata_io_out_bits_strobe[34]; // @[StreamController.scala 97:28:@53701.4]
  assign io_dram_wdata_bits_wstrb_30 = wdata_io_out_bits_strobe[33]; // @[StreamController.scala 97:28:@53702.4]
  assign io_dram_wdata_bits_wstrb_31 = wdata_io_out_bits_strobe[32]; // @[StreamController.scala 97:28:@53703.4]
  assign io_dram_wdata_bits_wstrb_32 = wdata_io_out_bits_strobe[31]; // @[StreamController.scala 97:28:@53704.4]
  assign io_dram_wdata_bits_wstrb_33 = wdata_io_out_bits_strobe[30]; // @[StreamController.scala 97:28:@53705.4]
  assign io_dram_wdata_bits_wstrb_34 = wdata_io_out_bits_strobe[29]; // @[StreamController.scala 97:28:@53706.4]
  assign io_dram_wdata_bits_wstrb_35 = wdata_io_out_bits_strobe[28]; // @[StreamController.scala 97:28:@53707.4]
  assign io_dram_wdata_bits_wstrb_36 = wdata_io_out_bits_strobe[27]; // @[StreamController.scala 97:28:@53708.4]
  assign io_dram_wdata_bits_wstrb_37 = wdata_io_out_bits_strobe[26]; // @[StreamController.scala 97:28:@53709.4]
  assign io_dram_wdata_bits_wstrb_38 = wdata_io_out_bits_strobe[25]; // @[StreamController.scala 97:28:@53710.4]
  assign io_dram_wdata_bits_wstrb_39 = wdata_io_out_bits_strobe[24]; // @[StreamController.scala 97:28:@53711.4]
  assign io_dram_wdata_bits_wstrb_40 = wdata_io_out_bits_strobe[23]; // @[StreamController.scala 97:28:@53712.4]
  assign io_dram_wdata_bits_wstrb_41 = wdata_io_out_bits_strobe[22]; // @[StreamController.scala 97:28:@53713.4]
  assign io_dram_wdata_bits_wstrb_42 = wdata_io_out_bits_strobe[21]; // @[StreamController.scala 97:28:@53714.4]
  assign io_dram_wdata_bits_wstrb_43 = wdata_io_out_bits_strobe[20]; // @[StreamController.scala 97:28:@53715.4]
  assign io_dram_wdata_bits_wstrb_44 = wdata_io_out_bits_strobe[19]; // @[StreamController.scala 97:28:@53716.4]
  assign io_dram_wdata_bits_wstrb_45 = wdata_io_out_bits_strobe[18]; // @[StreamController.scala 97:28:@53717.4]
  assign io_dram_wdata_bits_wstrb_46 = wdata_io_out_bits_strobe[17]; // @[StreamController.scala 97:28:@53718.4]
  assign io_dram_wdata_bits_wstrb_47 = wdata_io_out_bits_strobe[16]; // @[StreamController.scala 97:28:@53719.4]
  assign io_dram_wdata_bits_wstrb_48 = wdata_io_out_bits_strobe[15]; // @[StreamController.scala 97:28:@53720.4]
  assign io_dram_wdata_bits_wstrb_49 = wdata_io_out_bits_strobe[14]; // @[StreamController.scala 97:28:@53721.4]
  assign io_dram_wdata_bits_wstrb_50 = wdata_io_out_bits_strobe[13]; // @[StreamController.scala 97:28:@53722.4]
  assign io_dram_wdata_bits_wstrb_51 = wdata_io_out_bits_strobe[12]; // @[StreamController.scala 97:28:@53723.4]
  assign io_dram_wdata_bits_wstrb_52 = wdata_io_out_bits_strobe[11]; // @[StreamController.scala 97:28:@53724.4]
  assign io_dram_wdata_bits_wstrb_53 = wdata_io_out_bits_strobe[10]; // @[StreamController.scala 97:28:@53725.4]
  assign io_dram_wdata_bits_wstrb_54 = wdata_io_out_bits_strobe[9]; // @[StreamController.scala 97:28:@53726.4]
  assign io_dram_wdata_bits_wstrb_55 = wdata_io_out_bits_strobe[8]; // @[StreamController.scala 97:28:@53727.4]
  assign io_dram_wdata_bits_wstrb_56 = wdata_io_out_bits_strobe[7]; // @[StreamController.scala 97:28:@53728.4]
  assign io_dram_wdata_bits_wstrb_57 = wdata_io_out_bits_strobe[6]; // @[StreamController.scala 97:28:@53729.4]
  assign io_dram_wdata_bits_wstrb_58 = wdata_io_out_bits_strobe[5]; // @[StreamController.scala 97:28:@53730.4]
  assign io_dram_wdata_bits_wstrb_59 = wdata_io_out_bits_strobe[4]; // @[StreamController.scala 97:28:@53731.4]
  assign io_dram_wdata_bits_wstrb_60 = wdata_io_out_bits_strobe[3]; // @[StreamController.scala 97:28:@53732.4]
  assign io_dram_wdata_bits_wstrb_61 = wdata_io_out_bits_strobe[2]; // @[StreamController.scala 97:28:@53733.4]
  assign io_dram_wdata_bits_wstrb_62 = wdata_io_out_bits_strobe[1]; // @[StreamController.scala 97:28:@53734.4]
  assign io_dram_wdata_bits_wstrb_63 = wdata_io_out_bits_strobe[0]; // @[StreamController.scala 97:28:@53735.4]
  assign io_dram_wresp_ready = wresp_io_in_ready; // @[StreamController.scala 104:23:@54004.4]
  assign io_store_cmd_ready = cmd_io_in_ready; // @[StreamController.scala 79:22:@53488.4]
  assign io_store_data_ready = wdata_io_in_ready; // @[StreamController.scala 93:23:@53525.4]
  assign io_store_wresp_valid = wresp_io_out_valid; // @[StreamController.scala 106:24:@54005.4]
  assign io_store_wresp_bits = wresp_io_out_bits; // @[StreamController.scala 107:23:@54006.4]
  assign cmd_clock = clock; // @[:@53091.4]
  assign cmd_reset = reset; // @[:@53092.4]
  assign cmd_io_in_valid = io_store_cmd_valid; // @[StreamController.scala 77:19:@53485.4]
  assign cmd_io_in_bits_addr = io_store_cmd_bits_addr; // @[StreamController.scala 78:18:@53487.4]
  assign cmd_io_in_bits_size = io_store_cmd_bits_size; // @[StreamController.scala 78:18:@53486.4]
  assign cmd_io_out_ready = io_dram_cmd_ready; // @[StreamController.scala 80:20:@53489.4]
  assign wdata_clock = clock; // @[:@53497.4]
  assign wdata_reset = reset; // @[:@53498.4]
  assign wdata_io_in_valid = io_store_data_valid; // @[StreamController.scala 90:21:@53522.4]
  assign wdata_io_in_bits_data_0 = io_store_data_bits_wdata_0; // @[StreamController.scala 91:25:@53523.4]
  assign wdata_io_in_bits_strobe = io_store_data_bits_wstrb; // @[StreamController.scala 92:27:@53524.4]
  assign wdata_io_out_ready = io_dram_wdata_ready; // @[StreamController.scala 98:22:@53736.4]
  assign wresp_clock = clock; // @[:@53738.4]
  assign wresp_reset = reset; // @[:@53739.4]
  assign wresp_io_in_valid = io_dram_wresp_valid; // @[StreamController.scala 102:21:@54002.4]
  assign wresp_io_in_bits = 1'h1; // @[StreamController.scala 103:20:@54003.4]
  assign wresp_io_out_ready = io_store_wresp_ready; // @[StreamController.scala 108:22:@54007.4]
  assign wresp_io_banks_0_wdata_valid = 1'h0;
  assign wresp_io_banks_0_wdata_bits = 1'h0;
  assign wresp_io_banks_1_wdata_valid = 1'h0;
  assign wresp_io_banks_1_wdata_bits = 1'h0;
  assign wresp_io_banks_2_wdata_valid = 1'h0;
  assign wresp_io_banks_2_wdata_bits = 1'h0;
  assign wresp_io_banks_3_wdata_valid = 1'h0;
  assign wresp_io_banks_3_wdata_bits = 1'h0;
  assign wresp_io_banks_4_wdata_valid = 1'h0;
  assign wresp_io_banks_4_wdata_bits = 1'h0;
  assign wresp_io_banks_5_wdata_valid = 1'h0;
  assign wresp_io_banks_5_wdata_bits = 1'h0;
  assign wresp_io_banks_6_wdata_valid = 1'h0;
  assign wresp_io_banks_6_wdata_bits = 1'h0;
  assign wresp_io_banks_7_wdata_valid = 1'h0;
  assign wresp_io_banks_7_wdata_bits = 1'h0;
  assign wresp_io_banks_8_wdata_valid = 1'h0;
  assign wresp_io_banks_8_wdata_bits = 1'h0;
  assign wresp_io_banks_9_wdata_valid = 1'h0;
  assign wresp_io_banks_9_wdata_bits = 1'h0;
  assign wresp_io_banks_10_wdata_valid = 1'h0;
  assign wresp_io_banks_10_wdata_bits = 1'h0;
  assign wresp_io_banks_11_wdata_valid = 1'h0;
  assign wresp_io_banks_11_wdata_bits = 1'h0;
  assign wresp_io_banks_12_wdata_valid = 1'h0;
  assign wresp_io_banks_12_wdata_bits = 1'h0;
  assign wresp_io_banks_13_wdata_valid = 1'h0;
  assign wresp_io_banks_13_wdata_bits = 1'h0;
  assign wresp_io_banks_14_wdata_valid = 1'h0;
  assign wresp_io_banks_14_wdata_bits = 1'h0;
  assign wresp_io_banks_15_wdata_valid = 1'h0;
  assign wresp_io_banks_15_wdata_bits = 1'h0;
  assign wresp_io_banks_16_wdata_valid = 1'h0;
  assign wresp_io_banks_16_wdata_bits = 1'h0;
  assign wresp_io_banks_17_wdata_valid = 1'h0;
  assign wresp_io_banks_17_wdata_bits = 1'h0;
  assign wresp_io_banks_18_wdata_valid = 1'h0;
  assign wresp_io_banks_18_wdata_bits = 1'h0;
  assign wresp_io_banks_19_wdata_valid = 1'h0;
  assign wresp_io_banks_19_wdata_bits = 1'h0;
  assign wresp_io_banks_20_wdata_valid = 1'h0;
  assign wresp_io_banks_20_wdata_bits = 1'h0;
  assign wresp_io_banks_21_wdata_valid = 1'h0;
  assign wresp_io_banks_21_wdata_bits = 1'h0;
  assign wresp_io_banks_22_wdata_valid = 1'h0;
  assign wresp_io_banks_22_wdata_bits = 1'h0;
  assign wresp_io_banks_23_wdata_valid = 1'h0;
  assign wresp_io_banks_23_wdata_bits = 1'h0;
  assign wresp_io_banks_24_wdata_valid = 1'h0;
  assign wresp_io_banks_24_wdata_bits = 1'h0;
  assign wresp_io_banks_25_wdata_valid = 1'h0;
  assign wresp_io_banks_25_wdata_bits = 1'h0;
  assign wresp_io_banks_26_wdata_valid = 1'h0;
  assign wresp_io_banks_26_wdata_bits = 1'h0;
  assign wresp_io_banks_27_wdata_valid = 1'h0;
  assign wresp_io_banks_27_wdata_bits = 1'h0;
  assign wresp_io_banks_28_wdata_valid = 1'h0;
  assign wresp_io_banks_28_wdata_bits = 1'h0;
  assign wresp_io_banks_29_wdata_valid = 1'h0;
  assign wresp_io_banks_29_wdata_bits = 1'h0;
  assign wresp_io_banks_30_wdata_valid = 1'h0;
  assign wresp_io_banks_30_wdata_bits = 1'h0;
  assign wresp_io_banks_31_wdata_valid = 1'h0;
  assign wresp_io_banks_31_wdata_bits = 1'h0;
  assign wresp_io_banks_32_wdata_valid = 1'h0;
  assign wresp_io_banks_32_wdata_bits = 1'h0;
  assign wresp_io_banks_33_wdata_valid = 1'h0;
  assign wresp_io_banks_33_wdata_bits = 1'h0;
  assign wresp_io_banks_34_wdata_valid = 1'h0;
  assign wresp_io_banks_34_wdata_bits = 1'h0;
  assign wresp_io_banks_35_wdata_valid = 1'h0;
  assign wresp_io_banks_35_wdata_bits = 1'h0;
  assign wresp_io_banks_36_wdata_valid = 1'h0;
  assign wresp_io_banks_36_wdata_bits = 1'h0;
  assign wresp_io_banks_37_wdata_valid = 1'h0;
  assign wresp_io_banks_37_wdata_bits = 1'h0;
  assign wresp_io_banks_38_wdata_valid = 1'h0;
  assign wresp_io_banks_38_wdata_bits = 1'h0;
  assign wresp_io_banks_39_wdata_valid = 1'h0;
  assign wresp_io_banks_39_wdata_bits = 1'h0;
  assign wresp_io_banks_40_wdata_valid = 1'h0;
  assign wresp_io_banks_40_wdata_bits = 1'h0;
  assign wresp_io_banks_41_wdata_valid = 1'h0;
  assign wresp_io_banks_41_wdata_bits = 1'h0;
  assign wresp_io_banks_42_wdata_valid = 1'h0;
  assign wresp_io_banks_42_wdata_bits = 1'h0;
  assign wresp_io_banks_43_wdata_valid = 1'h0;
  assign wresp_io_banks_43_wdata_bits = 1'h0;
  assign wresp_io_banks_44_wdata_valid = 1'h0;
  assign wresp_io_banks_44_wdata_bits = 1'h0;
  assign wresp_io_banks_45_wdata_valid = 1'h0;
  assign wresp_io_banks_45_wdata_bits = 1'h0;
  assign wresp_io_banks_46_wdata_valid = 1'h0;
  assign wresp_io_banks_46_wdata_bits = 1'h0;
  assign wresp_io_banks_47_wdata_valid = 1'h0;
  assign wresp_io_banks_47_wdata_bits = 1'h0;
  assign wresp_io_banks_48_wdata_valid = 1'h0;
  assign wresp_io_banks_48_wdata_bits = 1'h0;
  assign wresp_io_banks_49_wdata_valid = 1'h0;
  assign wresp_io_banks_49_wdata_bits = 1'h0;
  assign wresp_io_banks_50_wdata_valid = 1'h0;
  assign wresp_io_banks_50_wdata_bits = 1'h0;
  assign wresp_io_banks_51_wdata_valid = 1'h0;
  assign wresp_io_banks_51_wdata_bits = 1'h0;
  assign wresp_io_banks_52_wdata_valid = 1'h0;
  assign wresp_io_banks_52_wdata_bits = 1'h0;
  assign wresp_io_banks_53_wdata_valid = 1'h0;
  assign wresp_io_banks_53_wdata_bits = 1'h0;
  assign wresp_io_banks_54_wdata_valid = 1'h0;
  assign wresp_io_banks_54_wdata_bits = 1'h0;
  assign wresp_io_banks_55_wdata_valid = 1'h0;
  assign wresp_io_banks_55_wdata_bits = 1'h0;
  assign wresp_io_banks_56_wdata_valid = 1'h0;
  assign wresp_io_banks_56_wdata_bits = 1'h0;
  assign wresp_io_banks_57_wdata_valid = 1'h0;
  assign wresp_io_banks_57_wdata_bits = 1'h0;
  assign wresp_io_banks_58_wdata_valid = 1'h0;
  assign wresp_io_banks_58_wdata_bits = 1'h0;
  assign wresp_io_banks_59_wdata_valid = 1'h0;
  assign wresp_io_banks_59_wdata_bits = 1'h0;
  assign wresp_io_banks_60_wdata_valid = 1'h0;
  assign wresp_io_banks_60_wdata_bits = 1'h0;
  assign wresp_io_banks_61_wdata_valid = 1'h0;
  assign wresp_io_banks_61_wdata_bits = 1'h0;
  assign wresp_io_banks_62_wdata_valid = 1'h0;
  assign wresp_io_banks_62_wdata_bits = 1'h0;
  assign wresp_io_banks_63_wdata_valid = 1'h0;
  assign wresp_io_banks_63_wdata_bits = 1'h0;
endmodule
module MuxPipe( // @[:@54073.2]
  output        io_in_ready, // @[:@54076.4]
  input         io_in_valid, // @[:@54076.4]
  input  [63:0] io_in_bits_0_addr, // @[:@54076.4]
  input  [31:0] io_in_bits_0_size, // @[:@54076.4]
  input         io_in_bits_0_isWr, // @[:@54076.4]
  input  [31:0] io_in_bits_0_tag, // @[:@54076.4]
  input         io_out_ready, // @[:@54076.4]
  output        io_out_valid, // @[:@54076.4]
  output [63:0] io_out_bits_addr, // @[:@54076.4]
  output [31:0] io_out_bits_size, // @[:@54076.4]
  output        io_out_bits_isWr, // @[:@54076.4]
  output [31:0] io_out_bits_tag // @[:@54076.4]
);
  wire  _T_42; // @[MuxN.scala 28:31:@54078.4]
  assign _T_42 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@54078.4]
  assign io_in_ready = io_out_ready | _T_42; // @[MuxN.scala 71:15:@54087.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@54086.4]
  assign io_out_bits_addr = io_in_bits_0_addr; // @[MuxN.scala 72:15:@54092.4]
  assign io_out_bits_size = io_in_bits_0_size; // @[MuxN.scala 72:15:@54091.4]
  assign io_out_bits_isWr = io_in_bits_0_isWr; // @[MuxN.scala 72:15:@54089.4]
  assign io_out_bits_tag = io_in_bits_0_tag; // @[MuxN.scala 72:15:@54088.4]
endmodule
module MuxPipe_1( // @[:@54094.2]
  output        io_in_ready, // @[:@54097.4]
  input         io_in_valid, // @[:@54097.4]
  input  [31:0] io_in_bits_0_wdata_0, // @[:@54097.4]
  input  [31:0] io_in_bits_0_wdata_1, // @[:@54097.4]
  input  [31:0] io_in_bits_0_wdata_2, // @[:@54097.4]
  input  [31:0] io_in_bits_0_wdata_3, // @[:@54097.4]
  input  [31:0] io_in_bits_0_wdata_4, // @[:@54097.4]
  input  [31:0] io_in_bits_0_wdata_5, // @[:@54097.4]
  input  [31:0] io_in_bits_0_wdata_6, // @[:@54097.4]
  input  [31:0] io_in_bits_0_wdata_7, // @[:@54097.4]
  input  [31:0] io_in_bits_0_wdata_8, // @[:@54097.4]
  input  [31:0] io_in_bits_0_wdata_9, // @[:@54097.4]
  input  [31:0] io_in_bits_0_wdata_10, // @[:@54097.4]
  input  [31:0] io_in_bits_0_wdata_11, // @[:@54097.4]
  input  [31:0] io_in_bits_0_wdata_12, // @[:@54097.4]
  input  [31:0] io_in_bits_0_wdata_13, // @[:@54097.4]
  input  [31:0] io_in_bits_0_wdata_14, // @[:@54097.4]
  input  [31:0] io_in_bits_0_wdata_15, // @[:@54097.4]
  input         io_in_bits_0_wstrb_0, // @[:@54097.4]
  input         io_in_bits_0_wstrb_1, // @[:@54097.4]
  input         io_in_bits_0_wstrb_2, // @[:@54097.4]
  input         io_in_bits_0_wstrb_3, // @[:@54097.4]
  input         io_in_bits_0_wstrb_4, // @[:@54097.4]
  input         io_in_bits_0_wstrb_5, // @[:@54097.4]
  input         io_in_bits_0_wstrb_6, // @[:@54097.4]
  input         io_in_bits_0_wstrb_7, // @[:@54097.4]
  input         io_in_bits_0_wstrb_8, // @[:@54097.4]
  input         io_in_bits_0_wstrb_9, // @[:@54097.4]
  input         io_in_bits_0_wstrb_10, // @[:@54097.4]
  input         io_in_bits_0_wstrb_11, // @[:@54097.4]
  input         io_in_bits_0_wstrb_12, // @[:@54097.4]
  input         io_in_bits_0_wstrb_13, // @[:@54097.4]
  input         io_in_bits_0_wstrb_14, // @[:@54097.4]
  input         io_in_bits_0_wstrb_15, // @[:@54097.4]
  input         io_in_bits_0_wstrb_16, // @[:@54097.4]
  input         io_in_bits_0_wstrb_17, // @[:@54097.4]
  input         io_in_bits_0_wstrb_18, // @[:@54097.4]
  input         io_in_bits_0_wstrb_19, // @[:@54097.4]
  input         io_in_bits_0_wstrb_20, // @[:@54097.4]
  input         io_in_bits_0_wstrb_21, // @[:@54097.4]
  input         io_in_bits_0_wstrb_22, // @[:@54097.4]
  input         io_in_bits_0_wstrb_23, // @[:@54097.4]
  input         io_in_bits_0_wstrb_24, // @[:@54097.4]
  input         io_in_bits_0_wstrb_25, // @[:@54097.4]
  input         io_in_bits_0_wstrb_26, // @[:@54097.4]
  input         io_in_bits_0_wstrb_27, // @[:@54097.4]
  input         io_in_bits_0_wstrb_28, // @[:@54097.4]
  input         io_in_bits_0_wstrb_29, // @[:@54097.4]
  input         io_in_bits_0_wstrb_30, // @[:@54097.4]
  input         io_in_bits_0_wstrb_31, // @[:@54097.4]
  input         io_in_bits_0_wstrb_32, // @[:@54097.4]
  input         io_in_bits_0_wstrb_33, // @[:@54097.4]
  input         io_in_bits_0_wstrb_34, // @[:@54097.4]
  input         io_in_bits_0_wstrb_35, // @[:@54097.4]
  input         io_in_bits_0_wstrb_36, // @[:@54097.4]
  input         io_in_bits_0_wstrb_37, // @[:@54097.4]
  input         io_in_bits_0_wstrb_38, // @[:@54097.4]
  input         io_in_bits_0_wstrb_39, // @[:@54097.4]
  input         io_in_bits_0_wstrb_40, // @[:@54097.4]
  input         io_in_bits_0_wstrb_41, // @[:@54097.4]
  input         io_in_bits_0_wstrb_42, // @[:@54097.4]
  input         io_in_bits_0_wstrb_43, // @[:@54097.4]
  input         io_in_bits_0_wstrb_44, // @[:@54097.4]
  input         io_in_bits_0_wstrb_45, // @[:@54097.4]
  input         io_in_bits_0_wstrb_46, // @[:@54097.4]
  input         io_in_bits_0_wstrb_47, // @[:@54097.4]
  input         io_in_bits_0_wstrb_48, // @[:@54097.4]
  input         io_in_bits_0_wstrb_49, // @[:@54097.4]
  input         io_in_bits_0_wstrb_50, // @[:@54097.4]
  input         io_in_bits_0_wstrb_51, // @[:@54097.4]
  input         io_in_bits_0_wstrb_52, // @[:@54097.4]
  input         io_in_bits_0_wstrb_53, // @[:@54097.4]
  input         io_in_bits_0_wstrb_54, // @[:@54097.4]
  input         io_in_bits_0_wstrb_55, // @[:@54097.4]
  input         io_in_bits_0_wstrb_56, // @[:@54097.4]
  input         io_in_bits_0_wstrb_57, // @[:@54097.4]
  input         io_in_bits_0_wstrb_58, // @[:@54097.4]
  input         io_in_bits_0_wstrb_59, // @[:@54097.4]
  input         io_in_bits_0_wstrb_60, // @[:@54097.4]
  input         io_in_bits_0_wstrb_61, // @[:@54097.4]
  input         io_in_bits_0_wstrb_62, // @[:@54097.4]
  input         io_in_bits_0_wstrb_63, // @[:@54097.4]
  input         io_out_ready, // @[:@54097.4]
  output        io_out_valid, // @[:@54097.4]
  output [31:0] io_out_bits_wdata_0, // @[:@54097.4]
  output [31:0] io_out_bits_wdata_1, // @[:@54097.4]
  output [31:0] io_out_bits_wdata_2, // @[:@54097.4]
  output [31:0] io_out_bits_wdata_3, // @[:@54097.4]
  output [31:0] io_out_bits_wdata_4, // @[:@54097.4]
  output [31:0] io_out_bits_wdata_5, // @[:@54097.4]
  output [31:0] io_out_bits_wdata_6, // @[:@54097.4]
  output [31:0] io_out_bits_wdata_7, // @[:@54097.4]
  output [31:0] io_out_bits_wdata_8, // @[:@54097.4]
  output [31:0] io_out_bits_wdata_9, // @[:@54097.4]
  output [31:0] io_out_bits_wdata_10, // @[:@54097.4]
  output [31:0] io_out_bits_wdata_11, // @[:@54097.4]
  output [31:0] io_out_bits_wdata_12, // @[:@54097.4]
  output [31:0] io_out_bits_wdata_13, // @[:@54097.4]
  output [31:0] io_out_bits_wdata_14, // @[:@54097.4]
  output [31:0] io_out_bits_wdata_15, // @[:@54097.4]
  output        io_out_bits_wstrb_0, // @[:@54097.4]
  output        io_out_bits_wstrb_1, // @[:@54097.4]
  output        io_out_bits_wstrb_2, // @[:@54097.4]
  output        io_out_bits_wstrb_3, // @[:@54097.4]
  output        io_out_bits_wstrb_4, // @[:@54097.4]
  output        io_out_bits_wstrb_5, // @[:@54097.4]
  output        io_out_bits_wstrb_6, // @[:@54097.4]
  output        io_out_bits_wstrb_7, // @[:@54097.4]
  output        io_out_bits_wstrb_8, // @[:@54097.4]
  output        io_out_bits_wstrb_9, // @[:@54097.4]
  output        io_out_bits_wstrb_10, // @[:@54097.4]
  output        io_out_bits_wstrb_11, // @[:@54097.4]
  output        io_out_bits_wstrb_12, // @[:@54097.4]
  output        io_out_bits_wstrb_13, // @[:@54097.4]
  output        io_out_bits_wstrb_14, // @[:@54097.4]
  output        io_out_bits_wstrb_15, // @[:@54097.4]
  output        io_out_bits_wstrb_16, // @[:@54097.4]
  output        io_out_bits_wstrb_17, // @[:@54097.4]
  output        io_out_bits_wstrb_18, // @[:@54097.4]
  output        io_out_bits_wstrb_19, // @[:@54097.4]
  output        io_out_bits_wstrb_20, // @[:@54097.4]
  output        io_out_bits_wstrb_21, // @[:@54097.4]
  output        io_out_bits_wstrb_22, // @[:@54097.4]
  output        io_out_bits_wstrb_23, // @[:@54097.4]
  output        io_out_bits_wstrb_24, // @[:@54097.4]
  output        io_out_bits_wstrb_25, // @[:@54097.4]
  output        io_out_bits_wstrb_26, // @[:@54097.4]
  output        io_out_bits_wstrb_27, // @[:@54097.4]
  output        io_out_bits_wstrb_28, // @[:@54097.4]
  output        io_out_bits_wstrb_29, // @[:@54097.4]
  output        io_out_bits_wstrb_30, // @[:@54097.4]
  output        io_out_bits_wstrb_31, // @[:@54097.4]
  output        io_out_bits_wstrb_32, // @[:@54097.4]
  output        io_out_bits_wstrb_33, // @[:@54097.4]
  output        io_out_bits_wstrb_34, // @[:@54097.4]
  output        io_out_bits_wstrb_35, // @[:@54097.4]
  output        io_out_bits_wstrb_36, // @[:@54097.4]
  output        io_out_bits_wstrb_37, // @[:@54097.4]
  output        io_out_bits_wstrb_38, // @[:@54097.4]
  output        io_out_bits_wstrb_39, // @[:@54097.4]
  output        io_out_bits_wstrb_40, // @[:@54097.4]
  output        io_out_bits_wstrb_41, // @[:@54097.4]
  output        io_out_bits_wstrb_42, // @[:@54097.4]
  output        io_out_bits_wstrb_43, // @[:@54097.4]
  output        io_out_bits_wstrb_44, // @[:@54097.4]
  output        io_out_bits_wstrb_45, // @[:@54097.4]
  output        io_out_bits_wstrb_46, // @[:@54097.4]
  output        io_out_bits_wstrb_47, // @[:@54097.4]
  output        io_out_bits_wstrb_48, // @[:@54097.4]
  output        io_out_bits_wstrb_49, // @[:@54097.4]
  output        io_out_bits_wstrb_50, // @[:@54097.4]
  output        io_out_bits_wstrb_51, // @[:@54097.4]
  output        io_out_bits_wstrb_52, // @[:@54097.4]
  output        io_out_bits_wstrb_53, // @[:@54097.4]
  output        io_out_bits_wstrb_54, // @[:@54097.4]
  output        io_out_bits_wstrb_55, // @[:@54097.4]
  output        io_out_bits_wstrb_56, // @[:@54097.4]
  output        io_out_bits_wstrb_57, // @[:@54097.4]
  output        io_out_bits_wstrb_58, // @[:@54097.4]
  output        io_out_bits_wstrb_59, // @[:@54097.4]
  output        io_out_bits_wstrb_60, // @[:@54097.4]
  output        io_out_bits_wstrb_61, // @[:@54097.4]
  output        io_out_bits_wstrb_62, // @[:@54097.4]
  output        io_out_bits_wstrb_63 // @[:@54097.4]
);
  wire  _T_146; // @[MuxN.scala 28:31:@54099.4]
  assign _T_146 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@54099.4]
  assign io_in_ready = io_out_ready | _T_146; // @[MuxN.scala 71:15:@54184.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@54183.4]
  assign io_out_bits_wdata_0 = io_in_bits_0_wdata_0; // @[MuxN.scala 72:15:@54250.4]
  assign io_out_bits_wdata_1 = io_in_bits_0_wdata_1; // @[MuxN.scala 72:15:@54251.4]
  assign io_out_bits_wdata_2 = io_in_bits_0_wdata_2; // @[MuxN.scala 72:15:@54252.4]
  assign io_out_bits_wdata_3 = io_in_bits_0_wdata_3; // @[MuxN.scala 72:15:@54253.4]
  assign io_out_bits_wdata_4 = io_in_bits_0_wdata_4; // @[MuxN.scala 72:15:@54254.4]
  assign io_out_bits_wdata_5 = io_in_bits_0_wdata_5; // @[MuxN.scala 72:15:@54255.4]
  assign io_out_bits_wdata_6 = io_in_bits_0_wdata_6; // @[MuxN.scala 72:15:@54256.4]
  assign io_out_bits_wdata_7 = io_in_bits_0_wdata_7; // @[MuxN.scala 72:15:@54257.4]
  assign io_out_bits_wdata_8 = io_in_bits_0_wdata_8; // @[MuxN.scala 72:15:@54258.4]
  assign io_out_bits_wdata_9 = io_in_bits_0_wdata_9; // @[MuxN.scala 72:15:@54259.4]
  assign io_out_bits_wdata_10 = io_in_bits_0_wdata_10; // @[MuxN.scala 72:15:@54260.4]
  assign io_out_bits_wdata_11 = io_in_bits_0_wdata_11; // @[MuxN.scala 72:15:@54261.4]
  assign io_out_bits_wdata_12 = io_in_bits_0_wdata_12; // @[MuxN.scala 72:15:@54262.4]
  assign io_out_bits_wdata_13 = io_in_bits_0_wdata_13; // @[MuxN.scala 72:15:@54263.4]
  assign io_out_bits_wdata_14 = io_in_bits_0_wdata_14; // @[MuxN.scala 72:15:@54264.4]
  assign io_out_bits_wdata_15 = io_in_bits_0_wdata_15; // @[MuxN.scala 72:15:@54265.4]
  assign io_out_bits_wstrb_0 = io_in_bits_0_wstrb_0; // @[MuxN.scala 72:15:@54186.4]
  assign io_out_bits_wstrb_1 = io_in_bits_0_wstrb_1; // @[MuxN.scala 72:15:@54187.4]
  assign io_out_bits_wstrb_2 = io_in_bits_0_wstrb_2; // @[MuxN.scala 72:15:@54188.4]
  assign io_out_bits_wstrb_3 = io_in_bits_0_wstrb_3; // @[MuxN.scala 72:15:@54189.4]
  assign io_out_bits_wstrb_4 = io_in_bits_0_wstrb_4; // @[MuxN.scala 72:15:@54190.4]
  assign io_out_bits_wstrb_5 = io_in_bits_0_wstrb_5; // @[MuxN.scala 72:15:@54191.4]
  assign io_out_bits_wstrb_6 = io_in_bits_0_wstrb_6; // @[MuxN.scala 72:15:@54192.4]
  assign io_out_bits_wstrb_7 = io_in_bits_0_wstrb_7; // @[MuxN.scala 72:15:@54193.4]
  assign io_out_bits_wstrb_8 = io_in_bits_0_wstrb_8; // @[MuxN.scala 72:15:@54194.4]
  assign io_out_bits_wstrb_9 = io_in_bits_0_wstrb_9; // @[MuxN.scala 72:15:@54195.4]
  assign io_out_bits_wstrb_10 = io_in_bits_0_wstrb_10; // @[MuxN.scala 72:15:@54196.4]
  assign io_out_bits_wstrb_11 = io_in_bits_0_wstrb_11; // @[MuxN.scala 72:15:@54197.4]
  assign io_out_bits_wstrb_12 = io_in_bits_0_wstrb_12; // @[MuxN.scala 72:15:@54198.4]
  assign io_out_bits_wstrb_13 = io_in_bits_0_wstrb_13; // @[MuxN.scala 72:15:@54199.4]
  assign io_out_bits_wstrb_14 = io_in_bits_0_wstrb_14; // @[MuxN.scala 72:15:@54200.4]
  assign io_out_bits_wstrb_15 = io_in_bits_0_wstrb_15; // @[MuxN.scala 72:15:@54201.4]
  assign io_out_bits_wstrb_16 = io_in_bits_0_wstrb_16; // @[MuxN.scala 72:15:@54202.4]
  assign io_out_bits_wstrb_17 = io_in_bits_0_wstrb_17; // @[MuxN.scala 72:15:@54203.4]
  assign io_out_bits_wstrb_18 = io_in_bits_0_wstrb_18; // @[MuxN.scala 72:15:@54204.4]
  assign io_out_bits_wstrb_19 = io_in_bits_0_wstrb_19; // @[MuxN.scala 72:15:@54205.4]
  assign io_out_bits_wstrb_20 = io_in_bits_0_wstrb_20; // @[MuxN.scala 72:15:@54206.4]
  assign io_out_bits_wstrb_21 = io_in_bits_0_wstrb_21; // @[MuxN.scala 72:15:@54207.4]
  assign io_out_bits_wstrb_22 = io_in_bits_0_wstrb_22; // @[MuxN.scala 72:15:@54208.4]
  assign io_out_bits_wstrb_23 = io_in_bits_0_wstrb_23; // @[MuxN.scala 72:15:@54209.4]
  assign io_out_bits_wstrb_24 = io_in_bits_0_wstrb_24; // @[MuxN.scala 72:15:@54210.4]
  assign io_out_bits_wstrb_25 = io_in_bits_0_wstrb_25; // @[MuxN.scala 72:15:@54211.4]
  assign io_out_bits_wstrb_26 = io_in_bits_0_wstrb_26; // @[MuxN.scala 72:15:@54212.4]
  assign io_out_bits_wstrb_27 = io_in_bits_0_wstrb_27; // @[MuxN.scala 72:15:@54213.4]
  assign io_out_bits_wstrb_28 = io_in_bits_0_wstrb_28; // @[MuxN.scala 72:15:@54214.4]
  assign io_out_bits_wstrb_29 = io_in_bits_0_wstrb_29; // @[MuxN.scala 72:15:@54215.4]
  assign io_out_bits_wstrb_30 = io_in_bits_0_wstrb_30; // @[MuxN.scala 72:15:@54216.4]
  assign io_out_bits_wstrb_31 = io_in_bits_0_wstrb_31; // @[MuxN.scala 72:15:@54217.4]
  assign io_out_bits_wstrb_32 = io_in_bits_0_wstrb_32; // @[MuxN.scala 72:15:@54218.4]
  assign io_out_bits_wstrb_33 = io_in_bits_0_wstrb_33; // @[MuxN.scala 72:15:@54219.4]
  assign io_out_bits_wstrb_34 = io_in_bits_0_wstrb_34; // @[MuxN.scala 72:15:@54220.4]
  assign io_out_bits_wstrb_35 = io_in_bits_0_wstrb_35; // @[MuxN.scala 72:15:@54221.4]
  assign io_out_bits_wstrb_36 = io_in_bits_0_wstrb_36; // @[MuxN.scala 72:15:@54222.4]
  assign io_out_bits_wstrb_37 = io_in_bits_0_wstrb_37; // @[MuxN.scala 72:15:@54223.4]
  assign io_out_bits_wstrb_38 = io_in_bits_0_wstrb_38; // @[MuxN.scala 72:15:@54224.4]
  assign io_out_bits_wstrb_39 = io_in_bits_0_wstrb_39; // @[MuxN.scala 72:15:@54225.4]
  assign io_out_bits_wstrb_40 = io_in_bits_0_wstrb_40; // @[MuxN.scala 72:15:@54226.4]
  assign io_out_bits_wstrb_41 = io_in_bits_0_wstrb_41; // @[MuxN.scala 72:15:@54227.4]
  assign io_out_bits_wstrb_42 = io_in_bits_0_wstrb_42; // @[MuxN.scala 72:15:@54228.4]
  assign io_out_bits_wstrb_43 = io_in_bits_0_wstrb_43; // @[MuxN.scala 72:15:@54229.4]
  assign io_out_bits_wstrb_44 = io_in_bits_0_wstrb_44; // @[MuxN.scala 72:15:@54230.4]
  assign io_out_bits_wstrb_45 = io_in_bits_0_wstrb_45; // @[MuxN.scala 72:15:@54231.4]
  assign io_out_bits_wstrb_46 = io_in_bits_0_wstrb_46; // @[MuxN.scala 72:15:@54232.4]
  assign io_out_bits_wstrb_47 = io_in_bits_0_wstrb_47; // @[MuxN.scala 72:15:@54233.4]
  assign io_out_bits_wstrb_48 = io_in_bits_0_wstrb_48; // @[MuxN.scala 72:15:@54234.4]
  assign io_out_bits_wstrb_49 = io_in_bits_0_wstrb_49; // @[MuxN.scala 72:15:@54235.4]
  assign io_out_bits_wstrb_50 = io_in_bits_0_wstrb_50; // @[MuxN.scala 72:15:@54236.4]
  assign io_out_bits_wstrb_51 = io_in_bits_0_wstrb_51; // @[MuxN.scala 72:15:@54237.4]
  assign io_out_bits_wstrb_52 = io_in_bits_0_wstrb_52; // @[MuxN.scala 72:15:@54238.4]
  assign io_out_bits_wstrb_53 = io_in_bits_0_wstrb_53; // @[MuxN.scala 72:15:@54239.4]
  assign io_out_bits_wstrb_54 = io_in_bits_0_wstrb_54; // @[MuxN.scala 72:15:@54240.4]
  assign io_out_bits_wstrb_55 = io_in_bits_0_wstrb_55; // @[MuxN.scala 72:15:@54241.4]
  assign io_out_bits_wstrb_56 = io_in_bits_0_wstrb_56; // @[MuxN.scala 72:15:@54242.4]
  assign io_out_bits_wstrb_57 = io_in_bits_0_wstrb_57; // @[MuxN.scala 72:15:@54243.4]
  assign io_out_bits_wstrb_58 = io_in_bits_0_wstrb_58; // @[MuxN.scala 72:15:@54244.4]
  assign io_out_bits_wstrb_59 = io_in_bits_0_wstrb_59; // @[MuxN.scala 72:15:@54245.4]
  assign io_out_bits_wstrb_60 = io_in_bits_0_wstrb_60; // @[MuxN.scala 72:15:@54246.4]
  assign io_out_bits_wstrb_61 = io_in_bits_0_wstrb_61; // @[MuxN.scala 72:15:@54247.4]
  assign io_out_bits_wstrb_62 = io_in_bits_0_wstrb_62; // @[MuxN.scala 72:15:@54248.4]
  assign io_out_bits_wstrb_63 = io_in_bits_0_wstrb_63; // @[MuxN.scala 72:15:@54249.4]
endmodule
module ElementCounter( // @[:@54267.2]
  input         clock, // @[:@54268.4]
  input         reset, // @[:@54269.4]
  input         io_reset, // @[:@54270.4]
  input         io_enable, // @[:@54270.4]
  output [31:0] io_out // @[:@54270.4]
);
  reg [31:0] count; // @[Counter.scala 37:22:@54272.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_14; // @[Counter.scala 39:24:@54273.4]
  wire [31:0] newCount; // @[Counter.scala 39:24:@54274.4]
  wire [31:0] _GEN_0; // @[Counter.scala 43:26:@54279.6]
  wire [31:0] _GEN_1; // @[Counter.scala 41:18:@54275.4]
  assign _T_14 = count + 32'h1; // @[Counter.scala 39:24:@54273.4]
  assign newCount = count + 32'h1; // @[Counter.scala 39:24:@54274.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 43:26:@54279.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 41:18:@54275.4]
  assign io_out = count; // @[Counter.scala 47:10:@54282.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module StreamArbiter( // @[:@54284.2]
  input         clock, // @[:@54285.4]
  input         reset, // @[:@54286.4]
  output        io_app_0_cmd_ready, // @[:@54287.4]
  input         io_app_0_cmd_valid, // @[:@54287.4]
  input  [63:0] io_app_0_cmd_bits_addr, // @[:@54287.4]
  input  [31:0] io_app_0_cmd_bits_size, // @[:@54287.4]
  input         io_app_0_cmd_bits_isWr, // @[:@54287.4]
  input  [31:0] io_app_0_cmd_bits_tag, // @[:@54287.4]
  output        io_app_0_wdata_ready, // @[:@54287.4]
  input         io_app_0_wdata_valid, // @[:@54287.4]
  input  [31:0] io_app_0_wdata_bits_wdata_0, // @[:@54287.4]
  input  [31:0] io_app_0_wdata_bits_wdata_1, // @[:@54287.4]
  input  [31:0] io_app_0_wdata_bits_wdata_2, // @[:@54287.4]
  input  [31:0] io_app_0_wdata_bits_wdata_3, // @[:@54287.4]
  input  [31:0] io_app_0_wdata_bits_wdata_4, // @[:@54287.4]
  input  [31:0] io_app_0_wdata_bits_wdata_5, // @[:@54287.4]
  input  [31:0] io_app_0_wdata_bits_wdata_6, // @[:@54287.4]
  input  [31:0] io_app_0_wdata_bits_wdata_7, // @[:@54287.4]
  input  [31:0] io_app_0_wdata_bits_wdata_8, // @[:@54287.4]
  input  [31:0] io_app_0_wdata_bits_wdata_9, // @[:@54287.4]
  input  [31:0] io_app_0_wdata_bits_wdata_10, // @[:@54287.4]
  input  [31:0] io_app_0_wdata_bits_wdata_11, // @[:@54287.4]
  input  [31:0] io_app_0_wdata_bits_wdata_12, // @[:@54287.4]
  input  [31:0] io_app_0_wdata_bits_wdata_13, // @[:@54287.4]
  input  [31:0] io_app_0_wdata_bits_wdata_14, // @[:@54287.4]
  input  [31:0] io_app_0_wdata_bits_wdata_15, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_0, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_1, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_2, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_3, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_4, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_5, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_6, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_7, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_8, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_9, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_10, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_11, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_12, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_13, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_14, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_15, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_16, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_17, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_18, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_19, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_20, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_21, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_22, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_23, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_24, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_25, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_26, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_27, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_28, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_29, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_30, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_31, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_32, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_33, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_34, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_35, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_36, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_37, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_38, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_39, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_40, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_41, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_42, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_43, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_44, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_45, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_46, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_47, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_48, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_49, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_50, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_51, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_52, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_53, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_54, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_55, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_56, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_57, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_58, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_59, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_60, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_61, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_62, // @[:@54287.4]
  input         io_app_0_wdata_bits_wstrb_63, // @[:@54287.4]
  input         io_app_0_rresp_ready, // @[:@54287.4]
  input         io_app_0_wresp_ready, // @[:@54287.4]
  output        io_app_0_wresp_valid, // @[:@54287.4]
  input         io_dram_cmd_ready, // @[:@54287.4]
  output        io_dram_cmd_valid, // @[:@54287.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@54287.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@54287.4]
  output        io_dram_cmd_bits_isWr, // @[:@54287.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@54287.4]
  input         io_dram_wdata_ready, // @[:@54287.4]
  output        io_dram_wdata_valid, // @[:@54287.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@54287.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@54287.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@54287.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@54287.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@54287.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@54287.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@54287.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@54287.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@54287.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@54287.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@54287.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@54287.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@54287.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@54287.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@54287.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@54287.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@54287.4]
  output        io_dram_rresp_ready, // @[:@54287.4]
  output        io_dram_wresp_ready, // @[:@54287.4]
  input         io_dram_wresp_valid, // @[:@54287.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@54287.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@54516.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@54516.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@54516.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@54516.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@54516.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@54523.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@54523.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@54523.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@54523.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@54523.4]
  wire  cmdMux_io_in_ready; // @[StreamArbiter.scala 25:22:@54533.4]
  wire  cmdMux_io_in_valid; // @[StreamArbiter.scala 25:22:@54533.4]
  wire [63:0] cmdMux_io_in_bits_0_addr; // @[StreamArbiter.scala 25:22:@54533.4]
  wire [31:0] cmdMux_io_in_bits_0_size; // @[StreamArbiter.scala 25:22:@54533.4]
  wire  cmdMux_io_in_bits_0_isWr; // @[StreamArbiter.scala 25:22:@54533.4]
  wire [31:0] cmdMux_io_in_bits_0_tag; // @[StreamArbiter.scala 25:22:@54533.4]
  wire  cmdMux_io_out_ready; // @[StreamArbiter.scala 25:22:@54533.4]
  wire  cmdMux_io_out_valid; // @[StreamArbiter.scala 25:22:@54533.4]
  wire [63:0] cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 25:22:@54533.4]
  wire [31:0] cmdMux_io_out_bits_size; // @[StreamArbiter.scala 25:22:@54533.4]
  wire  cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 25:22:@54533.4]
  wire [31:0] cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 25:22:@54533.4]
  wire  wdataMux_io_in_ready; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_valid; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_0; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_1; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_2; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_3; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_4; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_5; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_6; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_7; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_8; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_9; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_10; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_11; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_12; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_13; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_14; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_15; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_0; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_1; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_2; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_3; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_4; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_5; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_6; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_7; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_8; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_9; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_10; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_11; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_12; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_13; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_14; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_15; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_16; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_17; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_18; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_19; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_20; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_21; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_22; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_23; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_24; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_25; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_26; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_27; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_28; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_29; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_30; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_31; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_32; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_33; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_34; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_35; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_36; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_37; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_38; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_39; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_40; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_41; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_42; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_43; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_44; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_45; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_46; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_47; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_48; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_49; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_50; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_51; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_52; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_53; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_54; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_55; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_56; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_57; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_58; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_59; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_60; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_61; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_62; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_in_bits_0_wstrb_63; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_ready; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_valid; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 35:24:@54556.4]
  wire [31:0] wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 35:24:@54556.4]
  wire  elementCtr_clock; // @[StreamArbiter.scala 36:26:@54559.4]
  wire  elementCtr_reset; // @[StreamArbiter.scala 36:26:@54559.4]
  wire  elementCtr_io_reset; // @[StreamArbiter.scala 36:26:@54559.4]
  wire  elementCtr_io_enable; // @[StreamArbiter.scala 36:26:@54559.4]
  wire [31:0] elementCtr_io_out; // @[StreamArbiter.scala 36:26:@54559.4]
  wire  _T_346; // @[package.scala 96:25:@54528.4 package.scala 96:25:@54529.4]
  wire  cmdIdx; // @[StreamArbiter.scala 21:16:@54530.4]
  wire [1:0] cmdInDecoder; // @[OneHot.scala 45:35:@54532.4]
  wire  _T_355; // @[FringeBundles.scala 114:28:@54548.4]
  wire [22:0] _T_356; // @[FringeBundles.scala 114:28:@54550.4]
  wire [23:0] _T_358; // @[FringeBundles.scala 115:37:@54553.4]
  wire  _T_360; // @[StreamArbiter.scala 37:49:@54562.4]
  wire [31:0] _T_365; // @[:@54566.4 :@54567.4]
  wire [7:0] _T_366; // @[FringeBundles.scala 114:28:@54568.4]
  wire [255:0] cmdOutDecoder; // @[OneHot.scala 45:35:@54574.4]
  wire  _T_379; // @[StreamArbiter.scala 42:78:@54577.4]
  wire  _T_380; // @[StreamArbiter.scala 42:121:@54578.4]
  wire [7:0] _T_395; // @[FringeBundles.scala 140:28:@54765.4]
  wire [255:0] wrespDecoder; // @[OneHot.scala 45:35:@54772.4]
  wire  _T_400; // @[StreamArbiter.scala 61:55:@54777.4]
  wire  _T_403; // @[StreamArbiter.scala 62:85:@54781.4]
  wire  _T_404; // @[StreamArbiter.scala 62:70:@54782.4]
  wire  _T_409; // @[StreamArbiter.scala 67:58:@54806.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@54516.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@54523.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  MuxPipe cmdMux ( // @[StreamArbiter.scala 25:22:@54533.4]
    .io_in_ready(cmdMux_io_in_ready),
    .io_in_valid(cmdMux_io_in_valid),
    .io_in_bits_0_addr(cmdMux_io_in_bits_0_addr),
    .io_in_bits_0_size(cmdMux_io_in_bits_0_size),
    .io_in_bits_0_isWr(cmdMux_io_in_bits_0_isWr),
    .io_in_bits_0_tag(cmdMux_io_in_bits_0_tag),
    .io_out_ready(cmdMux_io_out_ready),
    .io_out_valid(cmdMux_io_out_valid),
    .io_out_bits_addr(cmdMux_io_out_bits_addr),
    .io_out_bits_size(cmdMux_io_out_bits_size),
    .io_out_bits_isWr(cmdMux_io_out_bits_isWr),
    .io_out_bits_tag(cmdMux_io_out_bits_tag)
  );
  MuxPipe_1 wdataMux ( // @[StreamArbiter.scala 35:24:@54556.4]
    .io_in_ready(wdataMux_io_in_ready),
    .io_in_valid(wdataMux_io_in_valid),
    .io_in_bits_0_wdata_0(wdataMux_io_in_bits_0_wdata_0),
    .io_in_bits_0_wdata_1(wdataMux_io_in_bits_0_wdata_1),
    .io_in_bits_0_wdata_2(wdataMux_io_in_bits_0_wdata_2),
    .io_in_bits_0_wdata_3(wdataMux_io_in_bits_0_wdata_3),
    .io_in_bits_0_wdata_4(wdataMux_io_in_bits_0_wdata_4),
    .io_in_bits_0_wdata_5(wdataMux_io_in_bits_0_wdata_5),
    .io_in_bits_0_wdata_6(wdataMux_io_in_bits_0_wdata_6),
    .io_in_bits_0_wdata_7(wdataMux_io_in_bits_0_wdata_7),
    .io_in_bits_0_wdata_8(wdataMux_io_in_bits_0_wdata_8),
    .io_in_bits_0_wdata_9(wdataMux_io_in_bits_0_wdata_9),
    .io_in_bits_0_wdata_10(wdataMux_io_in_bits_0_wdata_10),
    .io_in_bits_0_wdata_11(wdataMux_io_in_bits_0_wdata_11),
    .io_in_bits_0_wdata_12(wdataMux_io_in_bits_0_wdata_12),
    .io_in_bits_0_wdata_13(wdataMux_io_in_bits_0_wdata_13),
    .io_in_bits_0_wdata_14(wdataMux_io_in_bits_0_wdata_14),
    .io_in_bits_0_wdata_15(wdataMux_io_in_bits_0_wdata_15),
    .io_in_bits_0_wstrb_0(wdataMux_io_in_bits_0_wstrb_0),
    .io_in_bits_0_wstrb_1(wdataMux_io_in_bits_0_wstrb_1),
    .io_in_bits_0_wstrb_2(wdataMux_io_in_bits_0_wstrb_2),
    .io_in_bits_0_wstrb_3(wdataMux_io_in_bits_0_wstrb_3),
    .io_in_bits_0_wstrb_4(wdataMux_io_in_bits_0_wstrb_4),
    .io_in_bits_0_wstrb_5(wdataMux_io_in_bits_0_wstrb_5),
    .io_in_bits_0_wstrb_6(wdataMux_io_in_bits_0_wstrb_6),
    .io_in_bits_0_wstrb_7(wdataMux_io_in_bits_0_wstrb_7),
    .io_in_bits_0_wstrb_8(wdataMux_io_in_bits_0_wstrb_8),
    .io_in_bits_0_wstrb_9(wdataMux_io_in_bits_0_wstrb_9),
    .io_in_bits_0_wstrb_10(wdataMux_io_in_bits_0_wstrb_10),
    .io_in_bits_0_wstrb_11(wdataMux_io_in_bits_0_wstrb_11),
    .io_in_bits_0_wstrb_12(wdataMux_io_in_bits_0_wstrb_12),
    .io_in_bits_0_wstrb_13(wdataMux_io_in_bits_0_wstrb_13),
    .io_in_bits_0_wstrb_14(wdataMux_io_in_bits_0_wstrb_14),
    .io_in_bits_0_wstrb_15(wdataMux_io_in_bits_0_wstrb_15),
    .io_in_bits_0_wstrb_16(wdataMux_io_in_bits_0_wstrb_16),
    .io_in_bits_0_wstrb_17(wdataMux_io_in_bits_0_wstrb_17),
    .io_in_bits_0_wstrb_18(wdataMux_io_in_bits_0_wstrb_18),
    .io_in_bits_0_wstrb_19(wdataMux_io_in_bits_0_wstrb_19),
    .io_in_bits_0_wstrb_20(wdataMux_io_in_bits_0_wstrb_20),
    .io_in_bits_0_wstrb_21(wdataMux_io_in_bits_0_wstrb_21),
    .io_in_bits_0_wstrb_22(wdataMux_io_in_bits_0_wstrb_22),
    .io_in_bits_0_wstrb_23(wdataMux_io_in_bits_0_wstrb_23),
    .io_in_bits_0_wstrb_24(wdataMux_io_in_bits_0_wstrb_24),
    .io_in_bits_0_wstrb_25(wdataMux_io_in_bits_0_wstrb_25),
    .io_in_bits_0_wstrb_26(wdataMux_io_in_bits_0_wstrb_26),
    .io_in_bits_0_wstrb_27(wdataMux_io_in_bits_0_wstrb_27),
    .io_in_bits_0_wstrb_28(wdataMux_io_in_bits_0_wstrb_28),
    .io_in_bits_0_wstrb_29(wdataMux_io_in_bits_0_wstrb_29),
    .io_in_bits_0_wstrb_30(wdataMux_io_in_bits_0_wstrb_30),
    .io_in_bits_0_wstrb_31(wdataMux_io_in_bits_0_wstrb_31),
    .io_in_bits_0_wstrb_32(wdataMux_io_in_bits_0_wstrb_32),
    .io_in_bits_0_wstrb_33(wdataMux_io_in_bits_0_wstrb_33),
    .io_in_bits_0_wstrb_34(wdataMux_io_in_bits_0_wstrb_34),
    .io_in_bits_0_wstrb_35(wdataMux_io_in_bits_0_wstrb_35),
    .io_in_bits_0_wstrb_36(wdataMux_io_in_bits_0_wstrb_36),
    .io_in_bits_0_wstrb_37(wdataMux_io_in_bits_0_wstrb_37),
    .io_in_bits_0_wstrb_38(wdataMux_io_in_bits_0_wstrb_38),
    .io_in_bits_0_wstrb_39(wdataMux_io_in_bits_0_wstrb_39),
    .io_in_bits_0_wstrb_40(wdataMux_io_in_bits_0_wstrb_40),
    .io_in_bits_0_wstrb_41(wdataMux_io_in_bits_0_wstrb_41),
    .io_in_bits_0_wstrb_42(wdataMux_io_in_bits_0_wstrb_42),
    .io_in_bits_0_wstrb_43(wdataMux_io_in_bits_0_wstrb_43),
    .io_in_bits_0_wstrb_44(wdataMux_io_in_bits_0_wstrb_44),
    .io_in_bits_0_wstrb_45(wdataMux_io_in_bits_0_wstrb_45),
    .io_in_bits_0_wstrb_46(wdataMux_io_in_bits_0_wstrb_46),
    .io_in_bits_0_wstrb_47(wdataMux_io_in_bits_0_wstrb_47),
    .io_in_bits_0_wstrb_48(wdataMux_io_in_bits_0_wstrb_48),
    .io_in_bits_0_wstrb_49(wdataMux_io_in_bits_0_wstrb_49),
    .io_in_bits_0_wstrb_50(wdataMux_io_in_bits_0_wstrb_50),
    .io_in_bits_0_wstrb_51(wdataMux_io_in_bits_0_wstrb_51),
    .io_in_bits_0_wstrb_52(wdataMux_io_in_bits_0_wstrb_52),
    .io_in_bits_0_wstrb_53(wdataMux_io_in_bits_0_wstrb_53),
    .io_in_bits_0_wstrb_54(wdataMux_io_in_bits_0_wstrb_54),
    .io_in_bits_0_wstrb_55(wdataMux_io_in_bits_0_wstrb_55),
    .io_in_bits_0_wstrb_56(wdataMux_io_in_bits_0_wstrb_56),
    .io_in_bits_0_wstrb_57(wdataMux_io_in_bits_0_wstrb_57),
    .io_in_bits_0_wstrb_58(wdataMux_io_in_bits_0_wstrb_58),
    .io_in_bits_0_wstrb_59(wdataMux_io_in_bits_0_wstrb_59),
    .io_in_bits_0_wstrb_60(wdataMux_io_in_bits_0_wstrb_60),
    .io_in_bits_0_wstrb_61(wdataMux_io_in_bits_0_wstrb_61),
    .io_in_bits_0_wstrb_62(wdataMux_io_in_bits_0_wstrb_62),
    .io_in_bits_0_wstrb_63(wdataMux_io_in_bits_0_wstrb_63),
    .io_out_ready(wdataMux_io_out_ready),
    .io_out_valid(wdataMux_io_out_valid),
    .io_out_bits_wdata_0(wdataMux_io_out_bits_wdata_0),
    .io_out_bits_wdata_1(wdataMux_io_out_bits_wdata_1),
    .io_out_bits_wdata_2(wdataMux_io_out_bits_wdata_2),
    .io_out_bits_wdata_3(wdataMux_io_out_bits_wdata_3),
    .io_out_bits_wdata_4(wdataMux_io_out_bits_wdata_4),
    .io_out_bits_wdata_5(wdataMux_io_out_bits_wdata_5),
    .io_out_bits_wdata_6(wdataMux_io_out_bits_wdata_6),
    .io_out_bits_wdata_7(wdataMux_io_out_bits_wdata_7),
    .io_out_bits_wdata_8(wdataMux_io_out_bits_wdata_8),
    .io_out_bits_wdata_9(wdataMux_io_out_bits_wdata_9),
    .io_out_bits_wdata_10(wdataMux_io_out_bits_wdata_10),
    .io_out_bits_wdata_11(wdataMux_io_out_bits_wdata_11),
    .io_out_bits_wdata_12(wdataMux_io_out_bits_wdata_12),
    .io_out_bits_wdata_13(wdataMux_io_out_bits_wdata_13),
    .io_out_bits_wdata_14(wdataMux_io_out_bits_wdata_14),
    .io_out_bits_wdata_15(wdataMux_io_out_bits_wdata_15),
    .io_out_bits_wstrb_0(wdataMux_io_out_bits_wstrb_0),
    .io_out_bits_wstrb_1(wdataMux_io_out_bits_wstrb_1),
    .io_out_bits_wstrb_2(wdataMux_io_out_bits_wstrb_2),
    .io_out_bits_wstrb_3(wdataMux_io_out_bits_wstrb_3),
    .io_out_bits_wstrb_4(wdataMux_io_out_bits_wstrb_4),
    .io_out_bits_wstrb_5(wdataMux_io_out_bits_wstrb_5),
    .io_out_bits_wstrb_6(wdataMux_io_out_bits_wstrb_6),
    .io_out_bits_wstrb_7(wdataMux_io_out_bits_wstrb_7),
    .io_out_bits_wstrb_8(wdataMux_io_out_bits_wstrb_8),
    .io_out_bits_wstrb_9(wdataMux_io_out_bits_wstrb_9),
    .io_out_bits_wstrb_10(wdataMux_io_out_bits_wstrb_10),
    .io_out_bits_wstrb_11(wdataMux_io_out_bits_wstrb_11),
    .io_out_bits_wstrb_12(wdataMux_io_out_bits_wstrb_12),
    .io_out_bits_wstrb_13(wdataMux_io_out_bits_wstrb_13),
    .io_out_bits_wstrb_14(wdataMux_io_out_bits_wstrb_14),
    .io_out_bits_wstrb_15(wdataMux_io_out_bits_wstrb_15),
    .io_out_bits_wstrb_16(wdataMux_io_out_bits_wstrb_16),
    .io_out_bits_wstrb_17(wdataMux_io_out_bits_wstrb_17),
    .io_out_bits_wstrb_18(wdataMux_io_out_bits_wstrb_18),
    .io_out_bits_wstrb_19(wdataMux_io_out_bits_wstrb_19),
    .io_out_bits_wstrb_20(wdataMux_io_out_bits_wstrb_20),
    .io_out_bits_wstrb_21(wdataMux_io_out_bits_wstrb_21),
    .io_out_bits_wstrb_22(wdataMux_io_out_bits_wstrb_22),
    .io_out_bits_wstrb_23(wdataMux_io_out_bits_wstrb_23),
    .io_out_bits_wstrb_24(wdataMux_io_out_bits_wstrb_24),
    .io_out_bits_wstrb_25(wdataMux_io_out_bits_wstrb_25),
    .io_out_bits_wstrb_26(wdataMux_io_out_bits_wstrb_26),
    .io_out_bits_wstrb_27(wdataMux_io_out_bits_wstrb_27),
    .io_out_bits_wstrb_28(wdataMux_io_out_bits_wstrb_28),
    .io_out_bits_wstrb_29(wdataMux_io_out_bits_wstrb_29),
    .io_out_bits_wstrb_30(wdataMux_io_out_bits_wstrb_30),
    .io_out_bits_wstrb_31(wdataMux_io_out_bits_wstrb_31),
    .io_out_bits_wstrb_32(wdataMux_io_out_bits_wstrb_32),
    .io_out_bits_wstrb_33(wdataMux_io_out_bits_wstrb_33),
    .io_out_bits_wstrb_34(wdataMux_io_out_bits_wstrb_34),
    .io_out_bits_wstrb_35(wdataMux_io_out_bits_wstrb_35),
    .io_out_bits_wstrb_36(wdataMux_io_out_bits_wstrb_36),
    .io_out_bits_wstrb_37(wdataMux_io_out_bits_wstrb_37),
    .io_out_bits_wstrb_38(wdataMux_io_out_bits_wstrb_38),
    .io_out_bits_wstrb_39(wdataMux_io_out_bits_wstrb_39),
    .io_out_bits_wstrb_40(wdataMux_io_out_bits_wstrb_40),
    .io_out_bits_wstrb_41(wdataMux_io_out_bits_wstrb_41),
    .io_out_bits_wstrb_42(wdataMux_io_out_bits_wstrb_42),
    .io_out_bits_wstrb_43(wdataMux_io_out_bits_wstrb_43),
    .io_out_bits_wstrb_44(wdataMux_io_out_bits_wstrb_44),
    .io_out_bits_wstrb_45(wdataMux_io_out_bits_wstrb_45),
    .io_out_bits_wstrb_46(wdataMux_io_out_bits_wstrb_46),
    .io_out_bits_wstrb_47(wdataMux_io_out_bits_wstrb_47),
    .io_out_bits_wstrb_48(wdataMux_io_out_bits_wstrb_48),
    .io_out_bits_wstrb_49(wdataMux_io_out_bits_wstrb_49),
    .io_out_bits_wstrb_50(wdataMux_io_out_bits_wstrb_50),
    .io_out_bits_wstrb_51(wdataMux_io_out_bits_wstrb_51),
    .io_out_bits_wstrb_52(wdataMux_io_out_bits_wstrb_52),
    .io_out_bits_wstrb_53(wdataMux_io_out_bits_wstrb_53),
    .io_out_bits_wstrb_54(wdataMux_io_out_bits_wstrb_54),
    .io_out_bits_wstrb_55(wdataMux_io_out_bits_wstrb_55),
    .io_out_bits_wstrb_56(wdataMux_io_out_bits_wstrb_56),
    .io_out_bits_wstrb_57(wdataMux_io_out_bits_wstrb_57),
    .io_out_bits_wstrb_58(wdataMux_io_out_bits_wstrb_58),
    .io_out_bits_wstrb_59(wdataMux_io_out_bits_wstrb_59),
    .io_out_bits_wstrb_60(wdataMux_io_out_bits_wstrb_60),
    .io_out_bits_wstrb_61(wdataMux_io_out_bits_wstrb_61),
    .io_out_bits_wstrb_62(wdataMux_io_out_bits_wstrb_62),
    .io_out_bits_wstrb_63(wdataMux_io_out_bits_wstrb_63)
  );
  ElementCounter elementCtr ( // @[StreamArbiter.scala 36:26:@54559.4]
    .clock(elementCtr_clock),
    .reset(elementCtr_reset),
    .io_reset(elementCtr_io_reset),
    .io_enable(elementCtr_io_enable),
    .io_out(elementCtr_io_out)
  );
  assign _T_346 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@54528.4 package.scala 96:25:@54529.4]
  assign cmdIdx = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[StreamArbiter.scala 21:16:@54530.4]
  assign cmdInDecoder = 2'h1 << cmdIdx; // @[OneHot.scala 45:35:@54532.4]
  assign _T_355 = io_app_0_cmd_bits_tag[8]; // @[FringeBundles.scala 114:28:@54548.4]
  assign _T_356 = io_app_0_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@54550.4]
  assign _T_358 = {_T_356,_T_355}; // @[FringeBundles.scala 115:37:@54553.4]
  assign _T_360 = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:49:@54562.4]
  assign _T_365 = cmdMux_io_out_bits_tag; // @[:@54566.4 :@54567.4]
  assign _T_366 = _T_365[7:0]; // @[FringeBundles.scala 114:28:@54568.4]
  assign cmdOutDecoder = 256'h1 << _T_366; // @[OneHot.scala 45:35:@54574.4]
  assign _T_379 = io_app_0_wdata_valid & cmdMux_io_out_valid; // @[StreamArbiter.scala 42:78:@54577.4]
  assign _T_380 = elementCtr_io_out < cmdMux_io_out_bits_size; // @[StreamArbiter.scala 42:121:@54578.4]
  assign _T_395 = io_dram_wresp_bits_tag[7:0]; // @[FringeBundles.scala 140:28:@54765.4]
  assign wrespDecoder = 256'h1 << _T_395; // @[OneHot.scala 45:35:@54772.4]
  assign _T_400 = cmdInDecoder[0]; // @[StreamArbiter.scala 61:55:@54777.4]
  assign _T_403 = cmdOutDecoder[0]; // @[StreamArbiter.scala 62:85:@54781.4]
  assign _T_404 = _T_360 & _T_403; // @[StreamArbiter.scala 62:70:@54782.4]
  assign _T_409 = wrespDecoder[0]; // @[StreamArbiter.scala 67:58:@54806.4]
  assign io_app_0_cmd_ready = cmdMux_io_in_ready & _T_400; // @[StreamArbiter.scala 61:19:@54779.4]
  assign io_app_0_wdata_ready = _T_404 & _T_380; // @[StreamArbiter.scala 62:21:@54785.4]
  assign io_app_0_wresp_valid = io_dram_wresp_valid & _T_409; // @[StreamArbiter.scala 67:21:@54808.4]
  assign io_dram_cmd_valid = cmdMux_io_out_valid; // @[StreamArbiter.scala 46:15:@54668.4]
  assign io_dram_cmd_bits_addr = cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 46:15:@54667.4]
  assign io_dram_cmd_bits_size = cmdMux_io_out_bits_size; // @[StreamArbiter.scala 46:15:@54666.4]
  assign io_dram_cmd_bits_isWr = cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 46:15:@54664.4]
  assign io_dram_cmd_bits_tag = cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 46:15:@54663.4]
  assign io_dram_wdata_valid = wdataMux_io_out_valid; // @[StreamArbiter.scala 47:17:@54751.4]
  assign io_dram_wdata_bits_wdata_0 = wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 47:17:@54735.4]
  assign io_dram_wdata_bits_wdata_1 = wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 47:17:@54736.4]
  assign io_dram_wdata_bits_wdata_2 = wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 47:17:@54737.4]
  assign io_dram_wdata_bits_wdata_3 = wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 47:17:@54738.4]
  assign io_dram_wdata_bits_wdata_4 = wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 47:17:@54739.4]
  assign io_dram_wdata_bits_wdata_5 = wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 47:17:@54740.4]
  assign io_dram_wdata_bits_wdata_6 = wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 47:17:@54741.4]
  assign io_dram_wdata_bits_wdata_7 = wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 47:17:@54742.4]
  assign io_dram_wdata_bits_wdata_8 = wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 47:17:@54743.4]
  assign io_dram_wdata_bits_wdata_9 = wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 47:17:@54744.4]
  assign io_dram_wdata_bits_wdata_10 = wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 47:17:@54745.4]
  assign io_dram_wdata_bits_wdata_11 = wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 47:17:@54746.4]
  assign io_dram_wdata_bits_wdata_12 = wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 47:17:@54747.4]
  assign io_dram_wdata_bits_wdata_13 = wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 47:17:@54748.4]
  assign io_dram_wdata_bits_wdata_14 = wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 47:17:@54749.4]
  assign io_dram_wdata_bits_wdata_15 = wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 47:17:@54750.4]
  assign io_dram_wdata_bits_wstrb_0 = wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 47:17:@54671.4]
  assign io_dram_wdata_bits_wstrb_1 = wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 47:17:@54672.4]
  assign io_dram_wdata_bits_wstrb_2 = wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 47:17:@54673.4]
  assign io_dram_wdata_bits_wstrb_3 = wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 47:17:@54674.4]
  assign io_dram_wdata_bits_wstrb_4 = wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 47:17:@54675.4]
  assign io_dram_wdata_bits_wstrb_5 = wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 47:17:@54676.4]
  assign io_dram_wdata_bits_wstrb_6 = wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 47:17:@54677.4]
  assign io_dram_wdata_bits_wstrb_7 = wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 47:17:@54678.4]
  assign io_dram_wdata_bits_wstrb_8 = wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 47:17:@54679.4]
  assign io_dram_wdata_bits_wstrb_9 = wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 47:17:@54680.4]
  assign io_dram_wdata_bits_wstrb_10 = wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 47:17:@54681.4]
  assign io_dram_wdata_bits_wstrb_11 = wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 47:17:@54682.4]
  assign io_dram_wdata_bits_wstrb_12 = wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 47:17:@54683.4]
  assign io_dram_wdata_bits_wstrb_13 = wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 47:17:@54684.4]
  assign io_dram_wdata_bits_wstrb_14 = wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 47:17:@54685.4]
  assign io_dram_wdata_bits_wstrb_15 = wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 47:17:@54686.4]
  assign io_dram_wdata_bits_wstrb_16 = wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 47:17:@54687.4]
  assign io_dram_wdata_bits_wstrb_17 = wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 47:17:@54688.4]
  assign io_dram_wdata_bits_wstrb_18 = wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 47:17:@54689.4]
  assign io_dram_wdata_bits_wstrb_19 = wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 47:17:@54690.4]
  assign io_dram_wdata_bits_wstrb_20 = wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 47:17:@54691.4]
  assign io_dram_wdata_bits_wstrb_21 = wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 47:17:@54692.4]
  assign io_dram_wdata_bits_wstrb_22 = wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 47:17:@54693.4]
  assign io_dram_wdata_bits_wstrb_23 = wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 47:17:@54694.4]
  assign io_dram_wdata_bits_wstrb_24 = wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 47:17:@54695.4]
  assign io_dram_wdata_bits_wstrb_25 = wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 47:17:@54696.4]
  assign io_dram_wdata_bits_wstrb_26 = wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 47:17:@54697.4]
  assign io_dram_wdata_bits_wstrb_27 = wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 47:17:@54698.4]
  assign io_dram_wdata_bits_wstrb_28 = wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 47:17:@54699.4]
  assign io_dram_wdata_bits_wstrb_29 = wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 47:17:@54700.4]
  assign io_dram_wdata_bits_wstrb_30 = wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 47:17:@54701.4]
  assign io_dram_wdata_bits_wstrb_31 = wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 47:17:@54702.4]
  assign io_dram_wdata_bits_wstrb_32 = wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 47:17:@54703.4]
  assign io_dram_wdata_bits_wstrb_33 = wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 47:17:@54704.4]
  assign io_dram_wdata_bits_wstrb_34 = wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 47:17:@54705.4]
  assign io_dram_wdata_bits_wstrb_35 = wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 47:17:@54706.4]
  assign io_dram_wdata_bits_wstrb_36 = wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 47:17:@54707.4]
  assign io_dram_wdata_bits_wstrb_37 = wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 47:17:@54708.4]
  assign io_dram_wdata_bits_wstrb_38 = wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 47:17:@54709.4]
  assign io_dram_wdata_bits_wstrb_39 = wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 47:17:@54710.4]
  assign io_dram_wdata_bits_wstrb_40 = wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 47:17:@54711.4]
  assign io_dram_wdata_bits_wstrb_41 = wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 47:17:@54712.4]
  assign io_dram_wdata_bits_wstrb_42 = wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 47:17:@54713.4]
  assign io_dram_wdata_bits_wstrb_43 = wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 47:17:@54714.4]
  assign io_dram_wdata_bits_wstrb_44 = wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 47:17:@54715.4]
  assign io_dram_wdata_bits_wstrb_45 = wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 47:17:@54716.4]
  assign io_dram_wdata_bits_wstrb_46 = wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 47:17:@54717.4]
  assign io_dram_wdata_bits_wstrb_47 = wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 47:17:@54718.4]
  assign io_dram_wdata_bits_wstrb_48 = wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 47:17:@54719.4]
  assign io_dram_wdata_bits_wstrb_49 = wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 47:17:@54720.4]
  assign io_dram_wdata_bits_wstrb_50 = wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 47:17:@54721.4]
  assign io_dram_wdata_bits_wstrb_51 = wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 47:17:@54722.4]
  assign io_dram_wdata_bits_wstrb_52 = wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 47:17:@54723.4]
  assign io_dram_wdata_bits_wstrb_53 = wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 47:17:@54724.4]
  assign io_dram_wdata_bits_wstrb_54 = wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 47:17:@54725.4]
  assign io_dram_wdata_bits_wstrb_55 = wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 47:17:@54726.4]
  assign io_dram_wdata_bits_wstrb_56 = wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 47:17:@54727.4]
  assign io_dram_wdata_bits_wstrb_57 = wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 47:17:@54728.4]
  assign io_dram_wdata_bits_wstrb_58 = wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 47:17:@54729.4]
  assign io_dram_wdata_bits_wstrb_59 = wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 47:17:@54730.4]
  assign io_dram_wdata_bits_wstrb_60 = wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 47:17:@54731.4]
  assign io_dram_wdata_bits_wstrb_61 = wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 47:17:@54732.4]
  assign io_dram_wdata_bits_wstrb_62 = wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 47:17:@54733.4]
  assign io_dram_wdata_bits_wstrb_63 = wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 47:17:@54734.4]
  assign io_dram_rresp_ready = io_app_0_rresp_ready; // @[StreamArbiter.scala 72:23:@54812.4]
  assign io_dram_wresp_ready = io_app_0_wresp_ready; // @[StreamArbiter.scala 73:23:@54815.4]
  assign RetimeWrapper_clock = clock; // @[:@54517.4]
  assign RetimeWrapper_reset = reset; // @[:@54518.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@54520.4]
  assign RetimeWrapper_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@54519.4]
  assign RetimeWrapper_1_clock = clock; // @[:@54524.4]
  assign RetimeWrapper_1_reset = reset; // @[:@54525.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@54527.4]
  assign RetimeWrapper_1_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@54526.4]
  assign cmdMux_io_in_valid = io_app_0_cmd_valid; // @[StreamArbiter.scala 26:22:@54536.4]
  assign cmdMux_io_in_bits_0_addr = io_app_0_cmd_bits_addr; // @[StreamArbiter.scala 29:9:@54542.4]
  assign cmdMux_io_in_bits_0_size = io_app_0_cmd_bits_size; // @[StreamArbiter.scala 29:9:@54541.4]
  assign cmdMux_io_in_bits_0_isWr = io_app_0_cmd_bits_isWr; // @[StreamArbiter.scala 29:9:@54539.4]
  assign cmdMux_io_in_bits_0_tag = {_T_358,8'h0}; // @[StreamArbiter.scala 29:9:@54538.4 FringeBundles.scala 115:32:@54555.4]
  assign cmdMux_io_out_ready = io_dram_cmd_valid & io_dram_cmd_ready; // @[StreamArbiter.scala 46:15:@54669.4 StreamArbiter.scala 57:23:@54775.4]
  assign wdataMux_io_in_valid = _T_379 & _T_380; // @[StreamArbiter.scala 42:24:@54580.4]
  assign wdataMux_io_in_bits_0_wdata_0 = io_app_0_wdata_bits_wdata_0; // @[StreamArbiter.scala 44:23:@54647.4]
  assign wdataMux_io_in_bits_0_wdata_1 = io_app_0_wdata_bits_wdata_1; // @[StreamArbiter.scala 44:23:@54648.4]
  assign wdataMux_io_in_bits_0_wdata_2 = io_app_0_wdata_bits_wdata_2; // @[StreamArbiter.scala 44:23:@54649.4]
  assign wdataMux_io_in_bits_0_wdata_3 = io_app_0_wdata_bits_wdata_3; // @[StreamArbiter.scala 44:23:@54650.4]
  assign wdataMux_io_in_bits_0_wdata_4 = io_app_0_wdata_bits_wdata_4; // @[StreamArbiter.scala 44:23:@54651.4]
  assign wdataMux_io_in_bits_0_wdata_5 = io_app_0_wdata_bits_wdata_5; // @[StreamArbiter.scala 44:23:@54652.4]
  assign wdataMux_io_in_bits_0_wdata_6 = io_app_0_wdata_bits_wdata_6; // @[StreamArbiter.scala 44:23:@54653.4]
  assign wdataMux_io_in_bits_0_wdata_7 = io_app_0_wdata_bits_wdata_7; // @[StreamArbiter.scala 44:23:@54654.4]
  assign wdataMux_io_in_bits_0_wdata_8 = io_app_0_wdata_bits_wdata_8; // @[StreamArbiter.scala 44:23:@54655.4]
  assign wdataMux_io_in_bits_0_wdata_9 = io_app_0_wdata_bits_wdata_9; // @[StreamArbiter.scala 44:23:@54656.4]
  assign wdataMux_io_in_bits_0_wdata_10 = io_app_0_wdata_bits_wdata_10; // @[StreamArbiter.scala 44:23:@54657.4]
  assign wdataMux_io_in_bits_0_wdata_11 = io_app_0_wdata_bits_wdata_11; // @[StreamArbiter.scala 44:23:@54658.4]
  assign wdataMux_io_in_bits_0_wdata_12 = io_app_0_wdata_bits_wdata_12; // @[StreamArbiter.scala 44:23:@54659.4]
  assign wdataMux_io_in_bits_0_wdata_13 = io_app_0_wdata_bits_wdata_13; // @[StreamArbiter.scala 44:23:@54660.4]
  assign wdataMux_io_in_bits_0_wdata_14 = io_app_0_wdata_bits_wdata_14; // @[StreamArbiter.scala 44:23:@54661.4]
  assign wdataMux_io_in_bits_0_wdata_15 = io_app_0_wdata_bits_wdata_15; // @[StreamArbiter.scala 44:23:@54662.4]
  assign wdataMux_io_in_bits_0_wstrb_0 = io_app_0_wdata_bits_wstrb_0; // @[StreamArbiter.scala 44:23:@54583.4]
  assign wdataMux_io_in_bits_0_wstrb_1 = io_app_0_wdata_bits_wstrb_1; // @[StreamArbiter.scala 44:23:@54584.4]
  assign wdataMux_io_in_bits_0_wstrb_2 = io_app_0_wdata_bits_wstrb_2; // @[StreamArbiter.scala 44:23:@54585.4]
  assign wdataMux_io_in_bits_0_wstrb_3 = io_app_0_wdata_bits_wstrb_3; // @[StreamArbiter.scala 44:23:@54586.4]
  assign wdataMux_io_in_bits_0_wstrb_4 = io_app_0_wdata_bits_wstrb_4; // @[StreamArbiter.scala 44:23:@54587.4]
  assign wdataMux_io_in_bits_0_wstrb_5 = io_app_0_wdata_bits_wstrb_5; // @[StreamArbiter.scala 44:23:@54588.4]
  assign wdataMux_io_in_bits_0_wstrb_6 = io_app_0_wdata_bits_wstrb_6; // @[StreamArbiter.scala 44:23:@54589.4]
  assign wdataMux_io_in_bits_0_wstrb_7 = io_app_0_wdata_bits_wstrb_7; // @[StreamArbiter.scala 44:23:@54590.4]
  assign wdataMux_io_in_bits_0_wstrb_8 = io_app_0_wdata_bits_wstrb_8; // @[StreamArbiter.scala 44:23:@54591.4]
  assign wdataMux_io_in_bits_0_wstrb_9 = io_app_0_wdata_bits_wstrb_9; // @[StreamArbiter.scala 44:23:@54592.4]
  assign wdataMux_io_in_bits_0_wstrb_10 = io_app_0_wdata_bits_wstrb_10; // @[StreamArbiter.scala 44:23:@54593.4]
  assign wdataMux_io_in_bits_0_wstrb_11 = io_app_0_wdata_bits_wstrb_11; // @[StreamArbiter.scala 44:23:@54594.4]
  assign wdataMux_io_in_bits_0_wstrb_12 = io_app_0_wdata_bits_wstrb_12; // @[StreamArbiter.scala 44:23:@54595.4]
  assign wdataMux_io_in_bits_0_wstrb_13 = io_app_0_wdata_bits_wstrb_13; // @[StreamArbiter.scala 44:23:@54596.4]
  assign wdataMux_io_in_bits_0_wstrb_14 = io_app_0_wdata_bits_wstrb_14; // @[StreamArbiter.scala 44:23:@54597.4]
  assign wdataMux_io_in_bits_0_wstrb_15 = io_app_0_wdata_bits_wstrb_15; // @[StreamArbiter.scala 44:23:@54598.4]
  assign wdataMux_io_in_bits_0_wstrb_16 = io_app_0_wdata_bits_wstrb_16; // @[StreamArbiter.scala 44:23:@54599.4]
  assign wdataMux_io_in_bits_0_wstrb_17 = io_app_0_wdata_bits_wstrb_17; // @[StreamArbiter.scala 44:23:@54600.4]
  assign wdataMux_io_in_bits_0_wstrb_18 = io_app_0_wdata_bits_wstrb_18; // @[StreamArbiter.scala 44:23:@54601.4]
  assign wdataMux_io_in_bits_0_wstrb_19 = io_app_0_wdata_bits_wstrb_19; // @[StreamArbiter.scala 44:23:@54602.4]
  assign wdataMux_io_in_bits_0_wstrb_20 = io_app_0_wdata_bits_wstrb_20; // @[StreamArbiter.scala 44:23:@54603.4]
  assign wdataMux_io_in_bits_0_wstrb_21 = io_app_0_wdata_bits_wstrb_21; // @[StreamArbiter.scala 44:23:@54604.4]
  assign wdataMux_io_in_bits_0_wstrb_22 = io_app_0_wdata_bits_wstrb_22; // @[StreamArbiter.scala 44:23:@54605.4]
  assign wdataMux_io_in_bits_0_wstrb_23 = io_app_0_wdata_bits_wstrb_23; // @[StreamArbiter.scala 44:23:@54606.4]
  assign wdataMux_io_in_bits_0_wstrb_24 = io_app_0_wdata_bits_wstrb_24; // @[StreamArbiter.scala 44:23:@54607.4]
  assign wdataMux_io_in_bits_0_wstrb_25 = io_app_0_wdata_bits_wstrb_25; // @[StreamArbiter.scala 44:23:@54608.4]
  assign wdataMux_io_in_bits_0_wstrb_26 = io_app_0_wdata_bits_wstrb_26; // @[StreamArbiter.scala 44:23:@54609.4]
  assign wdataMux_io_in_bits_0_wstrb_27 = io_app_0_wdata_bits_wstrb_27; // @[StreamArbiter.scala 44:23:@54610.4]
  assign wdataMux_io_in_bits_0_wstrb_28 = io_app_0_wdata_bits_wstrb_28; // @[StreamArbiter.scala 44:23:@54611.4]
  assign wdataMux_io_in_bits_0_wstrb_29 = io_app_0_wdata_bits_wstrb_29; // @[StreamArbiter.scala 44:23:@54612.4]
  assign wdataMux_io_in_bits_0_wstrb_30 = io_app_0_wdata_bits_wstrb_30; // @[StreamArbiter.scala 44:23:@54613.4]
  assign wdataMux_io_in_bits_0_wstrb_31 = io_app_0_wdata_bits_wstrb_31; // @[StreamArbiter.scala 44:23:@54614.4]
  assign wdataMux_io_in_bits_0_wstrb_32 = io_app_0_wdata_bits_wstrb_32; // @[StreamArbiter.scala 44:23:@54615.4]
  assign wdataMux_io_in_bits_0_wstrb_33 = io_app_0_wdata_bits_wstrb_33; // @[StreamArbiter.scala 44:23:@54616.4]
  assign wdataMux_io_in_bits_0_wstrb_34 = io_app_0_wdata_bits_wstrb_34; // @[StreamArbiter.scala 44:23:@54617.4]
  assign wdataMux_io_in_bits_0_wstrb_35 = io_app_0_wdata_bits_wstrb_35; // @[StreamArbiter.scala 44:23:@54618.4]
  assign wdataMux_io_in_bits_0_wstrb_36 = io_app_0_wdata_bits_wstrb_36; // @[StreamArbiter.scala 44:23:@54619.4]
  assign wdataMux_io_in_bits_0_wstrb_37 = io_app_0_wdata_bits_wstrb_37; // @[StreamArbiter.scala 44:23:@54620.4]
  assign wdataMux_io_in_bits_0_wstrb_38 = io_app_0_wdata_bits_wstrb_38; // @[StreamArbiter.scala 44:23:@54621.4]
  assign wdataMux_io_in_bits_0_wstrb_39 = io_app_0_wdata_bits_wstrb_39; // @[StreamArbiter.scala 44:23:@54622.4]
  assign wdataMux_io_in_bits_0_wstrb_40 = io_app_0_wdata_bits_wstrb_40; // @[StreamArbiter.scala 44:23:@54623.4]
  assign wdataMux_io_in_bits_0_wstrb_41 = io_app_0_wdata_bits_wstrb_41; // @[StreamArbiter.scala 44:23:@54624.4]
  assign wdataMux_io_in_bits_0_wstrb_42 = io_app_0_wdata_bits_wstrb_42; // @[StreamArbiter.scala 44:23:@54625.4]
  assign wdataMux_io_in_bits_0_wstrb_43 = io_app_0_wdata_bits_wstrb_43; // @[StreamArbiter.scala 44:23:@54626.4]
  assign wdataMux_io_in_bits_0_wstrb_44 = io_app_0_wdata_bits_wstrb_44; // @[StreamArbiter.scala 44:23:@54627.4]
  assign wdataMux_io_in_bits_0_wstrb_45 = io_app_0_wdata_bits_wstrb_45; // @[StreamArbiter.scala 44:23:@54628.4]
  assign wdataMux_io_in_bits_0_wstrb_46 = io_app_0_wdata_bits_wstrb_46; // @[StreamArbiter.scala 44:23:@54629.4]
  assign wdataMux_io_in_bits_0_wstrb_47 = io_app_0_wdata_bits_wstrb_47; // @[StreamArbiter.scala 44:23:@54630.4]
  assign wdataMux_io_in_bits_0_wstrb_48 = io_app_0_wdata_bits_wstrb_48; // @[StreamArbiter.scala 44:23:@54631.4]
  assign wdataMux_io_in_bits_0_wstrb_49 = io_app_0_wdata_bits_wstrb_49; // @[StreamArbiter.scala 44:23:@54632.4]
  assign wdataMux_io_in_bits_0_wstrb_50 = io_app_0_wdata_bits_wstrb_50; // @[StreamArbiter.scala 44:23:@54633.4]
  assign wdataMux_io_in_bits_0_wstrb_51 = io_app_0_wdata_bits_wstrb_51; // @[StreamArbiter.scala 44:23:@54634.4]
  assign wdataMux_io_in_bits_0_wstrb_52 = io_app_0_wdata_bits_wstrb_52; // @[StreamArbiter.scala 44:23:@54635.4]
  assign wdataMux_io_in_bits_0_wstrb_53 = io_app_0_wdata_bits_wstrb_53; // @[StreamArbiter.scala 44:23:@54636.4]
  assign wdataMux_io_in_bits_0_wstrb_54 = io_app_0_wdata_bits_wstrb_54; // @[StreamArbiter.scala 44:23:@54637.4]
  assign wdataMux_io_in_bits_0_wstrb_55 = io_app_0_wdata_bits_wstrb_55; // @[StreamArbiter.scala 44:23:@54638.4]
  assign wdataMux_io_in_bits_0_wstrb_56 = io_app_0_wdata_bits_wstrb_56; // @[StreamArbiter.scala 44:23:@54639.4]
  assign wdataMux_io_in_bits_0_wstrb_57 = io_app_0_wdata_bits_wstrb_57; // @[StreamArbiter.scala 44:23:@54640.4]
  assign wdataMux_io_in_bits_0_wstrb_58 = io_app_0_wdata_bits_wstrb_58; // @[StreamArbiter.scala 44:23:@54641.4]
  assign wdataMux_io_in_bits_0_wstrb_59 = io_app_0_wdata_bits_wstrb_59; // @[StreamArbiter.scala 44:23:@54642.4]
  assign wdataMux_io_in_bits_0_wstrb_60 = io_app_0_wdata_bits_wstrb_60; // @[StreamArbiter.scala 44:23:@54643.4]
  assign wdataMux_io_in_bits_0_wstrb_61 = io_app_0_wdata_bits_wstrb_61; // @[StreamArbiter.scala 44:23:@54644.4]
  assign wdataMux_io_in_bits_0_wstrb_62 = io_app_0_wdata_bits_wstrb_62; // @[StreamArbiter.scala 44:23:@54645.4]
  assign wdataMux_io_in_bits_0_wstrb_63 = io_app_0_wdata_bits_wstrb_63; // @[StreamArbiter.scala 44:23:@54646.4]
  assign wdataMux_io_out_ready = io_dram_wdata_valid & io_dram_wdata_ready; // @[StreamArbiter.scala 47:17:@54752.4 StreamArbiter.scala 58:25:@54776.4]
  assign elementCtr_clock = clock; // @[:@54560.4]
  assign elementCtr_reset = reset; // @[:@54561.4]
  assign elementCtr_io_reset = cmdMux_io_out_ready; // @[StreamArbiter.scala 38:23:@54564.4]
  assign elementCtr_io_enable = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:24:@54563.4]
endmodule
module Counter_72( // @[:@54817.2]
  input         clock, // @[:@54818.4]
  input         reset, // @[:@54819.4]
  input         io_reset, // @[:@54820.4]
  input         io_enable, // @[:@54820.4]
  input  [31:0] io_stride, // @[:@54820.4]
  output [31:0] io_out, // @[:@54820.4]
  output [31:0] io_next // @[:@54820.4]
);
  reg [31:0] count; // @[Counter.scala 15:22:@54822.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_17; // @[Counter.scala 17:24:@54823.4]
  wire [31:0] newCount; // @[Counter.scala 17:24:@54824.4]
  wire [31:0] _GEN_0; // @[Counter.scala 21:26:@54829.6]
  wire [31:0] _GEN_1; // @[Counter.scala 19:18:@54825.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@54823.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@54824.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@54829.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 19:18:@54825.4]
  assign io_out = count; // @[Counter.scala 25:10:@54832.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@54833.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module AXICmdSplit( // @[:@54835.2]
  input         clock, // @[:@54836.4]
  input         reset, // @[:@54837.4]
  output        io_in_cmd_ready, // @[:@54838.4]
  input         io_in_cmd_valid, // @[:@54838.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@54838.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@54838.4]
  input         io_in_cmd_bits_isWr, // @[:@54838.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@54838.4]
  output        io_in_wdata_ready, // @[:@54838.4]
  input         io_in_wdata_valid, // @[:@54838.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@54838.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@54838.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@54838.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@54838.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@54838.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@54838.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@54838.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@54838.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@54838.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@54838.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@54838.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@54838.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@54838.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@54838.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@54838.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@54838.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@54838.4]
  input         io_in_rresp_ready, // @[:@54838.4]
  input         io_in_wresp_ready, // @[:@54838.4]
  output        io_in_wresp_valid, // @[:@54838.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@54838.4]
  input         io_out_cmd_ready, // @[:@54838.4]
  output        io_out_cmd_valid, // @[:@54838.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@54838.4]
  output [31:0] io_out_cmd_bits_size, // @[:@54838.4]
  output        io_out_cmd_bits_isWr, // @[:@54838.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@54838.4]
  input         io_out_wdata_ready, // @[:@54838.4]
  output        io_out_wdata_valid, // @[:@54838.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@54838.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@54838.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@54838.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@54838.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@54838.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@54838.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@54838.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@54838.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@54838.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@54838.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@54838.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@54838.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@54838.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@54838.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@54838.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@54838.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@54838.4]
  output        io_out_rresp_ready, // @[:@54838.4]
  output        io_out_wresp_ready, // @[:@54838.4]
  input         io_out_wresp_valid, // @[:@54838.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@54838.4]
);
  wire  cmdSizeCounter_clock; // @[AXIProtocol.scala 18:30:@54952.4]
  wire  cmdSizeCounter_reset; // @[AXIProtocol.scala 18:30:@54952.4]
  wire  cmdSizeCounter_io_reset; // @[AXIProtocol.scala 18:30:@54952.4]
  wire  cmdSizeCounter_io_enable; // @[AXIProtocol.scala 18:30:@54952.4]
  wire [31:0] cmdSizeCounter_io_stride; // @[AXIProtocol.scala 18:30:@54952.4]
  wire [31:0] cmdSizeCounter_io_out; // @[AXIProtocol.scala 18:30:@54952.4]
  wire [31:0] cmdSizeCounter_io_next; // @[AXIProtocol.scala 18:30:@54952.4]
  wire [32:0] _T_199; // @[AXIProtocol.scala 20:46:@54955.4]
  wire [32:0] _T_200; // @[AXIProtocol.scala 20:46:@54956.4]
  wire [31:0] cmdSizeRemaining; // @[AXIProtocol.scala 20:46:@54957.4]
  wire  lastCmd; // @[AXIProtocol.scala 23:35:@54958.4]
  wire [37:0] _GEN_0; // @[AXIProtocol.scala 27:47:@54961.4]
  wire [37:0] addrOffsetBytes; // @[AXIProtocol.scala 27:47:@54961.4]
  wire [63:0] _GEN_1; // @[AXIProtocol.scala 28:49:@54962.4]
  wire [64:0] _T_201; // @[AXIProtocol.scala 28:49:@54962.4]
  wire [63:0] cmdAddr_bits; // @[AXIProtocol.scala 28:49:@54963.4]
  wire [57:0] _T_204; // @[FringeBundles.scala 158:22:@54966.4]
  wire [7:0] cmdTag_streamID; // @[FringeBundles.scala 114:28:@54973.4]
  wire [22:0] cmdTag_uid; // @[FringeBundles.scala 114:28:@54977.4]
  wire [23:0] _T_214; // @[FringeBundles.scala 115:37:@54980.4]
  wire  cmdIssue; // @[AXIProtocol.scala 36:35:@54983.4]
  wire  _T_223; // @[FringeBundles.scala 140:28:@54994.4]
  Counter_72 cmdSizeCounter ( // @[AXIProtocol.scala 18:30:@54952.4]
    .clock(cmdSizeCounter_clock),
    .reset(cmdSizeCounter_reset),
    .io_reset(cmdSizeCounter_io_reset),
    .io_enable(cmdSizeCounter_io_enable),
    .io_stride(cmdSizeCounter_io_stride),
    .io_out(cmdSizeCounter_io_out),
    .io_next(cmdSizeCounter_io_next)
  );
  assign _T_199 = io_in_cmd_bits_size - cmdSizeCounter_io_out; // @[AXIProtocol.scala 20:46:@54955.4]
  assign _T_200 = $unsigned(_T_199); // @[AXIProtocol.scala 20:46:@54956.4]
  assign cmdSizeRemaining = _T_200[31:0]; // @[AXIProtocol.scala 20:46:@54957.4]
  assign lastCmd = cmdSizeRemaining <= 32'h100; // @[AXIProtocol.scala 23:35:@54958.4]
  assign _GEN_0 = {{6'd0}, cmdSizeCounter_io_out}; // @[AXIProtocol.scala 27:47:@54961.4]
  assign addrOffsetBytes = _GEN_0 << 6; // @[AXIProtocol.scala 27:47:@54961.4]
  assign _GEN_1 = {{26'd0}, addrOffsetBytes}; // @[AXIProtocol.scala 28:49:@54962.4]
  assign _T_201 = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@54962.4]
  assign cmdAddr_bits = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@54963.4]
  assign _T_204 = cmdAddr_bits[63:6]; // @[FringeBundles.scala 158:22:@54966.4]
  assign cmdTag_streamID = io_in_cmd_bits_tag[7:0]; // @[FringeBundles.scala 114:28:@54973.4]
  assign cmdTag_uid = io_in_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@54977.4]
  assign _T_214 = {cmdTag_uid,lastCmd}; // @[FringeBundles.scala 115:37:@54980.4]
  assign cmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 36:35:@54983.4]
  assign _T_223 = io_out_wresp_bits_tag[8]; // @[FringeBundles.scala 140:28:@54994.4]
  assign io_in_cmd_ready = lastCmd & cmdIssue; // @[AXIProtocol.scala 15:10:@54951.4 AXIProtocol.scala 38:19:@54985.4]
  assign io_in_wdata_ready = io_out_wdata_ready; // @[AXIProtocol.scala 15:10:@54944.4]
  assign io_in_wresp_valid = io_out_wresp_valid & _T_223; // @[AXIProtocol.scala 15:10:@54841.4 AXIProtocol.scala 46:21:@54999.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 15:10:@54840.4]
  assign io_out_cmd_valid = io_in_cmd_valid; // @[AXIProtocol.scala 15:10:@54950.4]
  assign io_out_cmd_bits_addr = {_T_204,6'h0}; // @[AXIProtocol.scala 15:10:@54949.4 AXIProtocol.scala 29:24:@54968.4]
  assign io_out_cmd_bits_size = lastCmd ? cmdSizeRemaining : 32'h100; // @[AXIProtocol.scala 15:10:@54948.4 AXIProtocol.scala 25:24:@54960.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 15:10:@54946.4]
  assign io_out_cmd_bits_tag = {_T_214,cmdTag_streamID}; // @[AXIProtocol.scala 15:10:@54945.4 FringeBundles.scala 115:32:@54982.4]
  assign io_out_wdata_valid = io_in_wdata_valid; // @[AXIProtocol.scala 15:10:@54943.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 15:10:@54927.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 15:10:@54928.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 15:10:@54929.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 15:10:@54930.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 15:10:@54931.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 15:10:@54932.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 15:10:@54933.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 15:10:@54934.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 15:10:@54935.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 15:10:@54936.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 15:10:@54937.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 15:10:@54938.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 15:10:@54939.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 15:10:@54940.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 15:10:@54941.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 15:10:@54942.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 15:10:@54863.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 15:10:@54864.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 15:10:@54865.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 15:10:@54866.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 15:10:@54867.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 15:10:@54868.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 15:10:@54869.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 15:10:@54870.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 15:10:@54871.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 15:10:@54872.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 15:10:@54873.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 15:10:@54874.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 15:10:@54875.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 15:10:@54876.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 15:10:@54877.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 15:10:@54878.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 15:10:@54879.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 15:10:@54880.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 15:10:@54881.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 15:10:@54882.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 15:10:@54883.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 15:10:@54884.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 15:10:@54885.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 15:10:@54886.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 15:10:@54887.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 15:10:@54888.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 15:10:@54889.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 15:10:@54890.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 15:10:@54891.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 15:10:@54892.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 15:10:@54893.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 15:10:@54894.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 15:10:@54895.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 15:10:@54896.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 15:10:@54897.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 15:10:@54898.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 15:10:@54899.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 15:10:@54900.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 15:10:@54901.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 15:10:@54902.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 15:10:@54903.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 15:10:@54904.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 15:10:@54905.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 15:10:@54906.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 15:10:@54907.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 15:10:@54908.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 15:10:@54909.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 15:10:@54910.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 15:10:@54911.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 15:10:@54912.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 15:10:@54913.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 15:10:@54914.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 15:10:@54915.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 15:10:@54916.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 15:10:@54917.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 15:10:@54918.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 15:10:@54919.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 15:10:@54920.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 15:10:@54921.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 15:10:@54922.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 15:10:@54923.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 15:10:@54924.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 15:10:@54925.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 15:10:@54926.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 15:10:@54861.4]
  assign io_out_wresp_ready = _T_223 ? io_in_wresp_ready : 1'h1; // @[AXIProtocol.scala 15:10:@54842.4 AXIProtocol.scala 47:22:@55001.4]
  assign cmdSizeCounter_clock = clock; // @[:@54953.4]
  assign cmdSizeCounter_reset = reset; // @[:@54954.4]
  assign cmdSizeCounter_io_reset = lastCmd & cmdIssue; // @[AXIProtocol.scala 40:27:@54986.4]
  assign cmdSizeCounter_io_enable = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 41:28:@54987.4]
  assign cmdSizeCounter_io_stride = 32'h100; // @[AXIProtocol.scala 42:28:@54988.4]
endmodule
module AXICmdIssue( // @[:@55021.2]
  input         clock, // @[:@55022.4]
  input         reset, // @[:@55023.4]
  output        io_in_cmd_ready, // @[:@55024.4]
  input         io_in_cmd_valid, // @[:@55024.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@55024.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@55024.4]
  input         io_in_cmd_bits_isWr, // @[:@55024.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@55024.4]
  output        io_in_wdata_ready, // @[:@55024.4]
  input         io_in_wdata_valid, // @[:@55024.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@55024.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@55024.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@55024.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@55024.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@55024.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@55024.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@55024.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@55024.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@55024.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@55024.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@55024.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@55024.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@55024.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@55024.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@55024.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@55024.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@55024.4]
  input         io_in_rresp_ready, // @[:@55024.4]
  input         io_in_wresp_ready, // @[:@55024.4]
  output        io_in_wresp_valid, // @[:@55024.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@55024.4]
  input         io_out_cmd_ready, // @[:@55024.4]
  output        io_out_cmd_valid, // @[:@55024.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@55024.4]
  output [31:0] io_out_cmd_bits_size, // @[:@55024.4]
  output        io_out_cmd_bits_isWr, // @[:@55024.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@55024.4]
  input         io_out_wdata_ready, // @[:@55024.4]
  output        io_out_wdata_valid, // @[:@55024.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@55024.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@55024.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@55024.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@55024.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@55024.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@55024.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@55024.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@55024.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@55024.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@55024.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@55024.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@55024.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@55024.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@55024.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@55024.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@55024.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@55024.4]
  output        io_out_wdata_bits_wlast, // @[:@55024.4]
  output        io_out_rresp_ready, // @[:@55024.4]
  output        io_out_wresp_ready, // @[:@55024.4]
  input         io_out_wresp_valid, // @[:@55024.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@55024.4]
);
  wire  wdataCounter_clock; // @[AXIProtocol.scala 59:28:@55138.4]
  wire  wdataCounter_reset; // @[AXIProtocol.scala 59:28:@55138.4]
  wire  wdataCounter_io_reset; // @[AXIProtocol.scala 59:28:@55138.4]
  wire  wdataCounter_io_enable; // @[AXIProtocol.scala 59:28:@55138.4]
  wire [31:0] wdataCounter_io_stride; // @[AXIProtocol.scala 59:28:@55138.4]
  wire [31:0] wdataCounter_io_out; // @[AXIProtocol.scala 59:28:@55138.4]
  wire [31:0] wdataCounter_io_next; // @[AXIProtocol.scala 59:28:@55138.4]
  reg  writeIssued; // @[AXIProtocol.scala 61:28:@55141.4]
  reg [31:0] _RAND_0;
  wire  dramCmdIssue; // @[AXIProtocol.scala 63:39:@55142.4]
  wire  dramWriteIssue; // @[AXIProtocol.scala 64:43:@55143.4]
  wire  _T_201; // @[AXIProtocol.scala 68:54:@55144.4]
  wire  wlast; // @[AXIProtocol.scala 68:30:@55145.4]
  wire  _T_203; // @[AXIProtocol.scala 72:28:@55151.6]
  wire  _GEN_0; // @[AXIProtocol.scala 72:40:@55152.6]
  wire  _GEN_1; // @[AXIProtocol.scala 70:15:@55147.4]
  wire  _T_208; // @[AXIProtocol.scala 84:55:@55161.4]
  wire  _T_210; // @[AXIProtocol.scala 84:44:@55162.4]
  Counter_72 wdataCounter ( // @[AXIProtocol.scala 59:28:@55138.4]
    .clock(wdataCounter_clock),
    .reset(wdataCounter_reset),
    .io_reset(wdataCounter_io_reset),
    .io_enable(wdataCounter_io_enable),
    .io_stride(wdataCounter_io_stride),
    .io_out(wdataCounter_io_out),
    .io_next(wdataCounter_io_next)
  );
  assign dramCmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 63:39:@55142.4]
  assign dramWriteIssue = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 64:43:@55143.4]
  assign _T_201 = wdataCounter_io_next == io_in_cmd_bits_size; // @[AXIProtocol.scala 68:54:@55144.4]
  assign wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 68:30:@55145.4]
  assign _T_203 = dramCmdIssue & io_in_cmd_bits_isWr; // @[AXIProtocol.scala 72:28:@55151.6]
  assign _GEN_0 = _T_203 ? 1'h1 : writeIssued; // @[AXIProtocol.scala 72:40:@55152.6]
  assign _GEN_1 = wlast ? 1'h0 : _GEN_0; // @[AXIProtocol.scala 70:15:@55147.4]
  assign _T_208 = writeIssued == 1'h0; // @[AXIProtocol.scala 84:55:@55161.4]
  assign _T_210 = io_in_cmd_bits_isWr ? _T_208 : 1'h1; // @[AXIProtocol.scala 84:44:@55162.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? wlast : dramCmdIssue; // @[AXIProtocol.scala 56:10:@55137.4 AXIProtocol.scala 81:19:@55159.4]
  assign io_in_wdata_ready = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 56:10:@55130.4 AXIProtocol.scala 82:21:@55160.4]
  assign io_in_wresp_valid = io_out_wresp_valid; // @[AXIProtocol.scala 56:10:@55027.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 56:10:@55026.4]
  assign io_out_cmd_valid = io_in_cmd_valid & _T_210; // @[AXIProtocol.scala 56:10:@55136.4 AXIProtocol.scala 84:20:@55164.4]
  assign io_out_cmd_bits_addr = io_in_cmd_bits_addr; // @[AXIProtocol.scala 56:10:@55135.4]
  assign io_out_cmd_bits_size = io_in_cmd_bits_size; // @[AXIProtocol.scala 56:10:@55134.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 56:10:@55132.4]
  assign io_out_cmd_bits_tag = io_in_cmd_bits_tag; // @[AXIProtocol.scala 56:10:@55131.4]
  assign io_out_wdata_valid = io_in_wdata_valid & writeIssued; // @[AXIProtocol.scala 56:10:@55129.4 AXIProtocol.scala 86:22:@55166.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 56:10:@55113.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 56:10:@55114.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 56:10:@55115.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 56:10:@55116.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 56:10:@55117.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 56:10:@55118.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 56:10:@55119.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 56:10:@55120.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 56:10:@55121.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 56:10:@55122.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 56:10:@55123.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 56:10:@55124.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 56:10:@55125.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 56:10:@55126.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 56:10:@55127.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 56:10:@55128.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 56:10:@55049.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 56:10:@55050.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 56:10:@55051.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 56:10:@55052.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 56:10:@55053.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 56:10:@55054.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 56:10:@55055.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 56:10:@55056.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 56:10:@55057.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 56:10:@55058.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 56:10:@55059.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 56:10:@55060.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 56:10:@55061.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 56:10:@55062.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 56:10:@55063.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 56:10:@55064.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 56:10:@55065.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 56:10:@55066.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 56:10:@55067.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 56:10:@55068.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 56:10:@55069.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 56:10:@55070.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 56:10:@55071.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 56:10:@55072.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 56:10:@55073.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 56:10:@55074.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 56:10:@55075.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 56:10:@55076.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 56:10:@55077.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 56:10:@55078.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 56:10:@55079.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 56:10:@55080.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 56:10:@55081.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 56:10:@55082.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 56:10:@55083.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 56:10:@55084.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 56:10:@55085.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 56:10:@55086.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 56:10:@55087.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 56:10:@55088.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 56:10:@55089.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 56:10:@55090.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 56:10:@55091.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 56:10:@55092.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 56:10:@55093.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 56:10:@55094.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 56:10:@55095.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 56:10:@55096.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 56:10:@55097.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 56:10:@55098.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 56:10:@55099.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 56:10:@55100.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 56:10:@55101.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 56:10:@55102.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 56:10:@55103.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 56:10:@55104.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 56:10:@55105.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 56:10:@55106.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 56:10:@55107.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 56:10:@55108.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 56:10:@55109.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 56:10:@55110.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 56:10:@55111.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 56:10:@55112.4]
  assign io_out_wdata_bits_wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 56:10:@55048.4 AXIProtocol.scala 87:27:@55167.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 56:10:@55047.4]
  assign io_out_wresp_ready = io_in_wresp_ready; // @[AXIProtocol.scala 56:10:@55028.4]
  assign wdataCounter_clock = clock; // @[:@55139.4]
  assign wdataCounter_reset = reset; // @[:@55140.4]
  assign wdataCounter_io_reset = dramWriteIssue & _T_201; // @[AXIProtocol.scala 76:25:@55155.4]
  assign wdataCounter_io_enable = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 77:26:@55156.4]
  assign wdataCounter_io_stride = 32'h1; // @[AXIProtocol.scala 78:26:@55157.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeIssued = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      writeIssued <= 1'h0;
    end else begin
      if (wlast) begin
        writeIssued <= 1'h0;
      end else begin
        if (_T_203) begin
          writeIssued <= 1'h1;
        end
      end
    end
  end
endmodule
module DRAMArbiter( // @[:@55169.2]
  input         clock, // @[:@55170.4]
  input         reset, // @[:@55171.4]
  input         io_enable, // @[:@55172.4]
  output        io_app_stores_0_cmd_ready, // @[:@55172.4]
  input         io_app_stores_0_cmd_valid, // @[:@55172.4]
  input  [63:0] io_app_stores_0_cmd_bits_addr, // @[:@55172.4]
  input  [31:0] io_app_stores_0_cmd_bits_size, // @[:@55172.4]
  output        io_app_stores_0_data_ready, // @[:@55172.4]
  input         io_app_stores_0_data_valid, // @[:@55172.4]
  input  [31:0] io_app_stores_0_data_bits_wdata_0, // @[:@55172.4]
  input         io_app_stores_0_data_bits_wstrb, // @[:@55172.4]
  input         io_app_stores_0_wresp_ready, // @[:@55172.4]
  output        io_app_stores_0_wresp_valid, // @[:@55172.4]
  output        io_app_stores_0_wresp_bits, // @[:@55172.4]
  input         io_dram_cmd_ready, // @[:@55172.4]
  output        io_dram_cmd_valid, // @[:@55172.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@55172.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@55172.4]
  output        io_dram_cmd_bits_isWr, // @[:@55172.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@55172.4]
  input         io_dram_wdata_ready, // @[:@55172.4]
  output        io_dram_wdata_valid, // @[:@55172.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@55172.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@55172.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@55172.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@55172.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@55172.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@55172.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@55172.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@55172.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@55172.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@55172.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@55172.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@55172.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@55172.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@55172.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@55172.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@55172.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@55172.4]
  output        io_dram_wdata_bits_wlast, // @[:@55172.4]
  output        io_dram_rresp_ready, // @[:@55172.4]
  output        io_dram_wresp_ready, // @[:@55172.4]
  input         io_dram_wresp_valid, // @[:@55172.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@55172.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@56058.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@56072.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@56300.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@56415.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@56415.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@56058.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@56072.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@56300.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@56415.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_app_stores_0_cmd_ready = StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 68:18:@56071.4]
  assign io_app_stores_0_data_ready = StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 68:18:@56067.4]
  assign io_app_stores_0_wresp_valid = StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 68:18:@56062.4]
  assign io_app_stores_0_wresp_bits = StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 68:18:@56061.4]
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@56640.4 DRAMArbiter.scala 100:23:@56643.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@56639.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@56638.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@56636.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@56635.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@56633.4 DRAMArbiter.scala 101:25:@56645.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@56617.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@56618.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@56619.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@56620.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@56621.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@56622.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@56623.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@56624.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@56625.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@56626.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@56627.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@56628.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@56629.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@56630.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@56631.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@56632.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@56553.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@56554.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@56555.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@56556.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@56557.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@56558.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@56559.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@56560.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@56561.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@56562.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@56563.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@56564.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@56565.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@56566.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@56567.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@56568.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@56569.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@56570.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@56571.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@56572.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@56573.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@56574.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@56575.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@56576.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@56577.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@56578.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@56579.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@56580.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@56581.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@56582.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@56583.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@56584.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@56585.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@56586.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@56587.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@56588.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@56589.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@56590.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@56591.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@56592.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@56593.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@56594.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@56595.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@56596.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@56597.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@56598.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@56599.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@56600.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@56601.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@56602.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@56603.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@56604.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@56605.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@56606.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@56607.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@56608.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@56609.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@56610.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@56611.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@56612.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@56613.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@56614.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@56615.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@56616.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@56552.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@56551.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@56532.4]
  assign StreamControllerStore_clock = clock; // @[:@56059.4]
  assign StreamControllerStore_reset = reset; // @[:@56060.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@56187.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@56180.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@56077.4]
  assign StreamControllerStore_io_store_cmd_valid = io_app_stores_0_cmd_valid; // @[DRAMArbiter.scala 68:18:@56070.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = io_app_stores_0_cmd_bits_addr; // @[DRAMArbiter.scala 68:18:@56069.4]
  assign StreamControllerStore_io_store_cmd_bits_size = io_app_stores_0_cmd_bits_size; // @[DRAMArbiter.scala 68:18:@56068.4]
  assign StreamControllerStore_io_store_data_valid = io_app_stores_0_data_valid; // @[DRAMArbiter.scala 68:18:@56066.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = io_app_stores_0_data_bits_wdata_0; // @[DRAMArbiter.scala 68:18:@56065.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = io_app_stores_0_data_bits_wstrb; // @[DRAMArbiter.scala 68:18:@56064.4]
  assign StreamControllerStore_io_store_wresp_ready = io_app_stores_0_wresp_ready; // @[DRAMArbiter.scala 68:18:@56063.4]
  assign StreamArbiter_clock = clock; // @[:@56073.4]
  assign StreamArbiter_reset = reset; // @[:@56074.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@56298.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@56297.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@56296.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@56294.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@56293.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@56291.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@56275.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@56276.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@56277.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@56278.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@56279.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@56280.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@56281.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@56282.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@56283.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@56284.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@56285.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@56286.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@56287.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@56288.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@56289.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@56290.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@56211.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@56212.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@56213.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@56214.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@56215.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@56216.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@56217.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@56218.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@56219.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@56220.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@56221.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@56222.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@56223.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@56224.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@56225.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@56226.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@56227.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@56228.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@56229.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@56230.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@56231.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@56232.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@56233.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@56234.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@56235.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@56236.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@56237.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@56238.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@56239.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@56240.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@56241.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@56242.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@56243.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@56244.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@56245.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@56246.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@56247.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@56248.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@56249.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@56250.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@56251.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@56252.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@56253.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@56254.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@56255.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@56256.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@56257.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@56258.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@56259.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@56260.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@56261.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@56262.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@56263.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@56264.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@56265.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@56266.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@56267.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@56268.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@56269.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@56270.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@56271.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@56272.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@56273.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@56274.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@56209.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@56190.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@56414.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@56407.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@56304.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@56303.4]
  assign AXICmdSplit_clock = clock; // @[:@56301.4]
  assign AXICmdSplit_reset = reset; // @[:@56302.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@56413.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@56412.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@56411.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@56409.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@56408.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@56406.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@56390.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@56391.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@56392.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@56393.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@56394.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@56395.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@56396.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@56397.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@56398.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@56399.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@56400.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@56401.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@56402.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@56403.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@56404.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@56405.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@56326.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@56327.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@56328.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@56329.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@56330.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@56331.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@56332.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@56333.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@56334.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@56335.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@56336.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@56337.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@56338.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@56339.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@56340.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@56341.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@56342.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@56343.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@56344.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@56345.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@56346.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@56347.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@56348.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@56349.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@56350.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@56351.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@56352.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@56353.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@56354.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@56355.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@56356.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@56357.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@56358.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@56359.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@56360.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@56361.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@56362.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@56363.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@56364.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@56365.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@56366.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@56367.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@56368.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@56369.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@56370.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@56371.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@56372.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@56373.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@56374.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@56375.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@56376.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@56377.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@56378.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@56379.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@56380.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@56381.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@56382.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@56383.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@56384.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@56385.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@56386.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@56387.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@56388.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@56389.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@56324.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@56305.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@56529.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@56522.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@56419.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@56418.4]
  assign AXICmdIssue_clock = clock; // @[:@56416.4]
  assign AXICmdIssue_reset = reset; // @[:@56417.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@56528.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@56527.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@56526.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@56524.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@56523.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@56521.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@56505.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@56506.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@56507.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@56508.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@56509.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@56510.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@56511.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@56512.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@56513.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@56514.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@56515.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@56516.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@56517.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@56518.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@56519.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@56520.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@56441.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@56442.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@56443.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@56444.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@56445.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@56446.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@56447.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@56448.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@56449.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@56450.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@56451.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@56452.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@56453.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@56454.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@56455.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@56456.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@56457.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@56458.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@56459.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@56460.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@56461.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@56462.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@56463.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@56464.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@56465.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@56466.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@56467.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@56468.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@56469.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@56470.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@56471.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@56472.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@56473.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@56474.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@56475.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@56476.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@56477.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@56478.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@56479.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@56480.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@56481.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@56482.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@56483.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@56484.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@56485.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@56486.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@56487.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@56488.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@56489.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@56490.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@56491.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@56492.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@56493.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@56494.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@56495.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@56496.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@56497.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@56498.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@56499.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@56500.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@56501.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@56502.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@56503.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@56504.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@56439.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@56420.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@56641.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@56634.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@56531.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@56530.4]
endmodule
module DRAMArbiter_1( // @[:@70870.2]
  input         clock, // @[:@70871.4]
  input         reset, // @[:@70872.4]
  input         io_enable, // @[:@70873.4]
  input         io_dram_cmd_ready, // @[:@70873.4]
  output        io_dram_cmd_valid, // @[:@70873.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@70873.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@70873.4]
  output        io_dram_cmd_bits_isWr, // @[:@70873.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@70873.4]
  input         io_dram_wdata_ready, // @[:@70873.4]
  output        io_dram_wdata_valid, // @[:@70873.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@70873.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@70873.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@70873.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@70873.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@70873.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@70873.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@70873.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@70873.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@70873.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@70873.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@70873.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@70873.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@70873.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@70873.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@70873.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@70873.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@70873.4]
  output        io_dram_wdata_bits_wlast, // @[:@70873.4]
  output        io_dram_rresp_ready, // @[:@70873.4]
  output        io_dram_wresp_ready, // @[:@70873.4]
  input         io_dram_wresp_valid, // @[:@70873.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@70873.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@71759.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@71773.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@72001.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@72116.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@72116.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@71759.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@71773.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@72001.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@72116.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@72341.4 DRAMArbiter.scala 100:23:@72344.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@72340.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@72339.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@72337.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@72336.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@72334.4 DRAMArbiter.scala 101:25:@72346.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@72318.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@72319.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@72320.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@72321.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@72322.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@72323.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@72324.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@72325.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@72326.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@72327.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@72328.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@72329.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@72330.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@72331.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@72332.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@72333.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@72254.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@72255.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@72256.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@72257.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@72258.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@72259.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@72260.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@72261.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@72262.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@72263.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@72264.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@72265.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@72266.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@72267.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@72268.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@72269.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@72270.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@72271.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@72272.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@72273.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@72274.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@72275.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@72276.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@72277.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@72278.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@72279.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@72280.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@72281.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@72282.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@72283.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@72284.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@72285.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@72286.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@72287.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@72288.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@72289.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@72290.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@72291.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@72292.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@72293.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@72294.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@72295.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@72296.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@72297.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@72298.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@72299.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@72300.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@72301.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@72302.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@72303.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@72304.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@72305.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@72306.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@72307.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@72308.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@72309.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@72310.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@72311.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@72312.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@72313.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@72314.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@72315.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@72316.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@72317.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@72253.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@72252.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@72233.4]
  assign StreamControllerStore_clock = clock; // @[:@71760.4]
  assign StreamControllerStore_reset = reset; // @[:@71761.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@71888.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@71881.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@71778.4]
  assign StreamControllerStore_io_store_cmd_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@71771.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = 64'h0; // @[DRAMArbiter.scala 68:18:@71770.4]
  assign StreamControllerStore_io_store_cmd_bits_size = 32'h0; // @[DRAMArbiter.scala 68:18:@71769.4]
  assign StreamControllerStore_io_store_data_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@71767.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = 32'h0; // @[DRAMArbiter.scala 68:18:@71766.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = 1'h0; // @[DRAMArbiter.scala 68:18:@71765.4]
  assign StreamControllerStore_io_store_wresp_ready = 1'h0; // @[DRAMArbiter.scala 68:18:@71764.4]
  assign StreamArbiter_clock = clock; // @[:@71774.4]
  assign StreamArbiter_reset = reset; // @[:@71775.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@71999.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@71998.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@71997.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@71995.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@71994.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@71992.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@71976.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@71977.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@71978.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@71979.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@71980.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@71981.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@71982.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@71983.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@71984.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@71985.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@71986.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@71987.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@71988.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@71989.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@71990.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@71991.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@71912.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@71913.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@71914.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@71915.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@71916.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@71917.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@71918.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@71919.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@71920.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@71921.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@71922.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@71923.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@71924.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@71925.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@71926.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@71927.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@71928.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@71929.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@71930.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@71931.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@71932.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@71933.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@71934.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@71935.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@71936.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@71937.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@71938.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@71939.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@71940.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@71941.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@71942.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@71943.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@71944.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@71945.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@71946.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@71947.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@71948.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@71949.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@71950.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@71951.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@71952.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@71953.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@71954.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@71955.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@71956.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@71957.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@71958.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@71959.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@71960.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@71961.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@71962.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@71963.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@71964.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@71965.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@71966.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@71967.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@71968.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@71969.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@71970.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@71971.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@71972.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@71973.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@71974.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@71975.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@71910.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@71891.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@72115.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@72108.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@72005.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@72004.4]
  assign AXICmdSplit_clock = clock; // @[:@72002.4]
  assign AXICmdSplit_reset = reset; // @[:@72003.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@72114.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@72113.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@72112.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@72110.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@72109.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@72107.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@72091.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@72092.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@72093.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@72094.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@72095.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@72096.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@72097.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@72098.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@72099.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@72100.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@72101.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@72102.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@72103.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@72104.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@72105.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@72106.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@72027.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@72028.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@72029.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@72030.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@72031.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@72032.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@72033.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@72034.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@72035.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@72036.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@72037.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@72038.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@72039.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@72040.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@72041.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@72042.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@72043.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@72044.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@72045.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@72046.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@72047.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@72048.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@72049.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@72050.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@72051.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@72052.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@72053.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@72054.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@72055.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@72056.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@72057.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@72058.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@72059.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@72060.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@72061.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@72062.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@72063.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@72064.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@72065.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@72066.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@72067.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@72068.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@72069.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@72070.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@72071.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@72072.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@72073.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@72074.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@72075.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@72076.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@72077.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@72078.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@72079.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@72080.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@72081.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@72082.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@72083.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@72084.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@72085.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@72086.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@72087.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@72088.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@72089.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@72090.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@72025.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@72006.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@72230.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@72223.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@72120.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@72119.4]
  assign AXICmdIssue_clock = clock; // @[:@72117.4]
  assign AXICmdIssue_reset = reset; // @[:@72118.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@72229.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@72228.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@72227.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@72225.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@72224.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@72222.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@72206.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@72207.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@72208.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@72209.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@72210.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@72211.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@72212.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@72213.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@72214.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@72215.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@72216.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@72217.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@72218.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@72219.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@72220.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@72221.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@72142.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@72143.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@72144.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@72145.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@72146.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@72147.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@72148.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@72149.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@72150.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@72151.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@72152.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@72153.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@72154.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@72155.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@72156.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@72157.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@72158.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@72159.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@72160.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@72161.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@72162.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@72163.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@72164.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@72165.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@72166.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@72167.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@72168.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@72169.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@72170.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@72171.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@72172.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@72173.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@72174.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@72175.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@72176.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@72177.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@72178.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@72179.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@72180.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@72181.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@72182.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@72183.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@72184.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@72185.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@72186.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@72187.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@72188.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@72189.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@72190.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@72191.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@72192.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@72193.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@72194.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@72195.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@72196.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@72197.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@72198.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@72199.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@72200.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@72201.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@72202.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@72203.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@72204.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@72205.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@72140.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@72121.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@72342.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@72335.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@72232.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@72231.4]
endmodule
module DRAMHeap( // @[:@102978.2]
  input         io_accel_0_req_valid, // @[:@102981.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@102981.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@102981.4]
  output        io_accel_0_resp_valid, // @[:@102981.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@102981.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@102981.4]
  output        io_host_0_req_valid, // @[:@102981.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@102981.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@102981.4]
  input         io_host_0_resp_valid, // @[:@102981.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@102981.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@102981.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@102988.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@102990.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@102989.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@102985.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@102984.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@102983.4]
endmodule
module FringeFF( // @[:@103024.2]
  input         clock, // @[:@103025.4]
  input         reset, // @[:@103026.4]
  input  [63:0] io_in, // @[:@103027.4]
  input         io_reset, // @[:@103027.4]
  output [63:0] io_out, // @[:@103027.4]
  input         io_enable // @[:@103027.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@103030.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@103030.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@103030.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@103030.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@103030.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@103035.4 package.scala 96:25:@103036.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@103041.6]
  RetimeWrapper_50 RetimeWrapper ( // @[package.scala 93:22:@103030.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@103035.4 package.scala 96:25:@103036.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@103041.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@103047.4]
  assign RetimeWrapper_clock = clock; // @[:@103031.4]
  assign RetimeWrapper_reset = reset; // @[:@103032.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@103034.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@103033.4]
endmodule
module MuxN( // @[:@131663.2]
  input  [63:0] io_ins_0, // @[:@131666.4]
  input  [63:0] io_ins_1, // @[:@131666.4]
  input  [63:0] io_ins_2, // @[:@131666.4]
  input  [63:0] io_ins_3, // @[:@131666.4]
  input  [63:0] io_ins_4, // @[:@131666.4]
  input  [63:0] io_ins_5, // @[:@131666.4]
  input  [63:0] io_ins_6, // @[:@131666.4]
  input  [63:0] io_ins_7, // @[:@131666.4]
  input  [63:0] io_ins_8, // @[:@131666.4]
  input  [63:0] io_ins_9, // @[:@131666.4]
  input  [63:0] io_ins_10, // @[:@131666.4]
  input  [63:0] io_ins_11, // @[:@131666.4]
  input  [63:0] io_ins_12, // @[:@131666.4]
  input  [63:0] io_ins_13, // @[:@131666.4]
  input  [63:0] io_ins_14, // @[:@131666.4]
  input  [63:0] io_ins_15, // @[:@131666.4]
  input  [63:0] io_ins_16, // @[:@131666.4]
  input  [63:0] io_ins_17, // @[:@131666.4]
  input  [63:0] io_ins_18, // @[:@131666.4]
  input  [63:0] io_ins_19, // @[:@131666.4]
  input  [63:0] io_ins_20, // @[:@131666.4]
  input  [63:0] io_ins_21, // @[:@131666.4]
  input  [63:0] io_ins_22, // @[:@131666.4]
  input  [63:0] io_ins_23, // @[:@131666.4]
  input  [63:0] io_ins_24, // @[:@131666.4]
  input  [63:0] io_ins_25, // @[:@131666.4]
  input  [63:0] io_ins_26, // @[:@131666.4]
  input  [63:0] io_ins_27, // @[:@131666.4]
  input  [63:0] io_ins_28, // @[:@131666.4]
  input  [63:0] io_ins_29, // @[:@131666.4]
  input  [63:0] io_ins_30, // @[:@131666.4]
  input  [63:0] io_ins_31, // @[:@131666.4]
  input  [63:0] io_ins_32, // @[:@131666.4]
  input  [63:0] io_ins_33, // @[:@131666.4]
  input  [63:0] io_ins_34, // @[:@131666.4]
  input  [63:0] io_ins_35, // @[:@131666.4]
  input  [63:0] io_ins_36, // @[:@131666.4]
  input  [63:0] io_ins_37, // @[:@131666.4]
  input  [63:0] io_ins_38, // @[:@131666.4]
  input  [63:0] io_ins_39, // @[:@131666.4]
  input  [63:0] io_ins_40, // @[:@131666.4]
  input  [63:0] io_ins_41, // @[:@131666.4]
  input  [63:0] io_ins_42, // @[:@131666.4]
  input  [63:0] io_ins_43, // @[:@131666.4]
  input  [63:0] io_ins_44, // @[:@131666.4]
  input  [63:0] io_ins_45, // @[:@131666.4]
  input  [63:0] io_ins_46, // @[:@131666.4]
  input  [63:0] io_ins_47, // @[:@131666.4]
  input  [63:0] io_ins_48, // @[:@131666.4]
  input  [63:0] io_ins_49, // @[:@131666.4]
  input  [63:0] io_ins_50, // @[:@131666.4]
  input  [63:0] io_ins_51, // @[:@131666.4]
  input  [63:0] io_ins_52, // @[:@131666.4]
  input  [63:0] io_ins_53, // @[:@131666.4]
  input  [63:0] io_ins_54, // @[:@131666.4]
  input  [63:0] io_ins_55, // @[:@131666.4]
  input  [63:0] io_ins_56, // @[:@131666.4]
  input  [63:0] io_ins_57, // @[:@131666.4]
  input  [63:0] io_ins_58, // @[:@131666.4]
  input  [63:0] io_ins_59, // @[:@131666.4]
  input  [63:0] io_ins_60, // @[:@131666.4]
  input  [63:0] io_ins_61, // @[:@131666.4]
  input  [63:0] io_ins_62, // @[:@131666.4]
  input  [63:0] io_ins_63, // @[:@131666.4]
  input  [63:0] io_ins_64, // @[:@131666.4]
  input  [63:0] io_ins_65, // @[:@131666.4]
  input  [63:0] io_ins_66, // @[:@131666.4]
  input  [63:0] io_ins_67, // @[:@131666.4]
  input  [63:0] io_ins_68, // @[:@131666.4]
  input  [63:0] io_ins_69, // @[:@131666.4]
  input  [63:0] io_ins_70, // @[:@131666.4]
  input  [63:0] io_ins_71, // @[:@131666.4]
  input  [63:0] io_ins_72, // @[:@131666.4]
  input  [63:0] io_ins_73, // @[:@131666.4]
  input  [63:0] io_ins_74, // @[:@131666.4]
  input  [63:0] io_ins_75, // @[:@131666.4]
  input  [63:0] io_ins_76, // @[:@131666.4]
  input  [63:0] io_ins_77, // @[:@131666.4]
  input  [63:0] io_ins_78, // @[:@131666.4]
  input  [63:0] io_ins_79, // @[:@131666.4]
  input  [63:0] io_ins_80, // @[:@131666.4]
  input  [63:0] io_ins_81, // @[:@131666.4]
  input  [63:0] io_ins_82, // @[:@131666.4]
  input  [63:0] io_ins_83, // @[:@131666.4]
  input  [63:0] io_ins_84, // @[:@131666.4]
  input  [63:0] io_ins_85, // @[:@131666.4]
  input  [63:0] io_ins_86, // @[:@131666.4]
  input  [63:0] io_ins_87, // @[:@131666.4]
  input  [63:0] io_ins_88, // @[:@131666.4]
  input  [63:0] io_ins_89, // @[:@131666.4]
  input  [63:0] io_ins_90, // @[:@131666.4]
  input  [63:0] io_ins_91, // @[:@131666.4]
  input  [63:0] io_ins_92, // @[:@131666.4]
  input  [63:0] io_ins_93, // @[:@131666.4]
  input  [63:0] io_ins_94, // @[:@131666.4]
  input  [63:0] io_ins_95, // @[:@131666.4]
  input  [63:0] io_ins_96, // @[:@131666.4]
  input  [63:0] io_ins_97, // @[:@131666.4]
  input  [63:0] io_ins_98, // @[:@131666.4]
  input  [63:0] io_ins_99, // @[:@131666.4]
  input  [63:0] io_ins_100, // @[:@131666.4]
  input  [63:0] io_ins_101, // @[:@131666.4]
  input  [63:0] io_ins_102, // @[:@131666.4]
  input  [63:0] io_ins_103, // @[:@131666.4]
  input  [63:0] io_ins_104, // @[:@131666.4]
  input  [63:0] io_ins_105, // @[:@131666.4]
  input  [63:0] io_ins_106, // @[:@131666.4]
  input  [63:0] io_ins_107, // @[:@131666.4]
  input  [63:0] io_ins_108, // @[:@131666.4]
  input  [63:0] io_ins_109, // @[:@131666.4]
  input  [63:0] io_ins_110, // @[:@131666.4]
  input  [63:0] io_ins_111, // @[:@131666.4]
  input  [63:0] io_ins_112, // @[:@131666.4]
  input  [63:0] io_ins_113, // @[:@131666.4]
  input  [63:0] io_ins_114, // @[:@131666.4]
  input  [63:0] io_ins_115, // @[:@131666.4]
  input  [63:0] io_ins_116, // @[:@131666.4]
  input  [63:0] io_ins_117, // @[:@131666.4]
  input  [63:0] io_ins_118, // @[:@131666.4]
  input  [63:0] io_ins_119, // @[:@131666.4]
  input  [63:0] io_ins_120, // @[:@131666.4]
  input  [63:0] io_ins_121, // @[:@131666.4]
  input  [63:0] io_ins_122, // @[:@131666.4]
  input  [63:0] io_ins_123, // @[:@131666.4]
  input  [63:0] io_ins_124, // @[:@131666.4]
  input  [63:0] io_ins_125, // @[:@131666.4]
  input  [63:0] io_ins_126, // @[:@131666.4]
  input  [63:0] io_ins_127, // @[:@131666.4]
  input  [63:0] io_ins_128, // @[:@131666.4]
  input  [63:0] io_ins_129, // @[:@131666.4]
  input  [63:0] io_ins_130, // @[:@131666.4]
  input  [63:0] io_ins_131, // @[:@131666.4]
  input  [63:0] io_ins_132, // @[:@131666.4]
  input  [63:0] io_ins_133, // @[:@131666.4]
  input  [63:0] io_ins_134, // @[:@131666.4]
  input  [63:0] io_ins_135, // @[:@131666.4]
  input  [63:0] io_ins_136, // @[:@131666.4]
  input  [63:0] io_ins_137, // @[:@131666.4]
  input  [63:0] io_ins_138, // @[:@131666.4]
  input  [63:0] io_ins_139, // @[:@131666.4]
  input  [63:0] io_ins_140, // @[:@131666.4]
  input  [63:0] io_ins_141, // @[:@131666.4]
  input  [63:0] io_ins_142, // @[:@131666.4]
  input  [63:0] io_ins_143, // @[:@131666.4]
  input  [63:0] io_ins_144, // @[:@131666.4]
  input  [63:0] io_ins_145, // @[:@131666.4]
  input  [63:0] io_ins_146, // @[:@131666.4]
  input  [63:0] io_ins_147, // @[:@131666.4]
  input  [63:0] io_ins_148, // @[:@131666.4]
  input  [63:0] io_ins_149, // @[:@131666.4]
  input  [63:0] io_ins_150, // @[:@131666.4]
  input  [63:0] io_ins_151, // @[:@131666.4]
  input  [63:0] io_ins_152, // @[:@131666.4]
  input  [63:0] io_ins_153, // @[:@131666.4]
  input  [63:0] io_ins_154, // @[:@131666.4]
  input  [63:0] io_ins_155, // @[:@131666.4]
  input  [63:0] io_ins_156, // @[:@131666.4]
  input  [63:0] io_ins_157, // @[:@131666.4]
  input  [63:0] io_ins_158, // @[:@131666.4]
  input  [63:0] io_ins_159, // @[:@131666.4]
  input  [63:0] io_ins_160, // @[:@131666.4]
  input  [63:0] io_ins_161, // @[:@131666.4]
  input  [63:0] io_ins_162, // @[:@131666.4]
  input  [63:0] io_ins_163, // @[:@131666.4]
  input  [63:0] io_ins_164, // @[:@131666.4]
  input  [63:0] io_ins_165, // @[:@131666.4]
  input  [63:0] io_ins_166, // @[:@131666.4]
  input  [63:0] io_ins_167, // @[:@131666.4]
  input  [63:0] io_ins_168, // @[:@131666.4]
  input  [63:0] io_ins_169, // @[:@131666.4]
  input  [63:0] io_ins_170, // @[:@131666.4]
  input  [63:0] io_ins_171, // @[:@131666.4]
  input  [63:0] io_ins_172, // @[:@131666.4]
  input  [63:0] io_ins_173, // @[:@131666.4]
  input  [63:0] io_ins_174, // @[:@131666.4]
  input  [63:0] io_ins_175, // @[:@131666.4]
  input  [63:0] io_ins_176, // @[:@131666.4]
  input  [63:0] io_ins_177, // @[:@131666.4]
  input  [63:0] io_ins_178, // @[:@131666.4]
  input  [63:0] io_ins_179, // @[:@131666.4]
  input  [63:0] io_ins_180, // @[:@131666.4]
  input  [63:0] io_ins_181, // @[:@131666.4]
  input  [63:0] io_ins_182, // @[:@131666.4]
  input  [63:0] io_ins_183, // @[:@131666.4]
  input  [63:0] io_ins_184, // @[:@131666.4]
  input  [63:0] io_ins_185, // @[:@131666.4]
  input  [63:0] io_ins_186, // @[:@131666.4]
  input  [63:0] io_ins_187, // @[:@131666.4]
  input  [63:0] io_ins_188, // @[:@131666.4]
  input  [63:0] io_ins_189, // @[:@131666.4]
  input  [63:0] io_ins_190, // @[:@131666.4]
  input  [63:0] io_ins_191, // @[:@131666.4]
  input  [63:0] io_ins_192, // @[:@131666.4]
  input  [63:0] io_ins_193, // @[:@131666.4]
  input  [63:0] io_ins_194, // @[:@131666.4]
  input  [63:0] io_ins_195, // @[:@131666.4]
  input  [63:0] io_ins_196, // @[:@131666.4]
  input  [63:0] io_ins_197, // @[:@131666.4]
  input  [63:0] io_ins_198, // @[:@131666.4]
  input  [63:0] io_ins_199, // @[:@131666.4]
  input  [63:0] io_ins_200, // @[:@131666.4]
  input  [63:0] io_ins_201, // @[:@131666.4]
  input  [63:0] io_ins_202, // @[:@131666.4]
  input  [63:0] io_ins_203, // @[:@131666.4]
  input  [63:0] io_ins_204, // @[:@131666.4]
  input  [63:0] io_ins_205, // @[:@131666.4]
  input  [63:0] io_ins_206, // @[:@131666.4]
  input  [63:0] io_ins_207, // @[:@131666.4]
  input  [63:0] io_ins_208, // @[:@131666.4]
  input  [63:0] io_ins_209, // @[:@131666.4]
  input  [63:0] io_ins_210, // @[:@131666.4]
  input  [63:0] io_ins_211, // @[:@131666.4]
  input  [63:0] io_ins_212, // @[:@131666.4]
  input  [63:0] io_ins_213, // @[:@131666.4]
  input  [63:0] io_ins_214, // @[:@131666.4]
  input  [63:0] io_ins_215, // @[:@131666.4]
  input  [63:0] io_ins_216, // @[:@131666.4]
  input  [63:0] io_ins_217, // @[:@131666.4]
  input  [63:0] io_ins_218, // @[:@131666.4]
  input  [63:0] io_ins_219, // @[:@131666.4]
  input  [63:0] io_ins_220, // @[:@131666.4]
  input  [63:0] io_ins_221, // @[:@131666.4]
  input  [63:0] io_ins_222, // @[:@131666.4]
  input  [63:0] io_ins_223, // @[:@131666.4]
  input  [63:0] io_ins_224, // @[:@131666.4]
  input  [63:0] io_ins_225, // @[:@131666.4]
  input  [63:0] io_ins_226, // @[:@131666.4]
  input  [63:0] io_ins_227, // @[:@131666.4]
  input  [63:0] io_ins_228, // @[:@131666.4]
  input  [63:0] io_ins_229, // @[:@131666.4]
  input  [63:0] io_ins_230, // @[:@131666.4]
  input  [63:0] io_ins_231, // @[:@131666.4]
  input  [63:0] io_ins_232, // @[:@131666.4]
  input  [63:0] io_ins_233, // @[:@131666.4]
  input  [63:0] io_ins_234, // @[:@131666.4]
  input  [63:0] io_ins_235, // @[:@131666.4]
  input  [63:0] io_ins_236, // @[:@131666.4]
  input  [63:0] io_ins_237, // @[:@131666.4]
  input  [63:0] io_ins_238, // @[:@131666.4]
  input  [63:0] io_ins_239, // @[:@131666.4]
  input  [63:0] io_ins_240, // @[:@131666.4]
  input  [63:0] io_ins_241, // @[:@131666.4]
  input  [63:0] io_ins_242, // @[:@131666.4]
  input  [63:0] io_ins_243, // @[:@131666.4]
  input  [63:0] io_ins_244, // @[:@131666.4]
  input  [63:0] io_ins_245, // @[:@131666.4]
  input  [63:0] io_ins_246, // @[:@131666.4]
  input  [63:0] io_ins_247, // @[:@131666.4]
  input  [63:0] io_ins_248, // @[:@131666.4]
  input  [63:0] io_ins_249, // @[:@131666.4]
  input  [63:0] io_ins_250, // @[:@131666.4]
  input  [63:0] io_ins_251, // @[:@131666.4]
  input  [63:0] io_ins_252, // @[:@131666.4]
  input  [63:0] io_ins_253, // @[:@131666.4]
  input  [63:0] io_ins_254, // @[:@131666.4]
  input  [63:0] io_ins_255, // @[:@131666.4]
  input  [63:0] io_ins_256, // @[:@131666.4]
  input  [63:0] io_ins_257, // @[:@131666.4]
  input  [63:0] io_ins_258, // @[:@131666.4]
  input  [63:0] io_ins_259, // @[:@131666.4]
  input  [63:0] io_ins_260, // @[:@131666.4]
  input  [63:0] io_ins_261, // @[:@131666.4]
  input  [63:0] io_ins_262, // @[:@131666.4]
  input  [63:0] io_ins_263, // @[:@131666.4]
  input  [63:0] io_ins_264, // @[:@131666.4]
  input  [63:0] io_ins_265, // @[:@131666.4]
  input  [63:0] io_ins_266, // @[:@131666.4]
  input  [63:0] io_ins_267, // @[:@131666.4]
  input  [63:0] io_ins_268, // @[:@131666.4]
  input  [63:0] io_ins_269, // @[:@131666.4]
  input  [63:0] io_ins_270, // @[:@131666.4]
  input  [63:0] io_ins_271, // @[:@131666.4]
  input  [63:0] io_ins_272, // @[:@131666.4]
  input  [63:0] io_ins_273, // @[:@131666.4]
  input  [63:0] io_ins_274, // @[:@131666.4]
  input  [63:0] io_ins_275, // @[:@131666.4]
  input  [63:0] io_ins_276, // @[:@131666.4]
  input  [63:0] io_ins_277, // @[:@131666.4]
  input  [63:0] io_ins_278, // @[:@131666.4]
  input  [63:0] io_ins_279, // @[:@131666.4]
  input  [63:0] io_ins_280, // @[:@131666.4]
  input  [63:0] io_ins_281, // @[:@131666.4]
  input  [63:0] io_ins_282, // @[:@131666.4]
  input  [63:0] io_ins_283, // @[:@131666.4]
  input  [63:0] io_ins_284, // @[:@131666.4]
  input  [63:0] io_ins_285, // @[:@131666.4]
  input  [63:0] io_ins_286, // @[:@131666.4]
  input  [63:0] io_ins_287, // @[:@131666.4]
  input  [63:0] io_ins_288, // @[:@131666.4]
  input  [63:0] io_ins_289, // @[:@131666.4]
  input  [63:0] io_ins_290, // @[:@131666.4]
  input  [63:0] io_ins_291, // @[:@131666.4]
  input  [63:0] io_ins_292, // @[:@131666.4]
  input  [63:0] io_ins_293, // @[:@131666.4]
  input  [63:0] io_ins_294, // @[:@131666.4]
  input  [63:0] io_ins_295, // @[:@131666.4]
  input  [63:0] io_ins_296, // @[:@131666.4]
  input  [63:0] io_ins_297, // @[:@131666.4]
  input  [63:0] io_ins_298, // @[:@131666.4]
  input  [63:0] io_ins_299, // @[:@131666.4]
  input  [63:0] io_ins_300, // @[:@131666.4]
  input  [63:0] io_ins_301, // @[:@131666.4]
  input  [63:0] io_ins_302, // @[:@131666.4]
  input  [63:0] io_ins_303, // @[:@131666.4]
  input  [63:0] io_ins_304, // @[:@131666.4]
  input  [63:0] io_ins_305, // @[:@131666.4]
  input  [63:0] io_ins_306, // @[:@131666.4]
  input  [63:0] io_ins_307, // @[:@131666.4]
  input  [63:0] io_ins_308, // @[:@131666.4]
  input  [63:0] io_ins_309, // @[:@131666.4]
  input  [63:0] io_ins_310, // @[:@131666.4]
  input  [63:0] io_ins_311, // @[:@131666.4]
  input  [63:0] io_ins_312, // @[:@131666.4]
  input  [63:0] io_ins_313, // @[:@131666.4]
  input  [63:0] io_ins_314, // @[:@131666.4]
  input  [63:0] io_ins_315, // @[:@131666.4]
  input  [63:0] io_ins_316, // @[:@131666.4]
  input  [63:0] io_ins_317, // @[:@131666.4]
  input  [63:0] io_ins_318, // @[:@131666.4]
  input  [63:0] io_ins_319, // @[:@131666.4]
  input  [63:0] io_ins_320, // @[:@131666.4]
  input  [63:0] io_ins_321, // @[:@131666.4]
  input  [63:0] io_ins_322, // @[:@131666.4]
  input  [63:0] io_ins_323, // @[:@131666.4]
  input  [63:0] io_ins_324, // @[:@131666.4]
  input  [63:0] io_ins_325, // @[:@131666.4]
  input  [63:0] io_ins_326, // @[:@131666.4]
  input  [63:0] io_ins_327, // @[:@131666.4]
  input  [63:0] io_ins_328, // @[:@131666.4]
  input  [63:0] io_ins_329, // @[:@131666.4]
  input  [63:0] io_ins_330, // @[:@131666.4]
  input  [63:0] io_ins_331, // @[:@131666.4]
  input  [63:0] io_ins_332, // @[:@131666.4]
  input  [63:0] io_ins_333, // @[:@131666.4]
  input  [63:0] io_ins_334, // @[:@131666.4]
  input  [63:0] io_ins_335, // @[:@131666.4]
  input  [63:0] io_ins_336, // @[:@131666.4]
  input  [63:0] io_ins_337, // @[:@131666.4]
  input  [63:0] io_ins_338, // @[:@131666.4]
  input  [63:0] io_ins_339, // @[:@131666.4]
  input  [63:0] io_ins_340, // @[:@131666.4]
  input  [63:0] io_ins_341, // @[:@131666.4]
  input  [63:0] io_ins_342, // @[:@131666.4]
  input  [63:0] io_ins_343, // @[:@131666.4]
  input  [63:0] io_ins_344, // @[:@131666.4]
  input  [63:0] io_ins_345, // @[:@131666.4]
  input  [63:0] io_ins_346, // @[:@131666.4]
  input  [63:0] io_ins_347, // @[:@131666.4]
  input  [63:0] io_ins_348, // @[:@131666.4]
  input  [63:0] io_ins_349, // @[:@131666.4]
  input  [63:0] io_ins_350, // @[:@131666.4]
  input  [63:0] io_ins_351, // @[:@131666.4]
  input  [63:0] io_ins_352, // @[:@131666.4]
  input  [63:0] io_ins_353, // @[:@131666.4]
  input  [63:0] io_ins_354, // @[:@131666.4]
  input  [63:0] io_ins_355, // @[:@131666.4]
  input  [63:0] io_ins_356, // @[:@131666.4]
  input  [63:0] io_ins_357, // @[:@131666.4]
  input  [63:0] io_ins_358, // @[:@131666.4]
  input  [63:0] io_ins_359, // @[:@131666.4]
  input  [63:0] io_ins_360, // @[:@131666.4]
  input  [63:0] io_ins_361, // @[:@131666.4]
  input  [63:0] io_ins_362, // @[:@131666.4]
  input  [63:0] io_ins_363, // @[:@131666.4]
  input  [63:0] io_ins_364, // @[:@131666.4]
  input  [63:0] io_ins_365, // @[:@131666.4]
  input  [63:0] io_ins_366, // @[:@131666.4]
  input  [63:0] io_ins_367, // @[:@131666.4]
  input  [63:0] io_ins_368, // @[:@131666.4]
  input  [63:0] io_ins_369, // @[:@131666.4]
  input  [63:0] io_ins_370, // @[:@131666.4]
  input  [63:0] io_ins_371, // @[:@131666.4]
  input  [63:0] io_ins_372, // @[:@131666.4]
  input  [63:0] io_ins_373, // @[:@131666.4]
  input  [63:0] io_ins_374, // @[:@131666.4]
  input  [63:0] io_ins_375, // @[:@131666.4]
  input  [63:0] io_ins_376, // @[:@131666.4]
  input  [63:0] io_ins_377, // @[:@131666.4]
  input  [63:0] io_ins_378, // @[:@131666.4]
  input  [63:0] io_ins_379, // @[:@131666.4]
  input  [63:0] io_ins_380, // @[:@131666.4]
  input  [63:0] io_ins_381, // @[:@131666.4]
  input  [63:0] io_ins_382, // @[:@131666.4]
  input  [63:0] io_ins_383, // @[:@131666.4]
  input  [63:0] io_ins_384, // @[:@131666.4]
  input  [63:0] io_ins_385, // @[:@131666.4]
  input  [63:0] io_ins_386, // @[:@131666.4]
  input  [63:0] io_ins_387, // @[:@131666.4]
  input  [63:0] io_ins_388, // @[:@131666.4]
  input  [63:0] io_ins_389, // @[:@131666.4]
  input  [63:0] io_ins_390, // @[:@131666.4]
  input  [63:0] io_ins_391, // @[:@131666.4]
  input  [63:0] io_ins_392, // @[:@131666.4]
  input  [63:0] io_ins_393, // @[:@131666.4]
  input  [63:0] io_ins_394, // @[:@131666.4]
  input  [63:0] io_ins_395, // @[:@131666.4]
  input  [63:0] io_ins_396, // @[:@131666.4]
  input  [63:0] io_ins_397, // @[:@131666.4]
  input  [63:0] io_ins_398, // @[:@131666.4]
  input  [63:0] io_ins_399, // @[:@131666.4]
  input  [63:0] io_ins_400, // @[:@131666.4]
  input  [63:0] io_ins_401, // @[:@131666.4]
  input  [63:0] io_ins_402, // @[:@131666.4]
  input  [63:0] io_ins_403, // @[:@131666.4]
  input  [63:0] io_ins_404, // @[:@131666.4]
  input  [63:0] io_ins_405, // @[:@131666.4]
  input  [63:0] io_ins_406, // @[:@131666.4]
  input  [63:0] io_ins_407, // @[:@131666.4]
  input  [63:0] io_ins_408, // @[:@131666.4]
  input  [63:0] io_ins_409, // @[:@131666.4]
  input  [63:0] io_ins_410, // @[:@131666.4]
  input  [63:0] io_ins_411, // @[:@131666.4]
  input  [63:0] io_ins_412, // @[:@131666.4]
  input  [63:0] io_ins_413, // @[:@131666.4]
  input  [63:0] io_ins_414, // @[:@131666.4]
  input  [63:0] io_ins_415, // @[:@131666.4]
  input  [63:0] io_ins_416, // @[:@131666.4]
  input  [63:0] io_ins_417, // @[:@131666.4]
  input  [63:0] io_ins_418, // @[:@131666.4]
  input  [63:0] io_ins_419, // @[:@131666.4]
  input  [63:0] io_ins_420, // @[:@131666.4]
  input  [63:0] io_ins_421, // @[:@131666.4]
  input  [63:0] io_ins_422, // @[:@131666.4]
  input  [63:0] io_ins_423, // @[:@131666.4]
  input  [63:0] io_ins_424, // @[:@131666.4]
  input  [63:0] io_ins_425, // @[:@131666.4]
  input  [63:0] io_ins_426, // @[:@131666.4]
  input  [63:0] io_ins_427, // @[:@131666.4]
  input  [63:0] io_ins_428, // @[:@131666.4]
  input  [63:0] io_ins_429, // @[:@131666.4]
  input  [63:0] io_ins_430, // @[:@131666.4]
  input  [63:0] io_ins_431, // @[:@131666.4]
  input  [63:0] io_ins_432, // @[:@131666.4]
  input  [63:0] io_ins_433, // @[:@131666.4]
  input  [63:0] io_ins_434, // @[:@131666.4]
  input  [63:0] io_ins_435, // @[:@131666.4]
  input  [63:0] io_ins_436, // @[:@131666.4]
  input  [63:0] io_ins_437, // @[:@131666.4]
  input  [63:0] io_ins_438, // @[:@131666.4]
  input  [63:0] io_ins_439, // @[:@131666.4]
  input  [63:0] io_ins_440, // @[:@131666.4]
  input  [63:0] io_ins_441, // @[:@131666.4]
  input  [63:0] io_ins_442, // @[:@131666.4]
  input  [63:0] io_ins_443, // @[:@131666.4]
  input  [63:0] io_ins_444, // @[:@131666.4]
  input  [63:0] io_ins_445, // @[:@131666.4]
  input  [63:0] io_ins_446, // @[:@131666.4]
  input  [63:0] io_ins_447, // @[:@131666.4]
  input  [63:0] io_ins_448, // @[:@131666.4]
  input  [63:0] io_ins_449, // @[:@131666.4]
  input  [63:0] io_ins_450, // @[:@131666.4]
  input  [63:0] io_ins_451, // @[:@131666.4]
  input  [63:0] io_ins_452, // @[:@131666.4]
  input  [63:0] io_ins_453, // @[:@131666.4]
  input  [63:0] io_ins_454, // @[:@131666.4]
  input  [63:0] io_ins_455, // @[:@131666.4]
  input  [63:0] io_ins_456, // @[:@131666.4]
  input  [63:0] io_ins_457, // @[:@131666.4]
  input  [63:0] io_ins_458, // @[:@131666.4]
  input  [63:0] io_ins_459, // @[:@131666.4]
  input  [63:0] io_ins_460, // @[:@131666.4]
  input  [63:0] io_ins_461, // @[:@131666.4]
  input  [63:0] io_ins_462, // @[:@131666.4]
  input  [63:0] io_ins_463, // @[:@131666.4]
  input  [63:0] io_ins_464, // @[:@131666.4]
  input  [63:0] io_ins_465, // @[:@131666.4]
  input  [63:0] io_ins_466, // @[:@131666.4]
  input  [63:0] io_ins_467, // @[:@131666.4]
  input  [63:0] io_ins_468, // @[:@131666.4]
  input  [63:0] io_ins_469, // @[:@131666.4]
  input  [63:0] io_ins_470, // @[:@131666.4]
  input  [63:0] io_ins_471, // @[:@131666.4]
  input  [63:0] io_ins_472, // @[:@131666.4]
  input  [63:0] io_ins_473, // @[:@131666.4]
  input  [63:0] io_ins_474, // @[:@131666.4]
  input  [63:0] io_ins_475, // @[:@131666.4]
  input  [63:0] io_ins_476, // @[:@131666.4]
  input  [63:0] io_ins_477, // @[:@131666.4]
  input  [63:0] io_ins_478, // @[:@131666.4]
  input  [63:0] io_ins_479, // @[:@131666.4]
  input  [63:0] io_ins_480, // @[:@131666.4]
  input  [63:0] io_ins_481, // @[:@131666.4]
  input  [63:0] io_ins_482, // @[:@131666.4]
  input  [63:0] io_ins_483, // @[:@131666.4]
  input  [63:0] io_ins_484, // @[:@131666.4]
  input  [63:0] io_ins_485, // @[:@131666.4]
  input  [63:0] io_ins_486, // @[:@131666.4]
  input  [63:0] io_ins_487, // @[:@131666.4]
  input  [63:0] io_ins_488, // @[:@131666.4]
  input  [63:0] io_ins_489, // @[:@131666.4]
  input  [63:0] io_ins_490, // @[:@131666.4]
  input  [63:0] io_ins_491, // @[:@131666.4]
  input  [63:0] io_ins_492, // @[:@131666.4]
  input  [63:0] io_ins_493, // @[:@131666.4]
  input  [63:0] io_ins_494, // @[:@131666.4]
  input  [63:0] io_ins_495, // @[:@131666.4]
  input  [63:0] io_ins_496, // @[:@131666.4]
  input  [63:0] io_ins_497, // @[:@131666.4]
  input  [63:0] io_ins_498, // @[:@131666.4]
  input  [63:0] io_ins_499, // @[:@131666.4]
  input  [63:0] io_ins_500, // @[:@131666.4]
  input  [63:0] io_ins_501, // @[:@131666.4]
  input  [63:0] io_ins_502, // @[:@131666.4]
  input  [8:0]  io_sel, // @[:@131666.4]
  output [63:0] io_out // @[:@131666.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@131668.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_1 = 9'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_2 = 9'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_3 = 9'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_4 = 9'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_5 = 9'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_6 = 9'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_7 = 9'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_8 = 9'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_9 = 9'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_10 = 9'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_11 = 9'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_12 = 9'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_13 = 9'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_14 = 9'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_15 = 9'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_16 = 9'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_17 = 9'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_18 = 9'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_19 = 9'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_20 = 9'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_21 = 9'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_22 = 9'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_23 = 9'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_24 = 9'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_25 = 9'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_26 = 9'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_27 = 9'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_28 = 9'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_29 = 9'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_30 = 9'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_31 = 9'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_32 = 9'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_33 = 9'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_34 = 9'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_35 = 9'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_36 = 9'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_37 = 9'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_38 = 9'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_39 = 9'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_40 = 9'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_41 = 9'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_42 = 9'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_43 = 9'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_44 = 9'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_45 = 9'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_46 = 9'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_47 = 9'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_48 = 9'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_49 = 9'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_50 = 9'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_51 = 9'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_52 = 9'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_53 = 9'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_54 = 9'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_55 = 9'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_56 = 9'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_57 = 9'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_58 = 9'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_59 = 9'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_60 = 9'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_61 = 9'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_62 = 9'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_63 = 9'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_64 = 9'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_65 = 9'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_66 = 9'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_67 = 9'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_68 = 9'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_69 = 9'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_70 = 9'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_71 = 9'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_72 = 9'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_73 = 9'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_74 = 9'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_75 = 9'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_76 = 9'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_77 = 9'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_78 = 9'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_79 = 9'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_80 = 9'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_81 = 9'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_82 = 9'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_83 = 9'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_84 = 9'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_85 = 9'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_86 = 9'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_87 = 9'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_88 = 9'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_89 = 9'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_90 = 9'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_91 = 9'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_92 = 9'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_93 = 9'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_94 = 9'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_95 = 9'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_96 = 9'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_97 = 9'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_98 = 9'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_99 = 9'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_100 = 9'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_101 = 9'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_102 = 9'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_103 = 9'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_104 = 9'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_105 = 9'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_106 = 9'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_107 = 9'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_108 = 9'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_109 = 9'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_110 = 9'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_111 = 9'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_112 = 9'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_113 = 9'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_114 = 9'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_115 = 9'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_116 = 9'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_117 = 9'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_118 = 9'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_119 = 9'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_120 = 9'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_121 = 9'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_122 = 9'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_123 = 9'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_124 = 9'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_125 = 9'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_126 = 9'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_127 = 9'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_128 = 9'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_129 = 9'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_130 = 9'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_131 = 9'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_132 = 9'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_133 = 9'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_134 = 9'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_135 = 9'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_136 = 9'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_137 = 9'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_138 = 9'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_139 = 9'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_140 = 9'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_141 = 9'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_142 = 9'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_143 = 9'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_144 = 9'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_145 = 9'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_146 = 9'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_147 = 9'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_148 = 9'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_149 = 9'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_150 = 9'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_151 = 9'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_152 = 9'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_153 = 9'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_154 = 9'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_155 = 9'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_156 = 9'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_157 = 9'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_158 = 9'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_159 = 9'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_160 = 9'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_161 = 9'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_162 = 9'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_163 = 9'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_164 = 9'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_165 = 9'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_166 = 9'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_167 = 9'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_168 = 9'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_169 = 9'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_170 = 9'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_171 = 9'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_172 = 9'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_173 = 9'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_174 = 9'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_175 = 9'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_176 = 9'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_177 = 9'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_178 = 9'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_179 = 9'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_180 = 9'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_181 = 9'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_182 = 9'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_183 = 9'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_184 = 9'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_185 = 9'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_186 = 9'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_187 = 9'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_188 = 9'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_189 = 9'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_190 = 9'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_191 = 9'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_192 = 9'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_193 = 9'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_194 = 9'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_195 = 9'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_196 = 9'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_197 = 9'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_198 = 9'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_199 = 9'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_200 = 9'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_201 = 9'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_202 = 9'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_203 = 9'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_204 = 9'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_205 = 9'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_206 = 9'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_207 = 9'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_208 = 9'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_209 = 9'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_210 = 9'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_211 = 9'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_212 = 9'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_213 = 9'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_214 = 9'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_215 = 9'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_216 = 9'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_217 = 9'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_218 = 9'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_219 = 9'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_220 = 9'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_221 = 9'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_222 = 9'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_223 = 9'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_224 = 9'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_225 = 9'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_226 = 9'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_227 = 9'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_228 = 9'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_229 = 9'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_230 = 9'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_231 = 9'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_232 = 9'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_233 = 9'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_234 = 9'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_235 = 9'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_236 = 9'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_237 = 9'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_238 = 9'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_239 = 9'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_240 = 9'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_241 = 9'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_242 = 9'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_243 = 9'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_244 = 9'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_245 = 9'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_246 = 9'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_247 = 9'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_248 = 9'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_249 = 9'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_250 = 9'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_251 = 9'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_252 = 9'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_253 = 9'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_254 = 9'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_255 = 9'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_256 = 9'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_257 = 9'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_258 = 9'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_259 = 9'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_260 = 9'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_261 = 9'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_262 = 9'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_263 = 9'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_264 = 9'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_265 = 9'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_266 = 9'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_267 = 9'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_268 = 9'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_269 = 9'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_270 = 9'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_271 = 9'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_272 = 9'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_273 = 9'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_274 = 9'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_275 = 9'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_276 = 9'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_277 = 9'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_278 = 9'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_279 = 9'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_280 = 9'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_281 = 9'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_282 = 9'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_283 = 9'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_284 = 9'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_285 = 9'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_286 = 9'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_287 = 9'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_288 = 9'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_289 = 9'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_290 = 9'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_291 = 9'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_292 = 9'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_293 = 9'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_294 = 9'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_295 = 9'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_296 = 9'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_297 = 9'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_298 = 9'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_299 = 9'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_300 = 9'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_301 = 9'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_302 = 9'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_303 = 9'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_304 = 9'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_305 = 9'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_306 = 9'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_307 = 9'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_308 = 9'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_309 = 9'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_310 = 9'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_311 = 9'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_312 = 9'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_313 = 9'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_314 = 9'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_315 = 9'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_316 = 9'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_317 = 9'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_318 = 9'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_319 = 9'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_320 = 9'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_321 = 9'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_322 = 9'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_323 = 9'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_324 = 9'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_325 = 9'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_326 = 9'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_327 = 9'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_328 = 9'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_329 = 9'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_330 = 9'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_331 = 9'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_332 = 9'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_333 = 9'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_334 = 9'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_335 = 9'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_336 = 9'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_337 = 9'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_338 = 9'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_339 = 9'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_340 = 9'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_341 = 9'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_342 = 9'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_343 = 9'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_344 = 9'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_345 = 9'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_346 = 9'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_347 = 9'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_348 = 9'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_349 = 9'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_350 = 9'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_351 = 9'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_352 = 9'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_353 = 9'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_354 = 9'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_355 = 9'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_356 = 9'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_357 = 9'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_358 = 9'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_359 = 9'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_360 = 9'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_361 = 9'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_362 = 9'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_363 = 9'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_364 = 9'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_365 = 9'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_366 = 9'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_367 = 9'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_368 = 9'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_369 = 9'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_370 = 9'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_371 = 9'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_372 = 9'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_373 = 9'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_374 = 9'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_375 = 9'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_376 = 9'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_377 = 9'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_378 = 9'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_379 = 9'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_380 = 9'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_381 = 9'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_382 = 9'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_383 = 9'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_384 = 9'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_385 = 9'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_386 = 9'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_387 = 9'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_388 = 9'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_389 = 9'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_390 = 9'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_391 = 9'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_392 = 9'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_393 = 9'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_394 = 9'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_395 = 9'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_396 = 9'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_397 = 9'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_398 = 9'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_399 = 9'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_400 = 9'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_401 = 9'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_402 = 9'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_403 = 9'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_404 = 9'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_405 = 9'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_406 = 9'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_407 = 9'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_408 = 9'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_409 = 9'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_410 = 9'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_411 = 9'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_412 = 9'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_413 = 9'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_414 = 9'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_415 = 9'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_416 = 9'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_417 = 9'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_418 = 9'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_419 = 9'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_420 = 9'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_421 = 9'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_422 = 9'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_423 = 9'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_424 = 9'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_425 = 9'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_426 = 9'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_427 = 9'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_428 = 9'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_429 = 9'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_430 = 9'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_431 = 9'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_432 = 9'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_433 = 9'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_434 = 9'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_435 = 9'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_436 = 9'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_437 = 9'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_438 = 9'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_439 = 9'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_440 = 9'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_441 = 9'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_442 = 9'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_443 = 9'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_444 = 9'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_445 = 9'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_446 = 9'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_447 = 9'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_448 = 9'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_449 = 9'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_450 = 9'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_451 = 9'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_452 = 9'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_453 = 9'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_454 = 9'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_455 = 9'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_456 = 9'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_457 = 9'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_458 = 9'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_459 = 9'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_460 = 9'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_461 = 9'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_462 = 9'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_463 = 9'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_464 = 9'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_465 = 9'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_466 = 9'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_467 = 9'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_468 = 9'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_469 = 9'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_470 = 9'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_471 = 9'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_472 = 9'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_473 = 9'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_474 = 9'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_475 = 9'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_476 = 9'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_477 = 9'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_478 = 9'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_479 = 9'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_480 = 9'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_481 = 9'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_482 = 9'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_483 = 9'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_484 = 9'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_485 = 9'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_486 = 9'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_487 = 9'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_488 = 9'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_489 = 9'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_490 = 9'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_491 = 9'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_492 = 9'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_493 = 9'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_494 = 9'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_495 = 9'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_496 = 9'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_497 = 9'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_498 = 9'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_499 = 9'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_500 = 9'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@131668.4]
  assign _GEN_501 = 9'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@131668.4]
  assign io_out = 9'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@131668.4]
endmodule
module RegFile( // @[:@131670.2]
  input         clock, // @[:@131671.4]
  input         reset, // @[:@131672.4]
  input  [31:0] io_raddr, // @[:@131673.4]
  input         io_wen, // @[:@131673.4]
  input  [31:0] io_waddr, // @[:@131673.4]
  input  [63:0] io_wdata, // @[:@131673.4]
  output [63:0] io_rdata, // @[:@131673.4]
  input         io_reset, // @[:@131673.4]
  output [63:0] io_argIns_0, // @[:@131673.4]
  output [63:0] io_argIns_1, // @[:@131673.4]
  output [63:0] io_argIns_2, // @[:@131673.4]
  output [63:0] io_argIns_3, // @[:@131673.4]
  input         io_argOuts_0_valid, // @[:@131673.4]
  input  [63:0] io_argOuts_0_bits, // @[:@131673.4]
  input         io_argOuts_1_valid, // @[:@131673.4]
  input  [63:0] io_argOuts_1_bits // @[:@131673.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@133683.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@133683.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@133683.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@133683.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@133683.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@133683.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@133695.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@133695.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@133695.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@133695.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@133695.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@133695.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@133714.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@133714.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@133714.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@133714.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@133714.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@133714.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@133726.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@133726.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@133726.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@133726.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@133726.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@133726.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@133738.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@133738.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@133738.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@133738.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@133738.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@133738.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@133752.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@133752.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@133752.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@133752.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@133752.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@133752.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@133766.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@133766.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@133766.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@133766.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@133766.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@133766.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@133780.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@133780.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@133780.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@133780.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@133780.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@133780.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@133794.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@133794.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@133794.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@133794.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@133794.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@133794.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@133808.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@133808.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@133808.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@133808.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@133808.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@133808.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@133822.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@133822.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@133822.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@133822.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@133822.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@133822.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@133836.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@133836.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@133836.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@133836.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@133836.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@133836.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@133850.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@133850.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@133850.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@133850.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@133850.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@133850.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@133864.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@133864.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@133864.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@133864.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@133864.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@133864.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@133878.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@133878.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@133878.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@133878.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@133878.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@133878.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@133892.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@133892.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@133892.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@133892.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@133892.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@133892.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@133906.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@133906.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@133906.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@133906.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@133906.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@133906.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@133920.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@133920.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@133920.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@133920.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@133920.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@133920.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@133934.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@133934.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@133934.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@133934.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@133934.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@133934.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@133948.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@133948.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@133948.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@133948.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@133948.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@133948.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@133962.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@133962.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@133962.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@133962.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@133962.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@133962.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@133976.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@133976.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@133976.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@133976.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@133976.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@133976.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@133990.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@133990.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@133990.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@133990.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@133990.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@133990.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@134004.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@134004.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@134004.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@134004.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@134004.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@134004.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@134018.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@134018.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@134018.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@134018.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@134018.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@134018.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@134032.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@134032.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@134032.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@134032.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@134032.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@134032.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@134046.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@134046.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@134046.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@134046.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@134046.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@134046.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@134060.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@134060.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@134060.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@134060.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@134060.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@134060.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@134074.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@134074.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@134074.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@134074.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@134074.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@134074.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@134088.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@134088.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@134088.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@134088.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@134088.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@134088.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@134102.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@134102.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@134102.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@134102.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@134102.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@134102.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@134116.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@134116.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@134116.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@134116.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@134116.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@134116.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@134130.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@134130.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@134130.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@134130.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@134130.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@134130.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@134144.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@134144.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@134144.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@134144.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@134144.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@134144.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@134158.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@134158.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@134158.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@134158.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@134158.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@134158.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@134172.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@134172.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@134172.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@134172.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@134172.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@134172.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@134186.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@134186.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@134186.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@134186.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@134186.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@134186.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@134200.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@134200.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@134200.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@134200.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@134200.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@134200.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@134214.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@134214.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@134214.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@134214.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@134214.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@134214.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@134228.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@134228.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@134228.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@134228.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@134228.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@134228.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@134242.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@134242.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@134242.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@134242.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@134242.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@134242.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@134256.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@134256.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@134256.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@134256.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@134256.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@134256.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@134270.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@134270.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@134270.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@134270.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@134270.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@134270.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@134284.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@134284.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@134284.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@134284.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@134284.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@134284.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@134298.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@134298.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@134298.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@134298.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@134298.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@134298.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@134312.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@134312.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@134312.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@134312.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@134312.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@134312.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@134326.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@134326.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@134326.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@134326.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@134326.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@134326.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@134340.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@134340.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@134340.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@134340.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@134340.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@134340.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@134354.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@134354.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@134354.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@134354.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@134354.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@134354.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@134368.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@134368.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@134368.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@134368.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@134368.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@134368.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@134382.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@134382.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@134382.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@134382.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@134382.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@134382.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@134396.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@134396.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@134396.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@134396.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@134396.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@134396.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@134410.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@134410.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@134410.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@134410.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@134410.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@134410.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@134424.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@134424.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@134424.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@134424.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@134424.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@134424.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@134438.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@134438.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@134438.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@134438.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@134438.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@134438.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@134452.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@134452.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@134452.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@134452.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@134452.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@134452.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@134466.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@134466.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@134466.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@134466.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@134466.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@134466.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@134480.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@134480.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@134480.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@134480.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@134480.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@134480.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@134494.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@134494.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@134494.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@134494.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@134494.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@134494.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@134508.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@134508.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@134508.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@134508.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@134508.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@134508.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@134522.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@134522.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@134522.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@134522.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@134522.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@134522.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@134536.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@134536.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@134536.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@134536.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@134536.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@134536.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@134550.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@134550.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@134550.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@134550.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@134550.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@134550.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@134564.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@134564.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@134564.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@134564.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@134564.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@134564.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@134578.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@134578.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@134578.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@134578.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@134578.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@134578.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@134592.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@134592.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@134592.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@134592.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@134592.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@134592.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@134606.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@134606.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@134606.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@134606.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@134606.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@134606.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@134620.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@134620.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@134620.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@134620.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@134620.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@134620.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@134634.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@134634.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@134634.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@134634.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@134634.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@134634.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@134648.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@134648.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@134648.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@134648.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@134648.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@134648.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@134662.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@134662.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@134662.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@134662.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@134662.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@134662.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@134676.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@134676.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@134676.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@134676.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@134676.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@134676.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@134690.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@134690.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@134690.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@134690.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@134690.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@134690.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@134704.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@134704.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@134704.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@134704.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@134704.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@134704.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@134718.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@134718.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@134718.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@134718.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@134718.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@134718.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@134732.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@134732.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@134732.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@134732.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@134732.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@134732.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@134746.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@134746.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@134746.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@134746.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@134746.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@134746.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@134760.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@134760.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@134760.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@134760.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@134760.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@134760.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@134774.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@134774.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@134774.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@134774.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@134774.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@134774.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@134788.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@134788.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@134788.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@134788.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@134788.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@134788.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@134802.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@134802.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@134802.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@134802.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@134802.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@134802.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@134816.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@134816.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@134816.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@134816.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@134816.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@134816.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@134830.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@134830.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@134830.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@134830.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@134830.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@134830.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@134844.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@134844.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@134844.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@134844.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@134844.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@134844.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@134858.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@134858.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@134858.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@134858.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@134858.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@134858.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@134872.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@134872.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@134872.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@134872.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@134872.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@134872.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@134886.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@134886.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@134886.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@134886.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@134886.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@134886.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@134900.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@134900.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@134900.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@134900.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@134900.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@134900.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@134914.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@134914.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@134914.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@134914.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@134914.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@134914.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@134928.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@134928.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@134928.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@134928.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@134928.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@134928.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@134942.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@134942.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@134942.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@134942.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@134942.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@134942.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@134956.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@134956.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@134956.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@134956.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@134956.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@134956.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@134970.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@134970.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@134970.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@134970.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@134970.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@134970.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@134984.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@134984.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@134984.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@134984.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@134984.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@134984.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@134998.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@134998.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@134998.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@134998.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@134998.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@134998.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@135012.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@135012.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@135012.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@135012.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@135012.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@135012.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@135026.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@135026.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@135026.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@135026.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@135026.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@135026.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@135040.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@135040.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@135040.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@135040.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@135040.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@135040.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@135054.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@135054.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@135054.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@135054.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@135054.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@135054.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@135068.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@135068.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@135068.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@135068.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@135068.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@135068.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@135082.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@135082.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@135082.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@135082.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@135082.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@135082.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@135096.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@135096.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@135096.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@135096.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@135096.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@135096.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@135110.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@135110.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@135110.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@135110.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@135110.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@135110.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@135124.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@135124.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@135124.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@135124.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@135124.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@135124.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@135138.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@135138.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@135138.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@135138.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@135138.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@135138.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@135152.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@135152.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@135152.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@135152.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@135152.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@135152.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@135166.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@135166.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@135166.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@135166.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@135166.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@135166.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@135180.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@135180.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@135180.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@135180.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@135180.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@135180.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@135194.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@135194.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@135194.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@135194.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@135194.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@135194.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@135208.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@135208.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@135208.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@135208.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@135208.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@135208.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@135222.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@135222.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@135222.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@135222.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@135222.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@135222.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@135236.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@135236.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@135236.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@135236.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@135236.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@135236.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@135250.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@135250.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@135250.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@135250.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@135250.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@135250.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@135264.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@135264.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@135264.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@135264.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@135264.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@135264.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@135278.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@135278.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@135278.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@135278.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@135278.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@135278.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@135292.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@135292.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@135292.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@135292.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@135292.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@135292.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@135306.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@135306.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@135306.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@135306.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@135306.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@135306.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@135320.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@135320.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@135320.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@135320.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@135320.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@135320.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@135334.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@135334.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@135334.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@135334.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@135334.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@135334.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@135348.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@135348.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@135348.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@135348.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@135348.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@135348.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@135362.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@135362.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@135362.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@135362.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@135362.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@135362.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@135376.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@135376.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@135376.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@135376.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@135376.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@135376.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@135390.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@135390.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@135390.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@135390.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@135390.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@135390.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@135404.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@135404.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@135404.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@135404.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@135404.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@135404.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@135418.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@135418.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@135418.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@135418.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@135418.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@135418.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@135432.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@135432.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@135432.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@135432.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@135432.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@135432.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@135446.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@135446.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@135446.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@135446.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@135446.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@135446.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@135460.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@135460.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@135460.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@135460.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@135460.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@135460.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@135474.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@135474.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@135474.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@135474.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@135474.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@135474.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@135488.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@135488.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@135488.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@135488.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@135488.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@135488.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@135502.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@135502.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@135502.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@135502.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@135502.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@135502.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@135516.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@135516.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@135516.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@135516.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@135516.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@135516.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@135530.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@135530.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@135530.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@135530.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@135530.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@135530.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@135544.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@135544.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@135544.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@135544.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@135544.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@135544.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@135558.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@135558.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@135558.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@135558.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@135558.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@135558.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@135572.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@135572.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@135572.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@135572.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@135572.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@135572.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@135586.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@135586.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@135586.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@135586.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@135586.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@135586.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@135600.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@135600.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@135600.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@135600.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@135600.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@135600.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@135614.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@135614.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@135614.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@135614.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@135614.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@135614.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@135628.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@135628.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@135628.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@135628.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@135628.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@135628.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@135642.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@135642.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@135642.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@135642.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@135642.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@135642.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@135656.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@135656.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@135656.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@135656.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@135656.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@135656.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@135670.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@135670.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@135670.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@135670.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@135670.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@135670.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@135684.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@135684.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@135684.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@135684.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@135684.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@135684.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@135698.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@135698.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@135698.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@135698.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@135698.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@135698.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@135712.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@135712.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@135712.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@135712.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@135712.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@135712.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@135726.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@135726.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@135726.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@135726.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@135726.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@135726.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@135740.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@135740.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@135740.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@135740.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@135740.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@135740.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@135754.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@135754.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@135754.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@135754.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@135754.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@135754.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@135768.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@135768.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@135768.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@135768.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@135768.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@135768.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@135782.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@135782.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@135782.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@135782.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@135782.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@135782.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@135796.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@135796.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@135796.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@135796.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@135796.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@135796.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@135810.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@135810.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@135810.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@135810.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@135810.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@135810.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@135824.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@135824.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@135824.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@135824.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@135824.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@135824.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@135838.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@135838.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@135838.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@135838.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@135838.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@135838.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@135852.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@135852.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@135852.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@135852.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@135852.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@135852.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@135866.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@135866.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@135866.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@135866.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@135866.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@135866.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@135880.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@135880.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@135880.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@135880.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@135880.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@135880.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@135894.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@135894.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@135894.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@135894.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@135894.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@135894.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@135908.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@135908.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@135908.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@135908.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@135908.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@135908.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@135922.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@135922.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@135922.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@135922.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@135922.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@135922.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@135936.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@135936.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@135936.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@135936.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@135936.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@135936.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@135950.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@135950.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@135950.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@135950.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@135950.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@135950.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@135964.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@135964.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@135964.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@135964.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@135964.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@135964.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@135978.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@135978.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@135978.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@135978.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@135978.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@135978.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@135992.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@135992.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@135992.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@135992.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@135992.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@135992.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@136006.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@136006.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@136006.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@136006.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@136006.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@136006.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@136020.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@136020.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@136020.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@136020.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@136020.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@136020.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@136034.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@136034.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@136034.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@136034.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@136034.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@136034.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@136048.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@136048.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@136048.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@136048.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@136048.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@136048.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@136062.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@136062.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@136062.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@136062.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@136062.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@136062.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@136076.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@136076.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@136076.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@136076.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@136076.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@136076.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@136090.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@136090.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@136090.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@136090.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@136090.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@136090.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@136104.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@136104.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@136104.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@136104.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@136104.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@136104.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@136118.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@136118.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@136118.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@136118.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@136118.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@136118.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@136132.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@136132.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@136132.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@136132.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@136132.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@136132.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@136146.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@136146.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@136146.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@136146.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@136146.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@136146.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@136160.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@136160.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@136160.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@136160.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@136160.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@136160.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@136174.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@136174.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@136174.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@136174.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@136174.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@136174.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@136188.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@136188.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@136188.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@136188.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@136188.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@136188.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@136202.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@136202.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@136202.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@136202.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@136202.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@136202.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@136216.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@136216.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@136216.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@136216.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@136216.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@136216.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@136230.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@136230.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@136230.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@136230.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@136230.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@136230.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@136244.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@136244.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@136244.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@136244.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@136244.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@136244.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@136258.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@136258.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@136258.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@136258.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@136258.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@136258.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@136272.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@136272.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@136272.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@136272.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@136272.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@136272.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@136286.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@136286.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@136286.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@136286.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@136286.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@136286.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@136300.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@136300.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@136300.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@136300.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@136300.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@136300.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@136314.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@136314.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@136314.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@136314.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@136314.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@136314.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@136328.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@136328.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@136328.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@136328.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@136328.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@136328.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@136342.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@136342.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@136342.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@136342.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@136342.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@136342.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@136356.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@136356.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@136356.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@136356.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@136356.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@136356.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@136370.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@136370.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@136370.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@136370.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@136370.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@136370.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@136384.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@136384.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@136384.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@136384.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@136384.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@136384.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@136398.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@136398.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@136398.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@136398.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@136398.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@136398.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@136412.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@136412.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@136412.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@136412.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@136412.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@136412.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@136426.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@136426.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@136426.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@136426.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@136426.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@136426.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@136440.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@136440.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@136440.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@136440.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@136440.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@136440.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@136454.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@136454.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@136454.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@136454.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@136454.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@136454.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@136468.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@136468.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@136468.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@136468.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@136468.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@136468.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@136482.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@136482.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@136482.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@136482.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@136482.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@136482.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@136496.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@136496.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@136496.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@136496.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@136496.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@136496.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@136510.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@136510.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@136510.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@136510.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@136510.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@136510.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@136524.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@136524.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@136524.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@136524.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@136524.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@136524.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@136538.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@136538.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@136538.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@136538.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@136538.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@136538.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@136552.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@136552.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@136552.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@136552.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@136552.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@136552.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@136566.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@136566.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@136566.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@136566.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@136566.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@136566.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@136580.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@136580.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@136580.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@136580.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@136580.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@136580.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@136594.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@136594.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@136594.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@136594.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@136594.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@136594.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@136608.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@136608.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@136608.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@136608.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@136608.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@136608.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@136622.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@136622.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@136622.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@136622.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@136622.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@136622.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@136636.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@136636.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@136636.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@136636.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@136636.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@136636.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@136650.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@136650.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@136650.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@136650.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@136650.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@136650.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@136664.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@136664.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@136664.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@136664.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@136664.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@136664.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@136678.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@136678.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@136678.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@136678.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@136678.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@136678.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@136692.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@136692.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@136692.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@136692.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@136692.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@136692.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@136706.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@136706.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@136706.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@136706.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@136706.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@136706.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@136720.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@136720.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@136720.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@136720.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@136720.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@136720.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@136734.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@136734.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@136734.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@136734.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@136734.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@136734.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@136748.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@136748.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@136748.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@136748.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@136748.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@136748.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@136762.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@136762.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@136762.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@136762.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@136762.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@136762.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@136776.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@136776.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@136776.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@136776.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@136776.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@136776.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@136790.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@136790.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@136790.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@136790.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@136790.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@136790.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@136804.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@136804.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@136804.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@136804.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@136804.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@136804.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@136818.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@136818.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@136818.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@136818.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@136818.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@136818.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@136832.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@136832.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@136832.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@136832.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@136832.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@136832.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@136846.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@136846.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@136846.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@136846.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@136846.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@136846.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@136860.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@136860.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@136860.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@136860.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@136860.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@136860.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@136874.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@136874.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@136874.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@136874.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@136874.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@136874.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@136888.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@136888.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@136888.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@136888.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@136888.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@136888.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@136902.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@136902.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@136902.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@136902.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@136902.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@136902.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@136916.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@136916.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@136916.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@136916.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@136916.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@136916.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@136930.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@136930.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@136930.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@136930.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@136930.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@136930.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@136944.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@136944.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@136944.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@136944.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@136944.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@136944.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@136958.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@136958.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@136958.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@136958.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@136958.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@136958.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@136972.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@136972.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@136972.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@136972.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@136972.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@136972.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@136986.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@136986.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@136986.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@136986.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@136986.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@136986.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@137000.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@137000.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@137000.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@137000.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@137000.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@137000.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@137014.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@137014.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@137014.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@137014.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@137014.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@137014.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@137028.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@137028.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@137028.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@137028.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@137028.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@137028.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@137042.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@137042.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@137042.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@137042.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@137042.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@137042.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@137056.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@137056.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@137056.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@137056.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@137056.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@137056.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@137070.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@137070.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@137070.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@137070.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@137070.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@137070.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@137084.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@137084.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@137084.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@137084.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@137084.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@137084.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@137098.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@137098.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@137098.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@137098.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@137098.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@137098.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@137112.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@137112.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@137112.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@137112.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@137112.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@137112.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@137126.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@137126.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@137126.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@137126.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@137126.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@137126.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@137140.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@137140.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@137140.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@137140.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@137140.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@137140.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@137154.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@137154.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@137154.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@137154.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@137154.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@137154.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@137168.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@137168.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@137168.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@137168.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@137168.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@137168.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@137182.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@137182.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@137182.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@137182.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@137182.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@137182.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@137196.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@137196.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@137196.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@137196.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@137196.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@137196.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@137210.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@137210.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@137210.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@137210.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@137210.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@137210.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@137224.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@137224.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@137224.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@137224.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@137224.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@137224.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@137238.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@137238.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@137238.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@137238.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@137238.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@137238.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@137252.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@137252.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@137252.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@137252.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@137252.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@137252.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@137266.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@137266.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@137266.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@137266.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@137266.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@137266.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@137280.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@137280.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@137280.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@137280.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@137280.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@137280.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@137294.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@137294.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@137294.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@137294.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@137294.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@137294.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@137308.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@137308.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@137308.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@137308.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@137308.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@137308.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@137322.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@137322.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@137322.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@137322.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@137322.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@137322.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@137336.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@137336.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@137336.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@137336.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@137336.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@137336.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@137350.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@137350.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@137350.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@137350.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@137350.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@137350.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@137364.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@137364.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@137364.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@137364.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@137364.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@137364.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@137378.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@137378.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@137378.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@137378.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@137378.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@137378.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@137392.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@137392.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@137392.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@137392.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@137392.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@137392.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@137406.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@137406.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@137406.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@137406.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@137406.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@137406.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@137420.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@137420.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@137420.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@137420.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@137420.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@137420.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@137434.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@137434.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@137434.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@137434.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@137434.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@137434.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@137448.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@137448.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@137448.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@137448.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@137448.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@137448.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@137462.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@137462.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@137462.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@137462.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@137462.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@137462.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@137476.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@137476.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@137476.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@137476.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@137476.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@137476.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@137490.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@137490.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@137490.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@137490.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@137490.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@137490.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@137504.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@137504.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@137504.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@137504.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@137504.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@137504.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@137518.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@137518.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@137518.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@137518.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@137518.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@137518.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@137532.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@137532.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@137532.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@137532.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@137532.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@137532.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@137546.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@137546.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@137546.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@137546.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@137546.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@137546.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@137560.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@137560.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@137560.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@137560.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@137560.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@137560.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@137574.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@137574.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@137574.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@137574.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@137574.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@137574.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@137588.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@137588.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@137588.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@137588.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@137588.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@137588.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@137602.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@137602.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@137602.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@137602.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@137602.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@137602.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@137616.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@137616.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@137616.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@137616.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@137616.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@137616.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@137630.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@137630.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@137630.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@137630.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@137630.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@137630.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@137644.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@137644.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@137644.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@137644.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@137644.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@137644.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@137658.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@137658.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@137658.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@137658.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@137658.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@137658.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@137672.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@137672.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@137672.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@137672.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@137672.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@137672.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@137686.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@137686.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@137686.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@137686.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@137686.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@137686.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@137700.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@137700.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@137700.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@137700.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@137700.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@137700.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@137714.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@137714.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@137714.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@137714.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@137714.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@137714.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@137728.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@137728.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@137728.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@137728.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@137728.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@137728.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@137742.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@137742.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@137742.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@137742.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@137742.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@137742.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@137756.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@137756.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@137756.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@137756.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@137756.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@137756.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@137770.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@137770.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@137770.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@137770.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@137770.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@137770.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@137784.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@137784.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@137784.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@137784.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@137784.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@137784.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@137798.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@137798.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@137798.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@137798.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@137798.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@137798.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@137812.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@137812.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@137812.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@137812.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@137812.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@137812.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@137826.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@137826.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@137826.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@137826.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@137826.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@137826.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@137840.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@137840.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@137840.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@137840.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@137840.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@137840.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@137854.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@137854.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@137854.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@137854.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@137854.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@137854.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@137868.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@137868.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@137868.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@137868.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@137868.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@137868.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@137882.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@137882.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@137882.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@137882.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@137882.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@137882.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@137896.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@137896.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@137896.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@137896.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@137896.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@137896.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@137910.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@137910.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@137910.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@137910.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@137910.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@137910.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@137924.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@137924.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@137924.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@137924.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@137924.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@137924.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@137938.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@137938.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@137938.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@137938.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@137938.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@137938.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@137952.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@137952.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@137952.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@137952.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@137952.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@137952.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@137966.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@137966.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@137966.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@137966.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@137966.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@137966.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@137980.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@137980.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@137980.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@137980.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@137980.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@137980.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@137994.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@137994.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@137994.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@137994.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@137994.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@137994.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@138008.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@138008.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@138008.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@138008.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@138008.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@138008.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@138022.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@138022.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@138022.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@138022.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@138022.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@138022.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@138036.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@138036.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@138036.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@138036.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@138036.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@138036.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@138050.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@138050.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@138050.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@138050.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@138050.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@138050.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@138064.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@138064.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@138064.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@138064.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@138064.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@138064.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@138078.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@138078.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@138078.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@138078.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@138078.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@138078.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@138092.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@138092.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@138092.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@138092.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@138092.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@138092.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@138106.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@138106.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@138106.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@138106.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@138106.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@138106.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@138120.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@138120.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@138120.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@138120.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@138120.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@138120.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@138134.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@138134.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@138134.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@138134.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@138134.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@138134.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@138148.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@138148.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@138148.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@138148.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@138148.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@138148.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@138162.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@138162.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@138162.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@138162.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@138162.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@138162.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@138176.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@138176.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@138176.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@138176.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@138176.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@138176.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@138190.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@138190.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@138190.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@138190.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@138190.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@138190.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@138204.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@138204.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@138204.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@138204.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@138204.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@138204.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@138218.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@138218.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@138218.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@138218.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@138218.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@138218.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@138232.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@138232.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@138232.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@138232.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@138232.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@138232.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@138246.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@138246.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@138246.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@138246.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@138246.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@138246.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@138260.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@138260.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@138260.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@138260.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@138260.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@138260.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@138274.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@138274.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@138274.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@138274.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@138274.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@138274.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@138288.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@138288.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@138288.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@138288.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@138288.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@138288.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@138302.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@138302.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@138302.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@138302.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@138302.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@138302.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@138316.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@138316.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@138316.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@138316.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@138316.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@138316.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@138330.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@138330.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@138330.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@138330.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@138330.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@138330.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@138344.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@138344.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@138344.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@138344.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@138344.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@138344.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@138358.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@138358.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@138358.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@138358.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@138358.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@138358.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@138372.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@138372.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@138372.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@138372.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@138372.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@138372.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@138386.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@138386.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@138386.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@138386.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@138386.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@138386.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@138400.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@138400.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@138400.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@138400.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@138400.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@138400.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@138414.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@138414.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@138414.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@138414.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@138414.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@138414.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@138428.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@138428.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@138428.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@138428.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@138428.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@138428.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@138442.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@138442.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@138442.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@138442.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@138442.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@138442.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@138456.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@138456.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@138456.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@138456.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@138456.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@138456.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@138470.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@138470.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@138470.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@138470.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@138470.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@138470.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@138484.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@138484.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@138484.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@138484.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@138484.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@138484.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@138498.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@138498.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@138498.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@138498.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@138498.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@138498.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@138512.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@138512.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@138512.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@138512.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@138512.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@138512.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@138526.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@138526.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@138526.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@138526.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@138526.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@138526.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@138540.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@138540.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@138540.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@138540.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@138540.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@138540.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@138554.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@138554.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@138554.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@138554.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@138554.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@138554.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@138568.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@138568.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@138568.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@138568.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@138568.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@138568.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@138582.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@138582.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@138582.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@138582.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@138582.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@138582.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@138596.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@138596.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@138596.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@138596.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@138596.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@138596.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@138610.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@138610.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@138610.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@138610.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@138610.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@138610.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@138624.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@138624.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@138624.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@138624.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@138624.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@138624.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@138638.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@138638.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@138638.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@138638.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@138638.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@138638.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@138652.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@138652.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@138652.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@138652.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@138652.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@138652.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@138666.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@138666.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@138666.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@138666.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@138666.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@138666.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@138680.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@138680.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@138680.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@138680.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@138680.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@138680.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@138694.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@138694.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@138694.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@138694.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@138694.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@138694.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@138708.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@138708.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@138708.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@138708.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@138708.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@138708.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@138722.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@138722.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@138722.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@138722.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@138722.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@138722.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@138736.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@138736.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@138736.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@138736.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@138736.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@138736.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@138750.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@138750.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@138750.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@138750.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@138750.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@138750.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@138764.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@138764.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@138764.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@138764.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@138764.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@138764.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@138778.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@138778.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@138778.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@138778.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@138778.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@138778.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@138792.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@138792.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@138792.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@138792.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@138792.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@138792.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@138806.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@138806.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@138806.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@138806.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@138806.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@138806.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@138820.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@138820.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@138820.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@138820.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@138820.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@138820.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@138834.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@138834.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@138834.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@138834.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@138834.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@138834.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@138848.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@138848.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@138848.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@138848.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@138848.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@138848.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@138862.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@138862.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@138862.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@138862.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@138862.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@138862.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@138876.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@138876.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@138876.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@138876.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@138876.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@138876.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@138890.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@138890.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@138890.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@138890.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@138890.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@138890.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@138904.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@138904.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@138904.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@138904.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@138904.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@138904.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@138918.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@138918.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@138918.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@138918.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@138918.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@138918.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@138932.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@138932.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@138932.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@138932.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@138932.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@138932.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@138946.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@138946.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@138946.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@138946.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@138946.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@138946.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@138960.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@138960.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@138960.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@138960.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@138960.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@138960.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@138974.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@138974.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@138974.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@138974.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@138974.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@138974.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@138988.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@138988.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@138988.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@138988.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@138988.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@138988.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@139002.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@139002.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@139002.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@139002.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@139002.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@139002.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@139016.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@139016.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@139016.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@139016.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@139016.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@139016.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@139030.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@139030.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@139030.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@139030.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@139030.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@139030.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@139044.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@139044.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@139044.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@139044.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@139044.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@139044.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@139058.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@139058.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@139058.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@139058.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@139058.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@139058.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@139072.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@139072.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@139072.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@139072.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@139072.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@139072.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@139086.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@139086.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@139086.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@139086.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@139086.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@139086.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@139100.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@139100.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@139100.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@139100.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@139100.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@139100.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@139114.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@139114.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@139114.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@139114.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@139114.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@139114.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@139128.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@139128.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@139128.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@139128.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@139128.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@139128.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@139142.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@139142.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@139142.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@139142.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@139142.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@139142.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@139156.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@139156.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@139156.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@139156.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@139156.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@139156.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@139170.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@139170.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@139170.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@139170.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@139170.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@139170.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@139184.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@139184.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@139184.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@139184.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@139184.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@139184.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@139198.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@139198.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@139198.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@139198.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@139198.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@139198.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@139212.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@139212.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@139212.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@139212.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@139212.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@139212.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@139226.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@139226.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@139226.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@139226.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@139226.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@139226.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@139240.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@139240.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@139240.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@139240.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@139240.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@139240.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@139254.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@139254.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@139254.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@139254.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@139254.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@139254.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@139268.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@139268.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@139268.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@139268.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@139268.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@139268.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@139282.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@139282.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@139282.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@139282.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@139282.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@139282.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@139296.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@139296.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@139296.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@139296.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@139296.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@139296.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@139310.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@139310.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@139310.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@139310.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@139310.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@139310.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@139324.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@139324.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@139324.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@139324.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@139324.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@139324.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@139338.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@139338.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@139338.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@139338.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@139338.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@139338.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@139352.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@139352.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@139352.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@139352.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@139352.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@139352.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@139366.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@139366.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@139366.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@139366.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@139366.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@139366.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@139380.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@139380.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@139380.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@139380.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@139380.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@139380.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@139394.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@139394.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@139394.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@139394.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@139394.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@139394.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@139408.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@139408.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@139408.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@139408.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@139408.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@139408.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@139422.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@139422.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@139422.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@139422.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@139422.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@139422.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@139436.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@139436.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@139436.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@139436.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@139436.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@139436.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@139450.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@139450.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@139450.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@139450.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@139450.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@139450.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@139464.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@139464.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@139464.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@139464.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@139464.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@139464.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@139478.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@139478.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@139478.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@139478.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@139478.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@139478.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@139492.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@139492.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@139492.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@139492.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@139492.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@139492.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@139506.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@139506.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@139506.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@139506.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@139506.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@139506.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@139520.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@139520.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@139520.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@139520.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@139520.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@139520.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@139534.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@139534.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@139534.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@139534.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@139534.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@139534.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@139548.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@139548.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@139548.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@139548.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@139548.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@139548.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@139562.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@139562.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@139562.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@139562.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@139562.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@139562.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@139576.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@139576.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@139576.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@139576.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@139576.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@139576.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@139590.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@139590.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@139590.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@139590.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@139590.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@139590.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@139604.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@139604.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@139604.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@139604.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@139604.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@139604.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@139618.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@139618.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@139618.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@139618.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@139618.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@139618.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@139632.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@139632.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@139632.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@139632.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@139632.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@139632.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@139646.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@139646.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@139646.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@139646.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@139646.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@139646.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@139660.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@139660.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@139660.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@139660.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@139660.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@139660.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@139674.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@139674.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@139674.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@139674.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@139674.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@139674.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@139688.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@139688.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@139688.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@139688.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@139688.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@139688.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@139702.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@139702.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@139702.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@139702.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@139702.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@139702.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@139716.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@139716.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@139716.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@139716.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@139716.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@139716.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@139730.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@139730.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@139730.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@139730.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@139730.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@139730.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@139744.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@139744.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@139744.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@139744.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@139744.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@139744.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@139758.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@139758.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@139758.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@139758.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@139758.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@139758.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@139772.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@139772.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@139772.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@139772.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@139772.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@139772.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@139786.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@139786.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@139786.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@139786.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@139786.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@139786.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@139800.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@139800.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@139800.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@139800.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@139800.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@139800.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@139814.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@139814.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@139814.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@139814.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@139814.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@139814.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@139828.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@139828.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@139828.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@139828.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@139828.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@139828.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@139842.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@139842.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@139842.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@139842.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@139842.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@139842.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@139856.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@139856.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@139856.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@139856.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@139856.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@139856.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@139870.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@139870.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@139870.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@139870.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@139870.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@139870.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@139884.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@139884.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@139884.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@139884.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@139884.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@139884.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@139898.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@139898.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@139898.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@139898.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@139898.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@139898.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@139912.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@139912.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@139912.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@139912.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@139912.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@139912.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@139926.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@139926.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@139926.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@139926.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@139926.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@139926.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@139940.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@139940.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@139940.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@139940.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@139940.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@139940.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@139954.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@139954.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@139954.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@139954.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@139954.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@139954.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@139968.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@139968.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@139968.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@139968.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@139968.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@139968.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@139982.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@139982.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@139982.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@139982.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@139982.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@139982.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@139996.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@139996.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@139996.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@139996.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@139996.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@139996.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@140010.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@140010.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@140010.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@140010.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@140010.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@140010.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@140024.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@140024.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@140024.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@140024.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@140024.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@140024.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@140038.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@140038.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@140038.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@140038.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@140038.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@140038.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@140052.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@140052.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@140052.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@140052.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@140052.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@140052.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@140066.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@140066.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@140066.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@140066.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@140066.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@140066.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@140080.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@140080.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@140080.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@140080.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@140080.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@140080.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@140094.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@140094.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@140094.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@140094.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@140094.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@140094.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@140108.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@140108.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@140108.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@140108.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@140108.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@140108.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@140122.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@140122.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@140122.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@140122.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@140122.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@140122.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@140136.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@140136.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@140136.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@140136.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@140136.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@140136.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@140150.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@140150.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@140150.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@140150.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@140150.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@140150.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@140164.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@140164.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@140164.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@140164.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@140164.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@140164.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@140178.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@140178.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@140178.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@140178.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@140178.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@140178.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@140192.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@140192.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@140192.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@140192.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@140192.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@140192.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@140206.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@140206.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@140206.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@140206.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@140206.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@140206.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@140220.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@140220.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@140220.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@140220.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@140220.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@140220.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@140234.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@140234.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@140234.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@140234.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@140234.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@140234.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@140248.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@140248.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@140248.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@140248.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@140248.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@140248.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@140262.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@140262.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@140262.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@140262.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@140262.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@140262.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@140276.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@140276.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@140276.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@140276.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@140276.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@140276.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@140290.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@140290.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@140290.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@140290.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@140290.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@140290.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@140304.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@140304.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@140304.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@140304.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@140304.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@140304.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@140318.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@140318.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@140318.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@140318.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@140318.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@140318.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@140332.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@140332.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@140332.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@140332.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@140332.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@140332.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@140346.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@140346.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@140346.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@140346.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@140346.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@140346.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@140360.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@140360.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@140360.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@140360.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@140360.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@140360.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@140374.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@140374.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@140374.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@140374.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@140374.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@140374.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@140388.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@140388.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@140388.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@140388.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@140388.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@140388.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@140402.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@140402.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@140402.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@140402.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@140402.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@140402.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@140416.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@140416.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@140416.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@140416.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@140416.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@140416.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@140430.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@140430.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@140430.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@140430.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@140430.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@140430.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@140444.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@140444.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@140444.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@140444.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@140444.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@140444.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@140458.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@140458.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@140458.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@140458.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@140458.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@140458.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@140472.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@140472.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@140472.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@140472.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@140472.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@140472.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@140486.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@140486.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@140486.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@140486.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@140486.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@140486.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@140500.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@140500.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@140500.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@140500.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@140500.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@140500.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@140514.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@140514.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@140514.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@140514.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@140514.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@140514.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@140528.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@140528.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@140528.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@140528.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@140528.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@140528.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@140542.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@140542.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@140542.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@140542.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@140542.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@140542.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@140556.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@140556.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@140556.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@140556.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@140556.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@140556.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@140570.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@140570.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@140570.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@140570.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@140570.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@140570.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@140584.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@140584.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@140584.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@140584.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@140584.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@140584.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@140598.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@140598.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@140598.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@140598.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@140598.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@140598.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@140612.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@140612.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@140612.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@140612.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@140612.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@140612.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@140626.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@140626.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@140626.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@140626.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@140626.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@140626.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@140640.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@140640.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@140640.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@140640.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@140640.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@140640.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@140654.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@140654.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@140654.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@140654.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@140654.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@140654.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@140668.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@140668.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@140668.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@140668.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@140668.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@140668.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@140682.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@140682.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@140682.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@140682.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@140682.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@140682.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@140696.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@140696.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@140696.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@140696.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@140696.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@140696.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@140710.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@140710.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@140710.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@140710.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@140710.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@140710.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@140724.4]
  wire [8:0] rport_io_sel; // @[RegFile.scala 95:21:@140724.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@140724.4]
  wire  _T_3078; // @[RegFile.scala 80:42:@133686.4]
  wire  _T_3084; // @[RegFile.scala 68:46:@133698.4]
  wire  _T_3085; // @[RegFile.scala 68:34:@133699.4]
  wire  _T_3098; // @[RegFile.scala 80:42:@133717.4]
  wire  _T_3104; // @[RegFile.scala 80:42:@133729.4]
  wire  _T_3110; // @[RegFile.scala 74:80:@133741.4]
  wire  _T_3111; // @[RegFile.scala 74:68:@133742.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@133683.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@133695.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@133714.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@133726.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@133738.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@133752.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@133766.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@133780.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@133794.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@133808.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@133822.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@133836.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@133850.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@133864.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@133878.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@133892.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@133906.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@133920.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@133934.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@133948.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@133962.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@133976.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@133990.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@134004.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@134018.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@134032.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@134046.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@134060.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@134074.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@134088.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@134102.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@134116.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@134130.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@134144.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@134158.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@134172.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@134186.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@134200.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@134214.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@134228.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@134242.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@134256.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@134270.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@134284.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@134298.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@134312.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@134326.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@134340.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@134354.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@134368.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@134382.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@134396.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@134410.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@134424.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@134438.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@134452.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@134466.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@134480.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@134494.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@134508.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@134522.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@134536.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@134550.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@134564.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@134578.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@134592.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@134606.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@134620.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@134634.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@134648.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@134662.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@134676.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@134690.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@134704.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@134718.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@134732.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@134746.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@134760.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@134774.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@134788.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@134802.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@134816.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@134830.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@134844.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@134858.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@134872.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@134886.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@134900.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@134914.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@134928.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@134942.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@134956.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@134970.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@134984.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@134998.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@135012.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@135026.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@135040.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@135054.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@135068.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@135082.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@135096.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@135110.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@135124.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@135138.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@135152.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@135166.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@135180.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@135194.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@135208.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@135222.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@135236.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@135250.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@135264.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@135278.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@135292.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@135306.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@135320.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@135334.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@135348.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@135362.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@135376.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@135390.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@135404.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@135418.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@135432.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@135446.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@135460.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@135474.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@135488.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@135502.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@135516.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@135530.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@135544.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@135558.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@135572.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@135586.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@135600.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@135614.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@135628.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@135642.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@135656.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@135670.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@135684.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@135698.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@135712.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@135726.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@135740.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@135754.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@135768.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@135782.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@135796.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@135810.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@135824.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@135838.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@135852.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@135866.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@135880.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@135894.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@135908.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@135922.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@135936.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@135950.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@135964.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@135978.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@135992.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@136006.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@136020.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@136034.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@136048.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@136062.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@136076.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@136090.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@136104.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@136118.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@136132.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@136146.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@136160.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@136174.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@136188.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@136202.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@136216.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@136230.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@136244.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@136258.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@136272.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@136286.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@136300.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@136314.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@136328.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@136342.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@136356.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@136370.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@136384.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@136398.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@136412.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@136426.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@136440.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@136454.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@136468.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@136482.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@136496.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@136510.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@136524.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@136538.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@136552.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@136566.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@136580.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@136594.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@136608.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@136622.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@136636.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@136650.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@136664.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@136678.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@136692.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@136706.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@136720.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@136734.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@136748.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@136762.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@136776.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@136790.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@136804.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@136818.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@136832.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@136846.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@136860.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@136874.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@136888.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@136902.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@136916.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@136930.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@136944.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@136958.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@136972.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@136986.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@137000.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@137014.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@137028.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@137042.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@137056.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@137070.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@137084.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@137098.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@137112.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@137126.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@137140.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@137154.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@137168.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@137182.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@137196.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@137210.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@137224.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@137238.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@137252.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@137266.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@137280.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@137294.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@137308.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@137322.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@137336.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@137350.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@137364.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@137378.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@137392.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@137406.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@137420.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@137434.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@137448.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@137462.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@137476.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@137490.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@137504.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@137518.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@137532.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@137546.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@137560.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@137574.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@137588.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@137602.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@137616.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@137630.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@137644.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@137658.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@137672.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@137686.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@137700.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@137714.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@137728.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@137742.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@137756.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@137770.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@137784.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@137798.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@137812.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@137826.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@137840.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@137854.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@137868.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@137882.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@137896.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@137910.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@137924.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@137938.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@137952.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@137966.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@137980.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@137994.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@138008.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@138022.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@138036.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@138050.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@138064.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@138078.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@138092.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@138106.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@138120.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@138134.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@138148.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@138162.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@138176.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@138190.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@138204.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@138218.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@138232.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@138246.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@138260.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@138274.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@138288.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@138302.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@138316.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@138330.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@138344.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@138358.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@138372.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@138386.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@138400.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@138414.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@138428.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@138442.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@138456.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@138470.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@138484.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@138498.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@138512.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@138526.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@138540.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@138554.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@138568.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@138582.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@138596.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@138610.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@138624.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@138638.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@138652.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@138666.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@138680.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@138694.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@138708.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@138722.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@138736.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@138750.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@138764.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@138778.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@138792.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@138806.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@138820.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@138834.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@138848.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@138862.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@138876.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@138890.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@138904.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@138918.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@138932.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@138946.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@138960.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@138974.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@138988.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@139002.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@139016.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@139030.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@139044.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@139058.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@139072.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@139086.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@139100.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@139114.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@139128.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@139142.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@139156.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@139170.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@139184.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@139198.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@139212.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@139226.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@139240.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@139254.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@139268.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@139282.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@139296.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@139310.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@139324.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@139338.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@139352.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@139366.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@139380.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@139394.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@139408.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@139422.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@139436.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@139450.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@139464.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@139478.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@139492.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@139506.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@139520.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@139534.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@139548.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@139562.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@139576.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@139590.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@139604.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@139618.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@139632.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@139646.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@139660.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@139674.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@139688.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@139702.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@139716.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@139730.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@139744.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@139758.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@139772.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@139786.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@139800.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@139814.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@139828.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@139842.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@139856.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@139870.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@139884.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@139898.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@139912.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@139926.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@139940.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@139954.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@139968.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@139982.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@139996.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@140010.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@140024.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@140038.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@140052.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@140066.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@140080.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@140094.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@140108.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@140122.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@140136.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@140150.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@140164.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@140178.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@140192.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@140206.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@140220.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@140234.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@140248.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@140262.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@140276.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@140290.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@140304.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@140318.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@140332.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@140346.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@140360.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@140374.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@140388.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@140402.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@140416.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@140430.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@140444.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@140458.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@140472.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@140486.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@140500.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@140514.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@140528.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@140542.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@140556.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@140570.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@140584.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@140598.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@140612.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@140626.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@140640.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@140654.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@140668.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@140682.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@140696.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@140710.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  MuxN rport ( // @[RegFile.scala 95:21:@140724.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3078 = io_waddr == 32'h0; // @[RegFile.scala 80:42:@133686.4]
  assign _T_3084 = io_waddr == 32'h1; // @[RegFile.scala 68:46:@133698.4]
  assign _T_3085 = io_wen & _T_3084; // @[RegFile.scala 68:34:@133699.4]
  assign _T_3098 = io_waddr == 32'h2; // @[RegFile.scala 80:42:@133717.4]
  assign _T_3104 = io_waddr == 32'h3; // @[RegFile.scala 80:42:@133729.4]
  assign _T_3110 = io_waddr == 32'h4; // @[RegFile.scala 74:80:@133741.4]
  assign _T_3111 = io_wen & _T_3110; // @[RegFile.scala 74:68:@133742.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@141735.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@141741.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@141742.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@141743.4]
  assign io_argIns_3 = regs_3_io_out; // @[RegFile.scala 111:13:@141744.4]
  assign regs_0_clock = clock; // @[:@133684.4]
  assign regs_0_reset = reset; // @[:@133685.4 RegFile.scala 82:16:@133691.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@133689.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@133693.4]
  assign regs_0_io_enable = io_wen & _T_3078; // @[RegFile.scala 80:20:@133688.4]
  assign regs_1_clock = clock; // @[:@133696.4]
  assign regs_1_reset = reset; // @[:@133697.4 RegFile.scala 70:16:@133709.4]
  assign regs_1_io_in = _T_3085 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@133707.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@133712.4]
  assign regs_1_io_enable = _T_3085 ? _T_3085 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@133703.4]
  assign regs_2_clock = clock; // @[:@133715.4]
  assign regs_2_reset = reset; // @[:@133716.4 RegFile.scala 82:16:@133722.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@133720.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@133724.4]
  assign regs_2_io_enable = io_wen & _T_3098; // @[RegFile.scala 80:20:@133719.4]
  assign regs_3_clock = clock; // @[:@133727.4]
  assign regs_3_reset = reset; // @[:@133728.4 RegFile.scala 82:16:@133734.4]
  assign regs_3_io_in = io_wdata; // @[RegFile.scala 81:16:@133732.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 83:19:@133736.4]
  assign regs_3_io_enable = io_wen & _T_3104; // @[RegFile.scala 80:20:@133731.4]
  assign regs_4_clock = clock; // @[:@133739.4]
  assign regs_4_reset = io_reset; // @[:@133740.4 RegFile.scala 76:16:@133747.4]
  assign regs_4_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@133746.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@133750.4]
  assign regs_4_io_enable = io_argOuts_1_valid | _T_3111; // @[RegFile.scala 74:20:@133744.4]
  assign regs_5_clock = clock; // @[:@133753.4]
  assign regs_5_reset = io_reset; // @[:@133754.4 RegFile.scala 76:16:@133761.4]
  assign regs_5_io_in = 64'h0; // @[RegFile.scala 75:16:@133760.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@133764.4]
  assign regs_5_io_enable = 1'h1; // @[RegFile.scala 74:20:@133758.4]
  assign regs_6_clock = clock; // @[:@133767.4]
  assign regs_6_reset = io_reset; // @[:@133768.4 RegFile.scala 76:16:@133775.4]
  assign regs_6_io_in = 64'h0; // @[RegFile.scala 75:16:@133774.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@133778.4]
  assign regs_6_io_enable = 1'h1; // @[RegFile.scala 74:20:@133772.4]
  assign regs_7_clock = clock; // @[:@133781.4]
  assign regs_7_reset = io_reset; // @[:@133782.4 RegFile.scala 76:16:@133789.4]
  assign regs_7_io_in = 64'h0; // @[RegFile.scala 75:16:@133788.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@133792.4]
  assign regs_7_io_enable = 1'h1; // @[RegFile.scala 74:20:@133786.4]
  assign regs_8_clock = clock; // @[:@133795.4]
  assign regs_8_reset = io_reset; // @[:@133796.4 RegFile.scala 76:16:@133803.4]
  assign regs_8_io_in = 64'h0; // @[RegFile.scala 75:16:@133802.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@133806.4]
  assign regs_8_io_enable = 1'h1; // @[RegFile.scala 74:20:@133800.4]
  assign regs_9_clock = clock; // @[:@133809.4]
  assign regs_9_reset = io_reset; // @[:@133810.4 RegFile.scala 76:16:@133817.4]
  assign regs_9_io_in = 64'h0; // @[RegFile.scala 75:16:@133816.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@133820.4]
  assign regs_9_io_enable = 1'h1; // @[RegFile.scala 74:20:@133814.4]
  assign regs_10_clock = clock; // @[:@133823.4]
  assign regs_10_reset = io_reset; // @[:@133824.4 RegFile.scala 76:16:@133831.4]
  assign regs_10_io_in = 64'h0; // @[RegFile.scala 75:16:@133830.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@133834.4]
  assign regs_10_io_enable = 1'h1; // @[RegFile.scala 74:20:@133828.4]
  assign regs_11_clock = clock; // @[:@133837.4]
  assign regs_11_reset = io_reset; // @[:@133838.4 RegFile.scala 76:16:@133845.4]
  assign regs_11_io_in = 64'h0; // @[RegFile.scala 75:16:@133844.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@133848.4]
  assign regs_11_io_enable = 1'h1; // @[RegFile.scala 74:20:@133842.4]
  assign regs_12_clock = clock; // @[:@133851.4]
  assign regs_12_reset = io_reset; // @[:@133852.4 RegFile.scala 76:16:@133859.4]
  assign regs_12_io_in = 64'h0; // @[RegFile.scala 75:16:@133858.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@133862.4]
  assign regs_12_io_enable = 1'h1; // @[RegFile.scala 74:20:@133856.4]
  assign regs_13_clock = clock; // @[:@133865.4]
  assign regs_13_reset = io_reset; // @[:@133866.4 RegFile.scala 76:16:@133873.4]
  assign regs_13_io_in = 64'h0; // @[RegFile.scala 75:16:@133872.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@133876.4]
  assign regs_13_io_enable = 1'h1; // @[RegFile.scala 74:20:@133870.4]
  assign regs_14_clock = clock; // @[:@133879.4]
  assign regs_14_reset = io_reset; // @[:@133880.4 RegFile.scala 76:16:@133887.4]
  assign regs_14_io_in = 64'h0; // @[RegFile.scala 75:16:@133886.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@133890.4]
  assign regs_14_io_enable = 1'h1; // @[RegFile.scala 74:20:@133884.4]
  assign regs_15_clock = clock; // @[:@133893.4]
  assign regs_15_reset = io_reset; // @[:@133894.4 RegFile.scala 76:16:@133901.4]
  assign regs_15_io_in = 64'h0; // @[RegFile.scala 75:16:@133900.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@133904.4]
  assign regs_15_io_enable = 1'h1; // @[RegFile.scala 74:20:@133898.4]
  assign regs_16_clock = clock; // @[:@133907.4]
  assign regs_16_reset = io_reset; // @[:@133908.4 RegFile.scala 76:16:@133915.4]
  assign regs_16_io_in = 64'h0; // @[RegFile.scala 75:16:@133914.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@133918.4]
  assign regs_16_io_enable = 1'h1; // @[RegFile.scala 74:20:@133912.4]
  assign regs_17_clock = clock; // @[:@133921.4]
  assign regs_17_reset = io_reset; // @[:@133922.4 RegFile.scala 76:16:@133929.4]
  assign regs_17_io_in = 64'h0; // @[RegFile.scala 75:16:@133928.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@133932.4]
  assign regs_17_io_enable = 1'h1; // @[RegFile.scala 74:20:@133926.4]
  assign regs_18_clock = clock; // @[:@133935.4]
  assign regs_18_reset = io_reset; // @[:@133936.4 RegFile.scala 76:16:@133943.4]
  assign regs_18_io_in = 64'h0; // @[RegFile.scala 75:16:@133942.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@133946.4]
  assign regs_18_io_enable = 1'h1; // @[RegFile.scala 74:20:@133940.4]
  assign regs_19_clock = clock; // @[:@133949.4]
  assign regs_19_reset = io_reset; // @[:@133950.4 RegFile.scala 76:16:@133957.4]
  assign regs_19_io_in = 64'h0; // @[RegFile.scala 75:16:@133956.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@133960.4]
  assign regs_19_io_enable = 1'h1; // @[RegFile.scala 74:20:@133954.4]
  assign regs_20_clock = clock; // @[:@133963.4]
  assign regs_20_reset = io_reset; // @[:@133964.4 RegFile.scala 76:16:@133971.4]
  assign regs_20_io_in = 64'h0; // @[RegFile.scala 75:16:@133970.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@133974.4]
  assign regs_20_io_enable = 1'h1; // @[RegFile.scala 74:20:@133968.4]
  assign regs_21_clock = clock; // @[:@133977.4]
  assign regs_21_reset = io_reset; // @[:@133978.4 RegFile.scala 76:16:@133985.4]
  assign regs_21_io_in = 64'h0; // @[RegFile.scala 75:16:@133984.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@133988.4]
  assign regs_21_io_enable = 1'h1; // @[RegFile.scala 74:20:@133982.4]
  assign regs_22_clock = clock; // @[:@133991.4]
  assign regs_22_reset = io_reset; // @[:@133992.4 RegFile.scala 76:16:@133999.4]
  assign regs_22_io_in = 64'h0; // @[RegFile.scala 75:16:@133998.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@134002.4]
  assign regs_22_io_enable = 1'h1; // @[RegFile.scala 74:20:@133996.4]
  assign regs_23_clock = clock; // @[:@134005.4]
  assign regs_23_reset = io_reset; // @[:@134006.4 RegFile.scala 76:16:@134013.4]
  assign regs_23_io_in = 64'h0; // @[RegFile.scala 75:16:@134012.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@134016.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 74:20:@134010.4]
  assign regs_24_clock = clock; // @[:@134019.4]
  assign regs_24_reset = io_reset; // @[:@134020.4 RegFile.scala 76:16:@134027.4]
  assign regs_24_io_in = 64'h0; // @[RegFile.scala 75:16:@134026.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@134030.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 74:20:@134024.4]
  assign regs_25_clock = clock; // @[:@134033.4]
  assign regs_25_reset = io_reset; // @[:@134034.4 RegFile.scala 76:16:@134041.4]
  assign regs_25_io_in = 64'h0; // @[RegFile.scala 75:16:@134040.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@134044.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 74:20:@134038.4]
  assign regs_26_clock = clock; // @[:@134047.4]
  assign regs_26_reset = io_reset; // @[:@134048.4 RegFile.scala 76:16:@134055.4]
  assign regs_26_io_in = 64'h0; // @[RegFile.scala 75:16:@134054.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@134058.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 74:20:@134052.4]
  assign regs_27_clock = clock; // @[:@134061.4]
  assign regs_27_reset = io_reset; // @[:@134062.4 RegFile.scala 76:16:@134069.4]
  assign regs_27_io_in = 64'h0; // @[RegFile.scala 75:16:@134068.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@134072.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 74:20:@134066.4]
  assign regs_28_clock = clock; // @[:@134075.4]
  assign regs_28_reset = io_reset; // @[:@134076.4 RegFile.scala 76:16:@134083.4]
  assign regs_28_io_in = 64'h0; // @[RegFile.scala 75:16:@134082.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@134086.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 74:20:@134080.4]
  assign regs_29_clock = clock; // @[:@134089.4]
  assign regs_29_reset = io_reset; // @[:@134090.4 RegFile.scala 76:16:@134097.4]
  assign regs_29_io_in = 64'h0; // @[RegFile.scala 75:16:@134096.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@134100.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 74:20:@134094.4]
  assign regs_30_clock = clock; // @[:@134103.4]
  assign regs_30_reset = io_reset; // @[:@134104.4 RegFile.scala 76:16:@134111.4]
  assign regs_30_io_in = 64'h0; // @[RegFile.scala 75:16:@134110.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@134114.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 74:20:@134108.4]
  assign regs_31_clock = clock; // @[:@134117.4]
  assign regs_31_reset = io_reset; // @[:@134118.4 RegFile.scala 76:16:@134125.4]
  assign regs_31_io_in = 64'h0; // @[RegFile.scala 75:16:@134124.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@134128.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 74:20:@134122.4]
  assign regs_32_clock = clock; // @[:@134131.4]
  assign regs_32_reset = io_reset; // @[:@134132.4 RegFile.scala 76:16:@134139.4]
  assign regs_32_io_in = 64'h0; // @[RegFile.scala 75:16:@134138.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@134142.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 74:20:@134136.4]
  assign regs_33_clock = clock; // @[:@134145.4]
  assign regs_33_reset = io_reset; // @[:@134146.4 RegFile.scala 76:16:@134153.4]
  assign regs_33_io_in = 64'h0; // @[RegFile.scala 75:16:@134152.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@134156.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 74:20:@134150.4]
  assign regs_34_clock = clock; // @[:@134159.4]
  assign regs_34_reset = io_reset; // @[:@134160.4 RegFile.scala 76:16:@134167.4]
  assign regs_34_io_in = 64'h0; // @[RegFile.scala 75:16:@134166.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@134170.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 74:20:@134164.4]
  assign regs_35_clock = clock; // @[:@134173.4]
  assign regs_35_reset = io_reset; // @[:@134174.4 RegFile.scala 76:16:@134181.4]
  assign regs_35_io_in = 64'h0; // @[RegFile.scala 75:16:@134180.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@134184.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@134178.4]
  assign regs_36_clock = clock; // @[:@134187.4]
  assign regs_36_reset = io_reset; // @[:@134188.4 RegFile.scala 76:16:@134195.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 75:16:@134194.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@134198.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@134192.4]
  assign regs_37_clock = clock; // @[:@134201.4]
  assign regs_37_reset = io_reset; // @[:@134202.4 RegFile.scala 76:16:@134209.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 75:16:@134208.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@134212.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@134206.4]
  assign regs_38_clock = clock; // @[:@134215.4]
  assign regs_38_reset = io_reset; // @[:@134216.4 RegFile.scala 76:16:@134223.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 75:16:@134222.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@134226.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@134220.4]
  assign regs_39_clock = clock; // @[:@134229.4]
  assign regs_39_reset = io_reset; // @[:@134230.4 RegFile.scala 76:16:@134237.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 75:16:@134236.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@134240.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@134234.4]
  assign regs_40_clock = clock; // @[:@134243.4]
  assign regs_40_reset = io_reset; // @[:@134244.4 RegFile.scala 76:16:@134251.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 75:16:@134250.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@134254.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@134248.4]
  assign regs_41_clock = clock; // @[:@134257.4]
  assign regs_41_reset = io_reset; // @[:@134258.4 RegFile.scala 76:16:@134265.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 75:16:@134264.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@134268.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@134262.4]
  assign regs_42_clock = clock; // @[:@134271.4]
  assign regs_42_reset = io_reset; // @[:@134272.4 RegFile.scala 76:16:@134279.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 75:16:@134278.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@134282.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@134276.4]
  assign regs_43_clock = clock; // @[:@134285.4]
  assign regs_43_reset = io_reset; // @[:@134286.4 RegFile.scala 76:16:@134293.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 75:16:@134292.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@134296.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@134290.4]
  assign regs_44_clock = clock; // @[:@134299.4]
  assign regs_44_reset = io_reset; // @[:@134300.4 RegFile.scala 76:16:@134307.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 75:16:@134306.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@134310.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@134304.4]
  assign regs_45_clock = clock; // @[:@134313.4]
  assign regs_45_reset = io_reset; // @[:@134314.4 RegFile.scala 76:16:@134321.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 75:16:@134320.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@134324.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@134318.4]
  assign regs_46_clock = clock; // @[:@134327.4]
  assign regs_46_reset = io_reset; // @[:@134328.4 RegFile.scala 76:16:@134335.4]
  assign regs_46_io_in = 64'h0; // @[RegFile.scala 75:16:@134334.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@134338.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@134332.4]
  assign regs_47_clock = clock; // @[:@134341.4]
  assign regs_47_reset = io_reset; // @[:@134342.4 RegFile.scala 76:16:@134349.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 75:16:@134348.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@134352.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@134346.4]
  assign regs_48_clock = clock; // @[:@134355.4]
  assign regs_48_reset = io_reset; // @[:@134356.4 RegFile.scala 76:16:@134363.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 75:16:@134362.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@134366.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@134360.4]
  assign regs_49_clock = clock; // @[:@134369.4]
  assign regs_49_reset = io_reset; // @[:@134370.4 RegFile.scala 76:16:@134377.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@134376.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@134380.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@134374.4]
  assign regs_50_clock = clock; // @[:@134383.4]
  assign regs_50_reset = io_reset; // @[:@134384.4 RegFile.scala 76:16:@134391.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@134390.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@134394.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@134388.4]
  assign regs_51_clock = clock; // @[:@134397.4]
  assign regs_51_reset = io_reset; // @[:@134398.4 RegFile.scala 76:16:@134405.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@134404.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@134408.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@134402.4]
  assign regs_52_clock = clock; // @[:@134411.4]
  assign regs_52_reset = io_reset; // @[:@134412.4 RegFile.scala 76:16:@134419.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@134418.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@134422.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@134416.4]
  assign regs_53_clock = clock; // @[:@134425.4]
  assign regs_53_reset = io_reset; // @[:@134426.4 RegFile.scala 76:16:@134433.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@134432.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@134436.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@134430.4]
  assign regs_54_clock = clock; // @[:@134439.4]
  assign regs_54_reset = io_reset; // @[:@134440.4 RegFile.scala 76:16:@134447.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@134446.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@134450.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@134444.4]
  assign regs_55_clock = clock; // @[:@134453.4]
  assign regs_55_reset = io_reset; // @[:@134454.4 RegFile.scala 76:16:@134461.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@134460.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@134464.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@134458.4]
  assign regs_56_clock = clock; // @[:@134467.4]
  assign regs_56_reset = io_reset; // @[:@134468.4 RegFile.scala 76:16:@134475.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@134474.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@134478.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@134472.4]
  assign regs_57_clock = clock; // @[:@134481.4]
  assign regs_57_reset = io_reset; // @[:@134482.4 RegFile.scala 76:16:@134489.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@134488.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@134492.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@134486.4]
  assign regs_58_clock = clock; // @[:@134495.4]
  assign regs_58_reset = io_reset; // @[:@134496.4 RegFile.scala 76:16:@134503.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@134502.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@134506.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@134500.4]
  assign regs_59_clock = clock; // @[:@134509.4]
  assign regs_59_reset = io_reset; // @[:@134510.4 RegFile.scala 76:16:@134517.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 75:16:@134516.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@134520.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@134514.4]
  assign regs_60_clock = clock; // @[:@134523.4]
  assign regs_60_reset = io_reset; // @[:@134524.4 RegFile.scala 76:16:@134531.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@134530.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@134534.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@134528.4]
  assign regs_61_clock = clock; // @[:@134537.4]
  assign regs_61_reset = io_reset; // @[:@134538.4 RegFile.scala 76:16:@134545.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@134544.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@134548.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@134542.4]
  assign regs_62_clock = clock; // @[:@134551.4]
  assign regs_62_reset = io_reset; // @[:@134552.4 RegFile.scala 76:16:@134559.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@134558.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@134562.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@134556.4]
  assign regs_63_clock = clock; // @[:@134565.4]
  assign regs_63_reset = io_reset; // @[:@134566.4 RegFile.scala 76:16:@134573.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@134572.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@134576.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@134570.4]
  assign regs_64_clock = clock; // @[:@134579.4]
  assign regs_64_reset = io_reset; // @[:@134580.4 RegFile.scala 76:16:@134587.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@134586.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@134590.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@134584.4]
  assign regs_65_clock = clock; // @[:@134593.4]
  assign regs_65_reset = io_reset; // @[:@134594.4 RegFile.scala 76:16:@134601.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@134600.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@134604.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@134598.4]
  assign regs_66_clock = clock; // @[:@134607.4]
  assign regs_66_reset = io_reset; // @[:@134608.4 RegFile.scala 76:16:@134615.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@134614.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@134618.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@134612.4]
  assign regs_67_clock = clock; // @[:@134621.4]
  assign regs_67_reset = io_reset; // @[:@134622.4 RegFile.scala 76:16:@134629.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@134628.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@134632.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@134626.4]
  assign regs_68_clock = clock; // @[:@134635.4]
  assign regs_68_reset = io_reset; // @[:@134636.4 RegFile.scala 76:16:@134643.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@134642.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@134646.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@134640.4]
  assign regs_69_clock = clock; // @[:@134649.4]
  assign regs_69_reset = io_reset; // @[:@134650.4 RegFile.scala 76:16:@134657.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@134656.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@134660.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@134654.4]
  assign regs_70_clock = clock; // @[:@134663.4]
  assign regs_70_reset = io_reset; // @[:@134664.4 RegFile.scala 76:16:@134671.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@134670.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@134674.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@134668.4]
  assign regs_71_clock = clock; // @[:@134677.4]
  assign regs_71_reset = io_reset; // @[:@134678.4 RegFile.scala 76:16:@134685.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@134684.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@134688.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@134682.4]
  assign regs_72_clock = clock; // @[:@134691.4]
  assign regs_72_reset = io_reset; // @[:@134692.4 RegFile.scala 76:16:@134699.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@134698.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@134702.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@134696.4]
  assign regs_73_clock = clock; // @[:@134705.4]
  assign regs_73_reset = io_reset; // @[:@134706.4 RegFile.scala 76:16:@134713.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@134712.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@134716.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@134710.4]
  assign regs_74_clock = clock; // @[:@134719.4]
  assign regs_74_reset = io_reset; // @[:@134720.4 RegFile.scala 76:16:@134727.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@134726.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@134730.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@134724.4]
  assign regs_75_clock = clock; // @[:@134733.4]
  assign regs_75_reset = io_reset; // @[:@134734.4 RegFile.scala 76:16:@134741.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@134740.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@134744.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@134738.4]
  assign regs_76_clock = clock; // @[:@134747.4]
  assign regs_76_reset = io_reset; // @[:@134748.4 RegFile.scala 76:16:@134755.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@134754.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@134758.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@134752.4]
  assign regs_77_clock = clock; // @[:@134761.4]
  assign regs_77_reset = io_reset; // @[:@134762.4 RegFile.scala 76:16:@134769.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@134768.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@134772.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@134766.4]
  assign regs_78_clock = clock; // @[:@134775.4]
  assign regs_78_reset = io_reset; // @[:@134776.4 RegFile.scala 76:16:@134783.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@134782.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@134786.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@134780.4]
  assign regs_79_clock = clock; // @[:@134789.4]
  assign regs_79_reset = io_reset; // @[:@134790.4 RegFile.scala 76:16:@134797.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@134796.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@134800.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@134794.4]
  assign regs_80_clock = clock; // @[:@134803.4]
  assign regs_80_reset = io_reset; // @[:@134804.4 RegFile.scala 76:16:@134811.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@134810.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@134814.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@134808.4]
  assign regs_81_clock = clock; // @[:@134817.4]
  assign regs_81_reset = io_reset; // @[:@134818.4 RegFile.scala 76:16:@134825.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@134824.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@134828.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@134822.4]
  assign regs_82_clock = clock; // @[:@134831.4]
  assign regs_82_reset = io_reset; // @[:@134832.4 RegFile.scala 76:16:@134839.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@134838.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@134842.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@134836.4]
  assign regs_83_clock = clock; // @[:@134845.4]
  assign regs_83_reset = io_reset; // @[:@134846.4 RegFile.scala 76:16:@134853.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@134852.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@134856.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@134850.4]
  assign regs_84_clock = clock; // @[:@134859.4]
  assign regs_84_reset = io_reset; // @[:@134860.4 RegFile.scala 76:16:@134867.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@134866.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@134870.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@134864.4]
  assign regs_85_clock = clock; // @[:@134873.4]
  assign regs_85_reset = io_reset; // @[:@134874.4 RegFile.scala 76:16:@134881.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@134880.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@134884.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@134878.4]
  assign regs_86_clock = clock; // @[:@134887.4]
  assign regs_86_reset = io_reset; // @[:@134888.4 RegFile.scala 76:16:@134895.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@134894.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@134898.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@134892.4]
  assign regs_87_clock = clock; // @[:@134901.4]
  assign regs_87_reset = io_reset; // @[:@134902.4 RegFile.scala 76:16:@134909.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@134908.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@134912.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@134906.4]
  assign regs_88_clock = clock; // @[:@134915.4]
  assign regs_88_reset = io_reset; // @[:@134916.4 RegFile.scala 76:16:@134923.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@134922.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@134926.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@134920.4]
  assign regs_89_clock = clock; // @[:@134929.4]
  assign regs_89_reset = io_reset; // @[:@134930.4 RegFile.scala 76:16:@134937.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@134936.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@134940.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@134934.4]
  assign regs_90_clock = clock; // @[:@134943.4]
  assign regs_90_reset = io_reset; // @[:@134944.4 RegFile.scala 76:16:@134951.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@134950.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@134954.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@134948.4]
  assign regs_91_clock = clock; // @[:@134957.4]
  assign regs_91_reset = io_reset; // @[:@134958.4 RegFile.scala 76:16:@134965.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@134964.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@134968.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@134962.4]
  assign regs_92_clock = clock; // @[:@134971.4]
  assign regs_92_reset = io_reset; // @[:@134972.4 RegFile.scala 76:16:@134979.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@134978.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@134982.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@134976.4]
  assign regs_93_clock = clock; // @[:@134985.4]
  assign regs_93_reset = io_reset; // @[:@134986.4 RegFile.scala 76:16:@134993.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@134992.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@134996.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@134990.4]
  assign regs_94_clock = clock; // @[:@134999.4]
  assign regs_94_reset = io_reset; // @[:@135000.4 RegFile.scala 76:16:@135007.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@135006.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@135010.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@135004.4]
  assign regs_95_clock = clock; // @[:@135013.4]
  assign regs_95_reset = io_reset; // @[:@135014.4 RegFile.scala 76:16:@135021.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@135020.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@135024.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@135018.4]
  assign regs_96_clock = clock; // @[:@135027.4]
  assign regs_96_reset = io_reset; // @[:@135028.4 RegFile.scala 76:16:@135035.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@135034.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@135038.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@135032.4]
  assign regs_97_clock = clock; // @[:@135041.4]
  assign regs_97_reset = io_reset; // @[:@135042.4 RegFile.scala 76:16:@135049.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@135048.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@135052.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@135046.4]
  assign regs_98_clock = clock; // @[:@135055.4]
  assign regs_98_reset = io_reset; // @[:@135056.4 RegFile.scala 76:16:@135063.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@135062.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@135066.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@135060.4]
  assign regs_99_clock = clock; // @[:@135069.4]
  assign regs_99_reset = io_reset; // @[:@135070.4 RegFile.scala 76:16:@135077.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@135076.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@135080.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@135074.4]
  assign regs_100_clock = clock; // @[:@135083.4]
  assign regs_100_reset = io_reset; // @[:@135084.4 RegFile.scala 76:16:@135091.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@135090.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@135094.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@135088.4]
  assign regs_101_clock = clock; // @[:@135097.4]
  assign regs_101_reset = io_reset; // @[:@135098.4 RegFile.scala 76:16:@135105.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@135104.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@135108.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@135102.4]
  assign regs_102_clock = clock; // @[:@135111.4]
  assign regs_102_reset = io_reset; // @[:@135112.4 RegFile.scala 76:16:@135119.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@135118.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@135122.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@135116.4]
  assign regs_103_clock = clock; // @[:@135125.4]
  assign regs_103_reset = io_reset; // @[:@135126.4 RegFile.scala 76:16:@135133.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@135132.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@135136.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@135130.4]
  assign regs_104_clock = clock; // @[:@135139.4]
  assign regs_104_reset = io_reset; // @[:@135140.4 RegFile.scala 76:16:@135147.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@135146.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@135150.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@135144.4]
  assign regs_105_clock = clock; // @[:@135153.4]
  assign regs_105_reset = io_reset; // @[:@135154.4 RegFile.scala 76:16:@135161.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@135160.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@135164.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@135158.4]
  assign regs_106_clock = clock; // @[:@135167.4]
  assign regs_106_reset = io_reset; // @[:@135168.4 RegFile.scala 76:16:@135175.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@135174.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@135178.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@135172.4]
  assign regs_107_clock = clock; // @[:@135181.4]
  assign regs_107_reset = io_reset; // @[:@135182.4 RegFile.scala 76:16:@135189.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@135188.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@135192.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@135186.4]
  assign regs_108_clock = clock; // @[:@135195.4]
  assign regs_108_reset = io_reset; // @[:@135196.4 RegFile.scala 76:16:@135203.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@135202.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@135206.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@135200.4]
  assign regs_109_clock = clock; // @[:@135209.4]
  assign regs_109_reset = io_reset; // @[:@135210.4 RegFile.scala 76:16:@135217.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@135216.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@135220.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@135214.4]
  assign regs_110_clock = clock; // @[:@135223.4]
  assign regs_110_reset = io_reset; // @[:@135224.4 RegFile.scala 76:16:@135231.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@135230.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@135234.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@135228.4]
  assign regs_111_clock = clock; // @[:@135237.4]
  assign regs_111_reset = io_reset; // @[:@135238.4 RegFile.scala 76:16:@135245.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@135244.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@135248.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@135242.4]
  assign regs_112_clock = clock; // @[:@135251.4]
  assign regs_112_reset = io_reset; // @[:@135252.4 RegFile.scala 76:16:@135259.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@135258.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@135262.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@135256.4]
  assign regs_113_clock = clock; // @[:@135265.4]
  assign regs_113_reset = io_reset; // @[:@135266.4 RegFile.scala 76:16:@135273.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@135272.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@135276.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@135270.4]
  assign regs_114_clock = clock; // @[:@135279.4]
  assign regs_114_reset = io_reset; // @[:@135280.4 RegFile.scala 76:16:@135287.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@135286.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@135290.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@135284.4]
  assign regs_115_clock = clock; // @[:@135293.4]
  assign regs_115_reset = io_reset; // @[:@135294.4 RegFile.scala 76:16:@135301.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@135300.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@135304.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@135298.4]
  assign regs_116_clock = clock; // @[:@135307.4]
  assign regs_116_reset = io_reset; // @[:@135308.4 RegFile.scala 76:16:@135315.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@135314.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@135318.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@135312.4]
  assign regs_117_clock = clock; // @[:@135321.4]
  assign regs_117_reset = io_reset; // @[:@135322.4 RegFile.scala 76:16:@135329.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@135328.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@135332.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@135326.4]
  assign regs_118_clock = clock; // @[:@135335.4]
  assign regs_118_reset = io_reset; // @[:@135336.4 RegFile.scala 76:16:@135343.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@135342.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@135346.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@135340.4]
  assign regs_119_clock = clock; // @[:@135349.4]
  assign regs_119_reset = io_reset; // @[:@135350.4 RegFile.scala 76:16:@135357.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@135356.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@135360.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@135354.4]
  assign regs_120_clock = clock; // @[:@135363.4]
  assign regs_120_reset = io_reset; // @[:@135364.4 RegFile.scala 76:16:@135371.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@135370.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@135374.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@135368.4]
  assign regs_121_clock = clock; // @[:@135377.4]
  assign regs_121_reset = io_reset; // @[:@135378.4 RegFile.scala 76:16:@135385.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@135384.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@135388.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@135382.4]
  assign regs_122_clock = clock; // @[:@135391.4]
  assign regs_122_reset = io_reset; // @[:@135392.4 RegFile.scala 76:16:@135399.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@135398.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@135402.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@135396.4]
  assign regs_123_clock = clock; // @[:@135405.4]
  assign regs_123_reset = io_reset; // @[:@135406.4 RegFile.scala 76:16:@135413.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@135412.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@135416.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@135410.4]
  assign regs_124_clock = clock; // @[:@135419.4]
  assign regs_124_reset = io_reset; // @[:@135420.4 RegFile.scala 76:16:@135427.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@135426.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@135430.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@135424.4]
  assign regs_125_clock = clock; // @[:@135433.4]
  assign regs_125_reset = io_reset; // @[:@135434.4 RegFile.scala 76:16:@135441.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@135440.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@135444.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@135438.4]
  assign regs_126_clock = clock; // @[:@135447.4]
  assign regs_126_reset = io_reset; // @[:@135448.4 RegFile.scala 76:16:@135455.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@135454.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@135458.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@135452.4]
  assign regs_127_clock = clock; // @[:@135461.4]
  assign regs_127_reset = io_reset; // @[:@135462.4 RegFile.scala 76:16:@135469.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@135468.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@135472.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@135466.4]
  assign regs_128_clock = clock; // @[:@135475.4]
  assign regs_128_reset = io_reset; // @[:@135476.4 RegFile.scala 76:16:@135483.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@135482.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@135486.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@135480.4]
  assign regs_129_clock = clock; // @[:@135489.4]
  assign regs_129_reset = io_reset; // @[:@135490.4 RegFile.scala 76:16:@135497.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@135496.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@135500.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@135494.4]
  assign regs_130_clock = clock; // @[:@135503.4]
  assign regs_130_reset = io_reset; // @[:@135504.4 RegFile.scala 76:16:@135511.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@135510.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@135514.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@135508.4]
  assign regs_131_clock = clock; // @[:@135517.4]
  assign regs_131_reset = io_reset; // @[:@135518.4 RegFile.scala 76:16:@135525.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@135524.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@135528.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@135522.4]
  assign regs_132_clock = clock; // @[:@135531.4]
  assign regs_132_reset = io_reset; // @[:@135532.4 RegFile.scala 76:16:@135539.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@135538.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@135542.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@135536.4]
  assign regs_133_clock = clock; // @[:@135545.4]
  assign regs_133_reset = io_reset; // @[:@135546.4 RegFile.scala 76:16:@135553.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@135552.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@135556.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@135550.4]
  assign regs_134_clock = clock; // @[:@135559.4]
  assign regs_134_reset = io_reset; // @[:@135560.4 RegFile.scala 76:16:@135567.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@135566.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@135570.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@135564.4]
  assign regs_135_clock = clock; // @[:@135573.4]
  assign regs_135_reset = io_reset; // @[:@135574.4 RegFile.scala 76:16:@135581.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@135580.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@135584.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@135578.4]
  assign regs_136_clock = clock; // @[:@135587.4]
  assign regs_136_reset = io_reset; // @[:@135588.4 RegFile.scala 76:16:@135595.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@135594.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@135598.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@135592.4]
  assign regs_137_clock = clock; // @[:@135601.4]
  assign regs_137_reset = io_reset; // @[:@135602.4 RegFile.scala 76:16:@135609.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@135608.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@135612.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@135606.4]
  assign regs_138_clock = clock; // @[:@135615.4]
  assign regs_138_reset = io_reset; // @[:@135616.4 RegFile.scala 76:16:@135623.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@135622.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@135626.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@135620.4]
  assign regs_139_clock = clock; // @[:@135629.4]
  assign regs_139_reset = io_reset; // @[:@135630.4 RegFile.scala 76:16:@135637.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@135636.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@135640.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@135634.4]
  assign regs_140_clock = clock; // @[:@135643.4]
  assign regs_140_reset = io_reset; // @[:@135644.4 RegFile.scala 76:16:@135651.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@135650.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@135654.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@135648.4]
  assign regs_141_clock = clock; // @[:@135657.4]
  assign regs_141_reset = io_reset; // @[:@135658.4 RegFile.scala 76:16:@135665.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@135664.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@135668.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@135662.4]
  assign regs_142_clock = clock; // @[:@135671.4]
  assign regs_142_reset = io_reset; // @[:@135672.4 RegFile.scala 76:16:@135679.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@135678.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@135682.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@135676.4]
  assign regs_143_clock = clock; // @[:@135685.4]
  assign regs_143_reset = io_reset; // @[:@135686.4 RegFile.scala 76:16:@135693.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@135692.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@135696.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@135690.4]
  assign regs_144_clock = clock; // @[:@135699.4]
  assign regs_144_reset = io_reset; // @[:@135700.4 RegFile.scala 76:16:@135707.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@135706.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@135710.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@135704.4]
  assign regs_145_clock = clock; // @[:@135713.4]
  assign regs_145_reset = io_reset; // @[:@135714.4 RegFile.scala 76:16:@135721.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@135720.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@135724.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@135718.4]
  assign regs_146_clock = clock; // @[:@135727.4]
  assign regs_146_reset = io_reset; // @[:@135728.4 RegFile.scala 76:16:@135735.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@135734.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@135738.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@135732.4]
  assign regs_147_clock = clock; // @[:@135741.4]
  assign regs_147_reset = io_reset; // @[:@135742.4 RegFile.scala 76:16:@135749.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@135748.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@135752.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@135746.4]
  assign regs_148_clock = clock; // @[:@135755.4]
  assign regs_148_reset = io_reset; // @[:@135756.4 RegFile.scala 76:16:@135763.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@135762.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@135766.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@135760.4]
  assign regs_149_clock = clock; // @[:@135769.4]
  assign regs_149_reset = io_reset; // @[:@135770.4 RegFile.scala 76:16:@135777.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@135776.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@135780.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@135774.4]
  assign regs_150_clock = clock; // @[:@135783.4]
  assign regs_150_reset = io_reset; // @[:@135784.4 RegFile.scala 76:16:@135791.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@135790.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@135794.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@135788.4]
  assign regs_151_clock = clock; // @[:@135797.4]
  assign regs_151_reset = io_reset; // @[:@135798.4 RegFile.scala 76:16:@135805.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@135804.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@135808.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@135802.4]
  assign regs_152_clock = clock; // @[:@135811.4]
  assign regs_152_reset = io_reset; // @[:@135812.4 RegFile.scala 76:16:@135819.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@135818.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@135822.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@135816.4]
  assign regs_153_clock = clock; // @[:@135825.4]
  assign regs_153_reset = io_reset; // @[:@135826.4 RegFile.scala 76:16:@135833.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@135832.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@135836.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@135830.4]
  assign regs_154_clock = clock; // @[:@135839.4]
  assign regs_154_reset = io_reset; // @[:@135840.4 RegFile.scala 76:16:@135847.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@135846.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@135850.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@135844.4]
  assign regs_155_clock = clock; // @[:@135853.4]
  assign regs_155_reset = io_reset; // @[:@135854.4 RegFile.scala 76:16:@135861.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@135860.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@135864.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@135858.4]
  assign regs_156_clock = clock; // @[:@135867.4]
  assign regs_156_reset = io_reset; // @[:@135868.4 RegFile.scala 76:16:@135875.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@135874.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@135878.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@135872.4]
  assign regs_157_clock = clock; // @[:@135881.4]
  assign regs_157_reset = io_reset; // @[:@135882.4 RegFile.scala 76:16:@135889.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@135888.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@135892.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@135886.4]
  assign regs_158_clock = clock; // @[:@135895.4]
  assign regs_158_reset = io_reset; // @[:@135896.4 RegFile.scala 76:16:@135903.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@135902.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@135906.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@135900.4]
  assign regs_159_clock = clock; // @[:@135909.4]
  assign regs_159_reset = io_reset; // @[:@135910.4 RegFile.scala 76:16:@135917.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@135916.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@135920.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@135914.4]
  assign regs_160_clock = clock; // @[:@135923.4]
  assign regs_160_reset = io_reset; // @[:@135924.4 RegFile.scala 76:16:@135931.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@135930.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@135934.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@135928.4]
  assign regs_161_clock = clock; // @[:@135937.4]
  assign regs_161_reset = io_reset; // @[:@135938.4 RegFile.scala 76:16:@135945.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@135944.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@135948.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@135942.4]
  assign regs_162_clock = clock; // @[:@135951.4]
  assign regs_162_reset = io_reset; // @[:@135952.4 RegFile.scala 76:16:@135959.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@135958.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@135962.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@135956.4]
  assign regs_163_clock = clock; // @[:@135965.4]
  assign regs_163_reset = io_reset; // @[:@135966.4 RegFile.scala 76:16:@135973.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@135972.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@135976.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@135970.4]
  assign regs_164_clock = clock; // @[:@135979.4]
  assign regs_164_reset = io_reset; // @[:@135980.4 RegFile.scala 76:16:@135987.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@135986.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@135990.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@135984.4]
  assign regs_165_clock = clock; // @[:@135993.4]
  assign regs_165_reset = io_reset; // @[:@135994.4 RegFile.scala 76:16:@136001.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@136000.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@136004.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@135998.4]
  assign regs_166_clock = clock; // @[:@136007.4]
  assign regs_166_reset = io_reset; // @[:@136008.4 RegFile.scala 76:16:@136015.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@136014.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@136018.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@136012.4]
  assign regs_167_clock = clock; // @[:@136021.4]
  assign regs_167_reset = io_reset; // @[:@136022.4 RegFile.scala 76:16:@136029.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@136028.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@136032.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@136026.4]
  assign regs_168_clock = clock; // @[:@136035.4]
  assign regs_168_reset = io_reset; // @[:@136036.4 RegFile.scala 76:16:@136043.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@136042.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@136046.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@136040.4]
  assign regs_169_clock = clock; // @[:@136049.4]
  assign regs_169_reset = io_reset; // @[:@136050.4 RegFile.scala 76:16:@136057.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@136056.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@136060.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@136054.4]
  assign regs_170_clock = clock; // @[:@136063.4]
  assign regs_170_reset = io_reset; // @[:@136064.4 RegFile.scala 76:16:@136071.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@136070.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@136074.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@136068.4]
  assign regs_171_clock = clock; // @[:@136077.4]
  assign regs_171_reset = io_reset; // @[:@136078.4 RegFile.scala 76:16:@136085.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@136084.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@136088.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@136082.4]
  assign regs_172_clock = clock; // @[:@136091.4]
  assign regs_172_reset = io_reset; // @[:@136092.4 RegFile.scala 76:16:@136099.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@136098.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@136102.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@136096.4]
  assign regs_173_clock = clock; // @[:@136105.4]
  assign regs_173_reset = io_reset; // @[:@136106.4 RegFile.scala 76:16:@136113.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@136112.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@136116.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@136110.4]
  assign regs_174_clock = clock; // @[:@136119.4]
  assign regs_174_reset = io_reset; // @[:@136120.4 RegFile.scala 76:16:@136127.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@136126.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@136130.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@136124.4]
  assign regs_175_clock = clock; // @[:@136133.4]
  assign regs_175_reset = io_reset; // @[:@136134.4 RegFile.scala 76:16:@136141.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@136140.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@136144.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@136138.4]
  assign regs_176_clock = clock; // @[:@136147.4]
  assign regs_176_reset = io_reset; // @[:@136148.4 RegFile.scala 76:16:@136155.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@136154.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@136158.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@136152.4]
  assign regs_177_clock = clock; // @[:@136161.4]
  assign regs_177_reset = io_reset; // @[:@136162.4 RegFile.scala 76:16:@136169.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@136168.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@136172.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@136166.4]
  assign regs_178_clock = clock; // @[:@136175.4]
  assign regs_178_reset = io_reset; // @[:@136176.4 RegFile.scala 76:16:@136183.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@136182.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@136186.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@136180.4]
  assign regs_179_clock = clock; // @[:@136189.4]
  assign regs_179_reset = io_reset; // @[:@136190.4 RegFile.scala 76:16:@136197.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@136196.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@136200.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@136194.4]
  assign regs_180_clock = clock; // @[:@136203.4]
  assign regs_180_reset = io_reset; // @[:@136204.4 RegFile.scala 76:16:@136211.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@136210.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@136214.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@136208.4]
  assign regs_181_clock = clock; // @[:@136217.4]
  assign regs_181_reset = io_reset; // @[:@136218.4 RegFile.scala 76:16:@136225.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@136224.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@136228.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@136222.4]
  assign regs_182_clock = clock; // @[:@136231.4]
  assign regs_182_reset = io_reset; // @[:@136232.4 RegFile.scala 76:16:@136239.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@136238.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@136242.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@136236.4]
  assign regs_183_clock = clock; // @[:@136245.4]
  assign regs_183_reset = io_reset; // @[:@136246.4 RegFile.scala 76:16:@136253.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@136252.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@136256.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@136250.4]
  assign regs_184_clock = clock; // @[:@136259.4]
  assign regs_184_reset = io_reset; // @[:@136260.4 RegFile.scala 76:16:@136267.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@136266.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@136270.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@136264.4]
  assign regs_185_clock = clock; // @[:@136273.4]
  assign regs_185_reset = io_reset; // @[:@136274.4 RegFile.scala 76:16:@136281.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@136280.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@136284.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@136278.4]
  assign regs_186_clock = clock; // @[:@136287.4]
  assign regs_186_reset = io_reset; // @[:@136288.4 RegFile.scala 76:16:@136295.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@136294.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@136298.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@136292.4]
  assign regs_187_clock = clock; // @[:@136301.4]
  assign regs_187_reset = io_reset; // @[:@136302.4 RegFile.scala 76:16:@136309.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@136308.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@136312.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@136306.4]
  assign regs_188_clock = clock; // @[:@136315.4]
  assign regs_188_reset = io_reset; // @[:@136316.4 RegFile.scala 76:16:@136323.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@136322.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@136326.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@136320.4]
  assign regs_189_clock = clock; // @[:@136329.4]
  assign regs_189_reset = io_reset; // @[:@136330.4 RegFile.scala 76:16:@136337.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@136336.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@136340.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@136334.4]
  assign regs_190_clock = clock; // @[:@136343.4]
  assign regs_190_reset = io_reset; // @[:@136344.4 RegFile.scala 76:16:@136351.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@136350.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@136354.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@136348.4]
  assign regs_191_clock = clock; // @[:@136357.4]
  assign regs_191_reset = io_reset; // @[:@136358.4 RegFile.scala 76:16:@136365.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@136364.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@136368.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@136362.4]
  assign regs_192_clock = clock; // @[:@136371.4]
  assign regs_192_reset = io_reset; // @[:@136372.4 RegFile.scala 76:16:@136379.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@136378.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@136382.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@136376.4]
  assign regs_193_clock = clock; // @[:@136385.4]
  assign regs_193_reset = io_reset; // @[:@136386.4 RegFile.scala 76:16:@136393.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@136392.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@136396.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@136390.4]
  assign regs_194_clock = clock; // @[:@136399.4]
  assign regs_194_reset = io_reset; // @[:@136400.4 RegFile.scala 76:16:@136407.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@136406.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@136410.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@136404.4]
  assign regs_195_clock = clock; // @[:@136413.4]
  assign regs_195_reset = io_reset; // @[:@136414.4 RegFile.scala 76:16:@136421.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@136420.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@136424.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@136418.4]
  assign regs_196_clock = clock; // @[:@136427.4]
  assign regs_196_reset = io_reset; // @[:@136428.4 RegFile.scala 76:16:@136435.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@136434.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@136438.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@136432.4]
  assign regs_197_clock = clock; // @[:@136441.4]
  assign regs_197_reset = io_reset; // @[:@136442.4 RegFile.scala 76:16:@136449.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@136448.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@136452.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@136446.4]
  assign regs_198_clock = clock; // @[:@136455.4]
  assign regs_198_reset = io_reset; // @[:@136456.4 RegFile.scala 76:16:@136463.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@136462.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@136466.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@136460.4]
  assign regs_199_clock = clock; // @[:@136469.4]
  assign regs_199_reset = io_reset; // @[:@136470.4 RegFile.scala 76:16:@136477.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@136476.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@136480.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@136474.4]
  assign regs_200_clock = clock; // @[:@136483.4]
  assign regs_200_reset = io_reset; // @[:@136484.4 RegFile.scala 76:16:@136491.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@136490.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@136494.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@136488.4]
  assign regs_201_clock = clock; // @[:@136497.4]
  assign regs_201_reset = io_reset; // @[:@136498.4 RegFile.scala 76:16:@136505.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@136504.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@136508.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@136502.4]
  assign regs_202_clock = clock; // @[:@136511.4]
  assign regs_202_reset = io_reset; // @[:@136512.4 RegFile.scala 76:16:@136519.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@136518.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@136522.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@136516.4]
  assign regs_203_clock = clock; // @[:@136525.4]
  assign regs_203_reset = io_reset; // @[:@136526.4 RegFile.scala 76:16:@136533.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@136532.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@136536.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@136530.4]
  assign regs_204_clock = clock; // @[:@136539.4]
  assign regs_204_reset = io_reset; // @[:@136540.4 RegFile.scala 76:16:@136547.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@136546.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@136550.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@136544.4]
  assign regs_205_clock = clock; // @[:@136553.4]
  assign regs_205_reset = io_reset; // @[:@136554.4 RegFile.scala 76:16:@136561.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@136560.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@136564.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@136558.4]
  assign regs_206_clock = clock; // @[:@136567.4]
  assign regs_206_reset = io_reset; // @[:@136568.4 RegFile.scala 76:16:@136575.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@136574.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@136578.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@136572.4]
  assign regs_207_clock = clock; // @[:@136581.4]
  assign regs_207_reset = io_reset; // @[:@136582.4 RegFile.scala 76:16:@136589.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@136588.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@136592.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@136586.4]
  assign regs_208_clock = clock; // @[:@136595.4]
  assign regs_208_reset = io_reset; // @[:@136596.4 RegFile.scala 76:16:@136603.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@136602.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@136606.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@136600.4]
  assign regs_209_clock = clock; // @[:@136609.4]
  assign regs_209_reset = io_reset; // @[:@136610.4 RegFile.scala 76:16:@136617.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@136616.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@136620.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@136614.4]
  assign regs_210_clock = clock; // @[:@136623.4]
  assign regs_210_reset = io_reset; // @[:@136624.4 RegFile.scala 76:16:@136631.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@136630.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@136634.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@136628.4]
  assign regs_211_clock = clock; // @[:@136637.4]
  assign regs_211_reset = io_reset; // @[:@136638.4 RegFile.scala 76:16:@136645.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@136644.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@136648.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@136642.4]
  assign regs_212_clock = clock; // @[:@136651.4]
  assign regs_212_reset = io_reset; // @[:@136652.4 RegFile.scala 76:16:@136659.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@136658.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@136662.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@136656.4]
  assign regs_213_clock = clock; // @[:@136665.4]
  assign regs_213_reset = io_reset; // @[:@136666.4 RegFile.scala 76:16:@136673.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@136672.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@136676.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@136670.4]
  assign regs_214_clock = clock; // @[:@136679.4]
  assign regs_214_reset = io_reset; // @[:@136680.4 RegFile.scala 76:16:@136687.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@136686.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@136690.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@136684.4]
  assign regs_215_clock = clock; // @[:@136693.4]
  assign regs_215_reset = io_reset; // @[:@136694.4 RegFile.scala 76:16:@136701.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@136700.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@136704.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@136698.4]
  assign regs_216_clock = clock; // @[:@136707.4]
  assign regs_216_reset = io_reset; // @[:@136708.4 RegFile.scala 76:16:@136715.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@136714.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@136718.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@136712.4]
  assign regs_217_clock = clock; // @[:@136721.4]
  assign regs_217_reset = io_reset; // @[:@136722.4 RegFile.scala 76:16:@136729.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@136728.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@136732.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@136726.4]
  assign regs_218_clock = clock; // @[:@136735.4]
  assign regs_218_reset = io_reset; // @[:@136736.4 RegFile.scala 76:16:@136743.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@136742.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@136746.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@136740.4]
  assign regs_219_clock = clock; // @[:@136749.4]
  assign regs_219_reset = io_reset; // @[:@136750.4 RegFile.scala 76:16:@136757.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@136756.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@136760.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@136754.4]
  assign regs_220_clock = clock; // @[:@136763.4]
  assign regs_220_reset = io_reset; // @[:@136764.4 RegFile.scala 76:16:@136771.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@136770.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@136774.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@136768.4]
  assign regs_221_clock = clock; // @[:@136777.4]
  assign regs_221_reset = io_reset; // @[:@136778.4 RegFile.scala 76:16:@136785.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@136784.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@136788.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@136782.4]
  assign regs_222_clock = clock; // @[:@136791.4]
  assign regs_222_reset = io_reset; // @[:@136792.4 RegFile.scala 76:16:@136799.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@136798.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@136802.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@136796.4]
  assign regs_223_clock = clock; // @[:@136805.4]
  assign regs_223_reset = io_reset; // @[:@136806.4 RegFile.scala 76:16:@136813.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@136812.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@136816.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@136810.4]
  assign regs_224_clock = clock; // @[:@136819.4]
  assign regs_224_reset = io_reset; // @[:@136820.4 RegFile.scala 76:16:@136827.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@136826.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@136830.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@136824.4]
  assign regs_225_clock = clock; // @[:@136833.4]
  assign regs_225_reset = io_reset; // @[:@136834.4 RegFile.scala 76:16:@136841.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@136840.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@136844.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@136838.4]
  assign regs_226_clock = clock; // @[:@136847.4]
  assign regs_226_reset = io_reset; // @[:@136848.4 RegFile.scala 76:16:@136855.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@136854.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@136858.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@136852.4]
  assign regs_227_clock = clock; // @[:@136861.4]
  assign regs_227_reset = io_reset; // @[:@136862.4 RegFile.scala 76:16:@136869.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@136868.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@136872.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@136866.4]
  assign regs_228_clock = clock; // @[:@136875.4]
  assign regs_228_reset = io_reset; // @[:@136876.4 RegFile.scala 76:16:@136883.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@136882.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@136886.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@136880.4]
  assign regs_229_clock = clock; // @[:@136889.4]
  assign regs_229_reset = io_reset; // @[:@136890.4 RegFile.scala 76:16:@136897.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@136896.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@136900.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@136894.4]
  assign regs_230_clock = clock; // @[:@136903.4]
  assign regs_230_reset = io_reset; // @[:@136904.4 RegFile.scala 76:16:@136911.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@136910.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@136914.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@136908.4]
  assign regs_231_clock = clock; // @[:@136917.4]
  assign regs_231_reset = io_reset; // @[:@136918.4 RegFile.scala 76:16:@136925.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@136924.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@136928.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@136922.4]
  assign regs_232_clock = clock; // @[:@136931.4]
  assign regs_232_reset = io_reset; // @[:@136932.4 RegFile.scala 76:16:@136939.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@136938.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@136942.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@136936.4]
  assign regs_233_clock = clock; // @[:@136945.4]
  assign regs_233_reset = io_reset; // @[:@136946.4 RegFile.scala 76:16:@136953.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@136952.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@136956.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@136950.4]
  assign regs_234_clock = clock; // @[:@136959.4]
  assign regs_234_reset = io_reset; // @[:@136960.4 RegFile.scala 76:16:@136967.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@136966.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@136970.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@136964.4]
  assign regs_235_clock = clock; // @[:@136973.4]
  assign regs_235_reset = io_reset; // @[:@136974.4 RegFile.scala 76:16:@136981.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@136980.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@136984.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@136978.4]
  assign regs_236_clock = clock; // @[:@136987.4]
  assign regs_236_reset = io_reset; // @[:@136988.4 RegFile.scala 76:16:@136995.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@136994.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@136998.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@136992.4]
  assign regs_237_clock = clock; // @[:@137001.4]
  assign regs_237_reset = io_reset; // @[:@137002.4 RegFile.scala 76:16:@137009.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@137008.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@137012.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@137006.4]
  assign regs_238_clock = clock; // @[:@137015.4]
  assign regs_238_reset = io_reset; // @[:@137016.4 RegFile.scala 76:16:@137023.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@137022.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@137026.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@137020.4]
  assign regs_239_clock = clock; // @[:@137029.4]
  assign regs_239_reset = io_reset; // @[:@137030.4 RegFile.scala 76:16:@137037.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@137036.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@137040.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@137034.4]
  assign regs_240_clock = clock; // @[:@137043.4]
  assign regs_240_reset = io_reset; // @[:@137044.4 RegFile.scala 76:16:@137051.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@137050.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@137054.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@137048.4]
  assign regs_241_clock = clock; // @[:@137057.4]
  assign regs_241_reset = io_reset; // @[:@137058.4 RegFile.scala 76:16:@137065.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@137064.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@137068.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@137062.4]
  assign regs_242_clock = clock; // @[:@137071.4]
  assign regs_242_reset = io_reset; // @[:@137072.4 RegFile.scala 76:16:@137079.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@137078.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@137082.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@137076.4]
  assign regs_243_clock = clock; // @[:@137085.4]
  assign regs_243_reset = io_reset; // @[:@137086.4 RegFile.scala 76:16:@137093.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@137092.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@137096.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@137090.4]
  assign regs_244_clock = clock; // @[:@137099.4]
  assign regs_244_reset = io_reset; // @[:@137100.4 RegFile.scala 76:16:@137107.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@137106.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@137110.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@137104.4]
  assign regs_245_clock = clock; // @[:@137113.4]
  assign regs_245_reset = io_reset; // @[:@137114.4 RegFile.scala 76:16:@137121.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@137120.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@137124.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@137118.4]
  assign regs_246_clock = clock; // @[:@137127.4]
  assign regs_246_reset = io_reset; // @[:@137128.4 RegFile.scala 76:16:@137135.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@137134.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@137138.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@137132.4]
  assign regs_247_clock = clock; // @[:@137141.4]
  assign regs_247_reset = io_reset; // @[:@137142.4 RegFile.scala 76:16:@137149.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@137148.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@137152.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@137146.4]
  assign regs_248_clock = clock; // @[:@137155.4]
  assign regs_248_reset = io_reset; // @[:@137156.4 RegFile.scala 76:16:@137163.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@137162.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@137166.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@137160.4]
  assign regs_249_clock = clock; // @[:@137169.4]
  assign regs_249_reset = io_reset; // @[:@137170.4 RegFile.scala 76:16:@137177.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@137176.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@137180.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@137174.4]
  assign regs_250_clock = clock; // @[:@137183.4]
  assign regs_250_reset = io_reset; // @[:@137184.4 RegFile.scala 76:16:@137191.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@137190.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@137194.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@137188.4]
  assign regs_251_clock = clock; // @[:@137197.4]
  assign regs_251_reset = io_reset; // @[:@137198.4 RegFile.scala 76:16:@137205.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@137204.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@137208.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@137202.4]
  assign regs_252_clock = clock; // @[:@137211.4]
  assign regs_252_reset = io_reset; // @[:@137212.4 RegFile.scala 76:16:@137219.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@137218.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@137222.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@137216.4]
  assign regs_253_clock = clock; // @[:@137225.4]
  assign regs_253_reset = io_reset; // @[:@137226.4 RegFile.scala 76:16:@137233.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@137232.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@137236.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@137230.4]
  assign regs_254_clock = clock; // @[:@137239.4]
  assign regs_254_reset = io_reset; // @[:@137240.4 RegFile.scala 76:16:@137247.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@137246.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@137250.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@137244.4]
  assign regs_255_clock = clock; // @[:@137253.4]
  assign regs_255_reset = io_reset; // @[:@137254.4 RegFile.scala 76:16:@137261.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@137260.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@137264.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@137258.4]
  assign regs_256_clock = clock; // @[:@137267.4]
  assign regs_256_reset = io_reset; // @[:@137268.4 RegFile.scala 76:16:@137275.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@137274.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@137278.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@137272.4]
  assign regs_257_clock = clock; // @[:@137281.4]
  assign regs_257_reset = io_reset; // @[:@137282.4 RegFile.scala 76:16:@137289.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@137288.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@137292.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@137286.4]
  assign regs_258_clock = clock; // @[:@137295.4]
  assign regs_258_reset = io_reset; // @[:@137296.4 RegFile.scala 76:16:@137303.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@137302.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@137306.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@137300.4]
  assign regs_259_clock = clock; // @[:@137309.4]
  assign regs_259_reset = io_reset; // @[:@137310.4 RegFile.scala 76:16:@137317.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@137316.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@137320.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@137314.4]
  assign regs_260_clock = clock; // @[:@137323.4]
  assign regs_260_reset = io_reset; // @[:@137324.4 RegFile.scala 76:16:@137331.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@137330.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@137334.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@137328.4]
  assign regs_261_clock = clock; // @[:@137337.4]
  assign regs_261_reset = io_reset; // @[:@137338.4 RegFile.scala 76:16:@137345.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@137344.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@137348.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@137342.4]
  assign regs_262_clock = clock; // @[:@137351.4]
  assign regs_262_reset = io_reset; // @[:@137352.4 RegFile.scala 76:16:@137359.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@137358.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@137362.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@137356.4]
  assign regs_263_clock = clock; // @[:@137365.4]
  assign regs_263_reset = io_reset; // @[:@137366.4 RegFile.scala 76:16:@137373.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@137372.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@137376.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@137370.4]
  assign regs_264_clock = clock; // @[:@137379.4]
  assign regs_264_reset = io_reset; // @[:@137380.4 RegFile.scala 76:16:@137387.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@137386.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@137390.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@137384.4]
  assign regs_265_clock = clock; // @[:@137393.4]
  assign regs_265_reset = io_reset; // @[:@137394.4 RegFile.scala 76:16:@137401.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@137400.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@137404.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@137398.4]
  assign regs_266_clock = clock; // @[:@137407.4]
  assign regs_266_reset = io_reset; // @[:@137408.4 RegFile.scala 76:16:@137415.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@137414.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@137418.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@137412.4]
  assign regs_267_clock = clock; // @[:@137421.4]
  assign regs_267_reset = io_reset; // @[:@137422.4 RegFile.scala 76:16:@137429.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@137428.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@137432.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@137426.4]
  assign regs_268_clock = clock; // @[:@137435.4]
  assign regs_268_reset = io_reset; // @[:@137436.4 RegFile.scala 76:16:@137443.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@137442.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@137446.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@137440.4]
  assign regs_269_clock = clock; // @[:@137449.4]
  assign regs_269_reset = io_reset; // @[:@137450.4 RegFile.scala 76:16:@137457.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@137456.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@137460.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@137454.4]
  assign regs_270_clock = clock; // @[:@137463.4]
  assign regs_270_reset = io_reset; // @[:@137464.4 RegFile.scala 76:16:@137471.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@137470.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@137474.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@137468.4]
  assign regs_271_clock = clock; // @[:@137477.4]
  assign regs_271_reset = io_reset; // @[:@137478.4 RegFile.scala 76:16:@137485.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@137484.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@137488.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@137482.4]
  assign regs_272_clock = clock; // @[:@137491.4]
  assign regs_272_reset = io_reset; // @[:@137492.4 RegFile.scala 76:16:@137499.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@137498.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@137502.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@137496.4]
  assign regs_273_clock = clock; // @[:@137505.4]
  assign regs_273_reset = io_reset; // @[:@137506.4 RegFile.scala 76:16:@137513.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@137512.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@137516.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@137510.4]
  assign regs_274_clock = clock; // @[:@137519.4]
  assign regs_274_reset = io_reset; // @[:@137520.4 RegFile.scala 76:16:@137527.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@137526.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@137530.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@137524.4]
  assign regs_275_clock = clock; // @[:@137533.4]
  assign regs_275_reset = io_reset; // @[:@137534.4 RegFile.scala 76:16:@137541.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@137540.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@137544.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@137538.4]
  assign regs_276_clock = clock; // @[:@137547.4]
  assign regs_276_reset = io_reset; // @[:@137548.4 RegFile.scala 76:16:@137555.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@137554.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@137558.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@137552.4]
  assign regs_277_clock = clock; // @[:@137561.4]
  assign regs_277_reset = io_reset; // @[:@137562.4 RegFile.scala 76:16:@137569.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@137568.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@137572.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@137566.4]
  assign regs_278_clock = clock; // @[:@137575.4]
  assign regs_278_reset = io_reset; // @[:@137576.4 RegFile.scala 76:16:@137583.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@137582.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@137586.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@137580.4]
  assign regs_279_clock = clock; // @[:@137589.4]
  assign regs_279_reset = io_reset; // @[:@137590.4 RegFile.scala 76:16:@137597.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@137596.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@137600.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@137594.4]
  assign regs_280_clock = clock; // @[:@137603.4]
  assign regs_280_reset = io_reset; // @[:@137604.4 RegFile.scala 76:16:@137611.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@137610.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@137614.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@137608.4]
  assign regs_281_clock = clock; // @[:@137617.4]
  assign regs_281_reset = io_reset; // @[:@137618.4 RegFile.scala 76:16:@137625.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@137624.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@137628.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@137622.4]
  assign regs_282_clock = clock; // @[:@137631.4]
  assign regs_282_reset = io_reset; // @[:@137632.4 RegFile.scala 76:16:@137639.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@137638.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@137642.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@137636.4]
  assign regs_283_clock = clock; // @[:@137645.4]
  assign regs_283_reset = io_reset; // @[:@137646.4 RegFile.scala 76:16:@137653.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@137652.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@137656.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@137650.4]
  assign regs_284_clock = clock; // @[:@137659.4]
  assign regs_284_reset = io_reset; // @[:@137660.4 RegFile.scala 76:16:@137667.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@137666.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@137670.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@137664.4]
  assign regs_285_clock = clock; // @[:@137673.4]
  assign regs_285_reset = io_reset; // @[:@137674.4 RegFile.scala 76:16:@137681.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@137680.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@137684.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@137678.4]
  assign regs_286_clock = clock; // @[:@137687.4]
  assign regs_286_reset = io_reset; // @[:@137688.4 RegFile.scala 76:16:@137695.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@137694.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@137698.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@137692.4]
  assign regs_287_clock = clock; // @[:@137701.4]
  assign regs_287_reset = io_reset; // @[:@137702.4 RegFile.scala 76:16:@137709.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@137708.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@137712.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@137706.4]
  assign regs_288_clock = clock; // @[:@137715.4]
  assign regs_288_reset = io_reset; // @[:@137716.4 RegFile.scala 76:16:@137723.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@137722.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@137726.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@137720.4]
  assign regs_289_clock = clock; // @[:@137729.4]
  assign regs_289_reset = io_reset; // @[:@137730.4 RegFile.scala 76:16:@137737.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@137736.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@137740.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@137734.4]
  assign regs_290_clock = clock; // @[:@137743.4]
  assign regs_290_reset = io_reset; // @[:@137744.4 RegFile.scala 76:16:@137751.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@137750.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@137754.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@137748.4]
  assign regs_291_clock = clock; // @[:@137757.4]
  assign regs_291_reset = io_reset; // @[:@137758.4 RegFile.scala 76:16:@137765.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@137764.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@137768.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@137762.4]
  assign regs_292_clock = clock; // @[:@137771.4]
  assign regs_292_reset = io_reset; // @[:@137772.4 RegFile.scala 76:16:@137779.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@137778.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@137782.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@137776.4]
  assign regs_293_clock = clock; // @[:@137785.4]
  assign regs_293_reset = io_reset; // @[:@137786.4 RegFile.scala 76:16:@137793.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@137792.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@137796.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@137790.4]
  assign regs_294_clock = clock; // @[:@137799.4]
  assign regs_294_reset = io_reset; // @[:@137800.4 RegFile.scala 76:16:@137807.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@137806.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@137810.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@137804.4]
  assign regs_295_clock = clock; // @[:@137813.4]
  assign regs_295_reset = io_reset; // @[:@137814.4 RegFile.scala 76:16:@137821.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@137820.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@137824.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@137818.4]
  assign regs_296_clock = clock; // @[:@137827.4]
  assign regs_296_reset = io_reset; // @[:@137828.4 RegFile.scala 76:16:@137835.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@137834.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@137838.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@137832.4]
  assign regs_297_clock = clock; // @[:@137841.4]
  assign regs_297_reset = io_reset; // @[:@137842.4 RegFile.scala 76:16:@137849.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@137848.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@137852.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@137846.4]
  assign regs_298_clock = clock; // @[:@137855.4]
  assign regs_298_reset = io_reset; // @[:@137856.4 RegFile.scala 76:16:@137863.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@137862.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@137866.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@137860.4]
  assign regs_299_clock = clock; // @[:@137869.4]
  assign regs_299_reset = io_reset; // @[:@137870.4 RegFile.scala 76:16:@137877.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@137876.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@137880.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@137874.4]
  assign regs_300_clock = clock; // @[:@137883.4]
  assign regs_300_reset = io_reset; // @[:@137884.4 RegFile.scala 76:16:@137891.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@137890.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@137894.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@137888.4]
  assign regs_301_clock = clock; // @[:@137897.4]
  assign regs_301_reset = io_reset; // @[:@137898.4 RegFile.scala 76:16:@137905.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@137904.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@137908.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@137902.4]
  assign regs_302_clock = clock; // @[:@137911.4]
  assign regs_302_reset = io_reset; // @[:@137912.4 RegFile.scala 76:16:@137919.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@137918.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@137922.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@137916.4]
  assign regs_303_clock = clock; // @[:@137925.4]
  assign regs_303_reset = io_reset; // @[:@137926.4 RegFile.scala 76:16:@137933.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@137932.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@137936.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@137930.4]
  assign regs_304_clock = clock; // @[:@137939.4]
  assign regs_304_reset = io_reset; // @[:@137940.4 RegFile.scala 76:16:@137947.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@137946.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@137950.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@137944.4]
  assign regs_305_clock = clock; // @[:@137953.4]
  assign regs_305_reset = io_reset; // @[:@137954.4 RegFile.scala 76:16:@137961.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@137960.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@137964.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@137958.4]
  assign regs_306_clock = clock; // @[:@137967.4]
  assign regs_306_reset = io_reset; // @[:@137968.4 RegFile.scala 76:16:@137975.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@137974.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@137978.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@137972.4]
  assign regs_307_clock = clock; // @[:@137981.4]
  assign regs_307_reset = io_reset; // @[:@137982.4 RegFile.scala 76:16:@137989.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@137988.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@137992.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@137986.4]
  assign regs_308_clock = clock; // @[:@137995.4]
  assign regs_308_reset = io_reset; // @[:@137996.4 RegFile.scala 76:16:@138003.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@138002.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@138006.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@138000.4]
  assign regs_309_clock = clock; // @[:@138009.4]
  assign regs_309_reset = io_reset; // @[:@138010.4 RegFile.scala 76:16:@138017.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@138016.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@138020.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@138014.4]
  assign regs_310_clock = clock; // @[:@138023.4]
  assign regs_310_reset = io_reset; // @[:@138024.4 RegFile.scala 76:16:@138031.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@138030.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@138034.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@138028.4]
  assign regs_311_clock = clock; // @[:@138037.4]
  assign regs_311_reset = io_reset; // @[:@138038.4 RegFile.scala 76:16:@138045.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@138044.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@138048.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@138042.4]
  assign regs_312_clock = clock; // @[:@138051.4]
  assign regs_312_reset = io_reset; // @[:@138052.4 RegFile.scala 76:16:@138059.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@138058.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@138062.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@138056.4]
  assign regs_313_clock = clock; // @[:@138065.4]
  assign regs_313_reset = io_reset; // @[:@138066.4 RegFile.scala 76:16:@138073.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@138072.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@138076.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@138070.4]
  assign regs_314_clock = clock; // @[:@138079.4]
  assign regs_314_reset = io_reset; // @[:@138080.4 RegFile.scala 76:16:@138087.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@138086.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@138090.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@138084.4]
  assign regs_315_clock = clock; // @[:@138093.4]
  assign regs_315_reset = io_reset; // @[:@138094.4 RegFile.scala 76:16:@138101.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@138100.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@138104.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@138098.4]
  assign regs_316_clock = clock; // @[:@138107.4]
  assign regs_316_reset = io_reset; // @[:@138108.4 RegFile.scala 76:16:@138115.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@138114.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@138118.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@138112.4]
  assign regs_317_clock = clock; // @[:@138121.4]
  assign regs_317_reset = io_reset; // @[:@138122.4 RegFile.scala 76:16:@138129.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@138128.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@138132.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@138126.4]
  assign regs_318_clock = clock; // @[:@138135.4]
  assign regs_318_reset = io_reset; // @[:@138136.4 RegFile.scala 76:16:@138143.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@138142.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@138146.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@138140.4]
  assign regs_319_clock = clock; // @[:@138149.4]
  assign regs_319_reset = io_reset; // @[:@138150.4 RegFile.scala 76:16:@138157.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@138156.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@138160.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@138154.4]
  assign regs_320_clock = clock; // @[:@138163.4]
  assign regs_320_reset = io_reset; // @[:@138164.4 RegFile.scala 76:16:@138171.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@138170.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@138174.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@138168.4]
  assign regs_321_clock = clock; // @[:@138177.4]
  assign regs_321_reset = io_reset; // @[:@138178.4 RegFile.scala 76:16:@138185.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@138184.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@138188.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@138182.4]
  assign regs_322_clock = clock; // @[:@138191.4]
  assign regs_322_reset = io_reset; // @[:@138192.4 RegFile.scala 76:16:@138199.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@138198.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@138202.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@138196.4]
  assign regs_323_clock = clock; // @[:@138205.4]
  assign regs_323_reset = io_reset; // @[:@138206.4 RegFile.scala 76:16:@138213.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@138212.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@138216.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@138210.4]
  assign regs_324_clock = clock; // @[:@138219.4]
  assign regs_324_reset = io_reset; // @[:@138220.4 RegFile.scala 76:16:@138227.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@138226.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@138230.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@138224.4]
  assign regs_325_clock = clock; // @[:@138233.4]
  assign regs_325_reset = io_reset; // @[:@138234.4 RegFile.scala 76:16:@138241.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@138240.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@138244.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@138238.4]
  assign regs_326_clock = clock; // @[:@138247.4]
  assign regs_326_reset = io_reset; // @[:@138248.4 RegFile.scala 76:16:@138255.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@138254.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@138258.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@138252.4]
  assign regs_327_clock = clock; // @[:@138261.4]
  assign regs_327_reset = io_reset; // @[:@138262.4 RegFile.scala 76:16:@138269.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@138268.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@138272.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@138266.4]
  assign regs_328_clock = clock; // @[:@138275.4]
  assign regs_328_reset = io_reset; // @[:@138276.4 RegFile.scala 76:16:@138283.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@138282.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@138286.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@138280.4]
  assign regs_329_clock = clock; // @[:@138289.4]
  assign regs_329_reset = io_reset; // @[:@138290.4 RegFile.scala 76:16:@138297.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@138296.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@138300.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@138294.4]
  assign regs_330_clock = clock; // @[:@138303.4]
  assign regs_330_reset = io_reset; // @[:@138304.4 RegFile.scala 76:16:@138311.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@138310.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@138314.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@138308.4]
  assign regs_331_clock = clock; // @[:@138317.4]
  assign regs_331_reset = io_reset; // @[:@138318.4 RegFile.scala 76:16:@138325.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@138324.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@138328.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@138322.4]
  assign regs_332_clock = clock; // @[:@138331.4]
  assign regs_332_reset = io_reset; // @[:@138332.4 RegFile.scala 76:16:@138339.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@138338.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@138342.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@138336.4]
  assign regs_333_clock = clock; // @[:@138345.4]
  assign regs_333_reset = io_reset; // @[:@138346.4 RegFile.scala 76:16:@138353.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@138352.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@138356.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@138350.4]
  assign regs_334_clock = clock; // @[:@138359.4]
  assign regs_334_reset = io_reset; // @[:@138360.4 RegFile.scala 76:16:@138367.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@138366.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@138370.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@138364.4]
  assign regs_335_clock = clock; // @[:@138373.4]
  assign regs_335_reset = io_reset; // @[:@138374.4 RegFile.scala 76:16:@138381.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@138380.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@138384.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@138378.4]
  assign regs_336_clock = clock; // @[:@138387.4]
  assign regs_336_reset = io_reset; // @[:@138388.4 RegFile.scala 76:16:@138395.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@138394.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@138398.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@138392.4]
  assign regs_337_clock = clock; // @[:@138401.4]
  assign regs_337_reset = io_reset; // @[:@138402.4 RegFile.scala 76:16:@138409.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@138408.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@138412.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@138406.4]
  assign regs_338_clock = clock; // @[:@138415.4]
  assign regs_338_reset = io_reset; // @[:@138416.4 RegFile.scala 76:16:@138423.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@138422.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@138426.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@138420.4]
  assign regs_339_clock = clock; // @[:@138429.4]
  assign regs_339_reset = io_reset; // @[:@138430.4 RegFile.scala 76:16:@138437.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@138436.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@138440.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@138434.4]
  assign regs_340_clock = clock; // @[:@138443.4]
  assign regs_340_reset = io_reset; // @[:@138444.4 RegFile.scala 76:16:@138451.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@138450.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@138454.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@138448.4]
  assign regs_341_clock = clock; // @[:@138457.4]
  assign regs_341_reset = io_reset; // @[:@138458.4 RegFile.scala 76:16:@138465.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@138464.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@138468.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@138462.4]
  assign regs_342_clock = clock; // @[:@138471.4]
  assign regs_342_reset = io_reset; // @[:@138472.4 RegFile.scala 76:16:@138479.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@138478.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@138482.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@138476.4]
  assign regs_343_clock = clock; // @[:@138485.4]
  assign regs_343_reset = io_reset; // @[:@138486.4 RegFile.scala 76:16:@138493.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@138492.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@138496.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@138490.4]
  assign regs_344_clock = clock; // @[:@138499.4]
  assign regs_344_reset = io_reset; // @[:@138500.4 RegFile.scala 76:16:@138507.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@138506.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@138510.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@138504.4]
  assign regs_345_clock = clock; // @[:@138513.4]
  assign regs_345_reset = io_reset; // @[:@138514.4 RegFile.scala 76:16:@138521.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@138520.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@138524.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@138518.4]
  assign regs_346_clock = clock; // @[:@138527.4]
  assign regs_346_reset = io_reset; // @[:@138528.4 RegFile.scala 76:16:@138535.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@138534.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@138538.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@138532.4]
  assign regs_347_clock = clock; // @[:@138541.4]
  assign regs_347_reset = io_reset; // @[:@138542.4 RegFile.scala 76:16:@138549.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@138548.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@138552.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@138546.4]
  assign regs_348_clock = clock; // @[:@138555.4]
  assign regs_348_reset = io_reset; // @[:@138556.4 RegFile.scala 76:16:@138563.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@138562.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@138566.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@138560.4]
  assign regs_349_clock = clock; // @[:@138569.4]
  assign regs_349_reset = io_reset; // @[:@138570.4 RegFile.scala 76:16:@138577.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@138576.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@138580.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@138574.4]
  assign regs_350_clock = clock; // @[:@138583.4]
  assign regs_350_reset = io_reset; // @[:@138584.4 RegFile.scala 76:16:@138591.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@138590.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@138594.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@138588.4]
  assign regs_351_clock = clock; // @[:@138597.4]
  assign regs_351_reset = io_reset; // @[:@138598.4 RegFile.scala 76:16:@138605.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@138604.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@138608.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@138602.4]
  assign regs_352_clock = clock; // @[:@138611.4]
  assign regs_352_reset = io_reset; // @[:@138612.4 RegFile.scala 76:16:@138619.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@138618.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@138622.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@138616.4]
  assign regs_353_clock = clock; // @[:@138625.4]
  assign regs_353_reset = io_reset; // @[:@138626.4 RegFile.scala 76:16:@138633.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@138632.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@138636.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@138630.4]
  assign regs_354_clock = clock; // @[:@138639.4]
  assign regs_354_reset = io_reset; // @[:@138640.4 RegFile.scala 76:16:@138647.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@138646.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@138650.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@138644.4]
  assign regs_355_clock = clock; // @[:@138653.4]
  assign regs_355_reset = io_reset; // @[:@138654.4 RegFile.scala 76:16:@138661.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@138660.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@138664.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@138658.4]
  assign regs_356_clock = clock; // @[:@138667.4]
  assign regs_356_reset = io_reset; // @[:@138668.4 RegFile.scala 76:16:@138675.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@138674.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@138678.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@138672.4]
  assign regs_357_clock = clock; // @[:@138681.4]
  assign regs_357_reset = io_reset; // @[:@138682.4 RegFile.scala 76:16:@138689.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@138688.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@138692.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@138686.4]
  assign regs_358_clock = clock; // @[:@138695.4]
  assign regs_358_reset = io_reset; // @[:@138696.4 RegFile.scala 76:16:@138703.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@138702.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@138706.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@138700.4]
  assign regs_359_clock = clock; // @[:@138709.4]
  assign regs_359_reset = io_reset; // @[:@138710.4 RegFile.scala 76:16:@138717.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@138716.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@138720.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@138714.4]
  assign regs_360_clock = clock; // @[:@138723.4]
  assign regs_360_reset = io_reset; // @[:@138724.4 RegFile.scala 76:16:@138731.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@138730.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@138734.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@138728.4]
  assign regs_361_clock = clock; // @[:@138737.4]
  assign regs_361_reset = io_reset; // @[:@138738.4 RegFile.scala 76:16:@138745.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@138744.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@138748.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@138742.4]
  assign regs_362_clock = clock; // @[:@138751.4]
  assign regs_362_reset = io_reset; // @[:@138752.4 RegFile.scala 76:16:@138759.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@138758.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@138762.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@138756.4]
  assign regs_363_clock = clock; // @[:@138765.4]
  assign regs_363_reset = io_reset; // @[:@138766.4 RegFile.scala 76:16:@138773.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@138772.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@138776.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@138770.4]
  assign regs_364_clock = clock; // @[:@138779.4]
  assign regs_364_reset = io_reset; // @[:@138780.4 RegFile.scala 76:16:@138787.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@138786.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@138790.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@138784.4]
  assign regs_365_clock = clock; // @[:@138793.4]
  assign regs_365_reset = io_reset; // @[:@138794.4 RegFile.scala 76:16:@138801.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@138800.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@138804.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@138798.4]
  assign regs_366_clock = clock; // @[:@138807.4]
  assign regs_366_reset = io_reset; // @[:@138808.4 RegFile.scala 76:16:@138815.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@138814.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@138818.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@138812.4]
  assign regs_367_clock = clock; // @[:@138821.4]
  assign regs_367_reset = io_reset; // @[:@138822.4 RegFile.scala 76:16:@138829.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@138828.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@138832.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@138826.4]
  assign regs_368_clock = clock; // @[:@138835.4]
  assign regs_368_reset = io_reset; // @[:@138836.4 RegFile.scala 76:16:@138843.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@138842.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@138846.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@138840.4]
  assign regs_369_clock = clock; // @[:@138849.4]
  assign regs_369_reset = io_reset; // @[:@138850.4 RegFile.scala 76:16:@138857.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@138856.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@138860.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@138854.4]
  assign regs_370_clock = clock; // @[:@138863.4]
  assign regs_370_reset = io_reset; // @[:@138864.4 RegFile.scala 76:16:@138871.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@138870.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@138874.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@138868.4]
  assign regs_371_clock = clock; // @[:@138877.4]
  assign regs_371_reset = io_reset; // @[:@138878.4 RegFile.scala 76:16:@138885.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@138884.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@138888.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@138882.4]
  assign regs_372_clock = clock; // @[:@138891.4]
  assign regs_372_reset = io_reset; // @[:@138892.4 RegFile.scala 76:16:@138899.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@138898.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@138902.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@138896.4]
  assign regs_373_clock = clock; // @[:@138905.4]
  assign regs_373_reset = io_reset; // @[:@138906.4 RegFile.scala 76:16:@138913.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@138912.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@138916.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@138910.4]
  assign regs_374_clock = clock; // @[:@138919.4]
  assign regs_374_reset = io_reset; // @[:@138920.4 RegFile.scala 76:16:@138927.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@138926.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@138930.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@138924.4]
  assign regs_375_clock = clock; // @[:@138933.4]
  assign regs_375_reset = io_reset; // @[:@138934.4 RegFile.scala 76:16:@138941.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@138940.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@138944.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@138938.4]
  assign regs_376_clock = clock; // @[:@138947.4]
  assign regs_376_reset = io_reset; // @[:@138948.4 RegFile.scala 76:16:@138955.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@138954.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@138958.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@138952.4]
  assign regs_377_clock = clock; // @[:@138961.4]
  assign regs_377_reset = io_reset; // @[:@138962.4 RegFile.scala 76:16:@138969.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@138968.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@138972.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@138966.4]
  assign regs_378_clock = clock; // @[:@138975.4]
  assign regs_378_reset = io_reset; // @[:@138976.4 RegFile.scala 76:16:@138983.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@138982.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@138986.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@138980.4]
  assign regs_379_clock = clock; // @[:@138989.4]
  assign regs_379_reset = io_reset; // @[:@138990.4 RegFile.scala 76:16:@138997.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@138996.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@139000.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@138994.4]
  assign regs_380_clock = clock; // @[:@139003.4]
  assign regs_380_reset = io_reset; // @[:@139004.4 RegFile.scala 76:16:@139011.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@139010.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@139014.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@139008.4]
  assign regs_381_clock = clock; // @[:@139017.4]
  assign regs_381_reset = io_reset; // @[:@139018.4 RegFile.scala 76:16:@139025.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@139024.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@139028.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@139022.4]
  assign regs_382_clock = clock; // @[:@139031.4]
  assign regs_382_reset = io_reset; // @[:@139032.4 RegFile.scala 76:16:@139039.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@139038.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@139042.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@139036.4]
  assign regs_383_clock = clock; // @[:@139045.4]
  assign regs_383_reset = io_reset; // @[:@139046.4 RegFile.scala 76:16:@139053.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@139052.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@139056.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@139050.4]
  assign regs_384_clock = clock; // @[:@139059.4]
  assign regs_384_reset = io_reset; // @[:@139060.4 RegFile.scala 76:16:@139067.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@139066.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@139070.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@139064.4]
  assign regs_385_clock = clock; // @[:@139073.4]
  assign regs_385_reset = io_reset; // @[:@139074.4 RegFile.scala 76:16:@139081.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@139080.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@139084.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@139078.4]
  assign regs_386_clock = clock; // @[:@139087.4]
  assign regs_386_reset = io_reset; // @[:@139088.4 RegFile.scala 76:16:@139095.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@139094.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@139098.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@139092.4]
  assign regs_387_clock = clock; // @[:@139101.4]
  assign regs_387_reset = io_reset; // @[:@139102.4 RegFile.scala 76:16:@139109.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@139108.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@139112.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@139106.4]
  assign regs_388_clock = clock; // @[:@139115.4]
  assign regs_388_reset = io_reset; // @[:@139116.4 RegFile.scala 76:16:@139123.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@139122.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@139126.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@139120.4]
  assign regs_389_clock = clock; // @[:@139129.4]
  assign regs_389_reset = io_reset; // @[:@139130.4 RegFile.scala 76:16:@139137.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@139136.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@139140.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@139134.4]
  assign regs_390_clock = clock; // @[:@139143.4]
  assign regs_390_reset = io_reset; // @[:@139144.4 RegFile.scala 76:16:@139151.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@139150.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@139154.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@139148.4]
  assign regs_391_clock = clock; // @[:@139157.4]
  assign regs_391_reset = io_reset; // @[:@139158.4 RegFile.scala 76:16:@139165.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@139164.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@139168.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@139162.4]
  assign regs_392_clock = clock; // @[:@139171.4]
  assign regs_392_reset = io_reset; // @[:@139172.4 RegFile.scala 76:16:@139179.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@139178.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@139182.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@139176.4]
  assign regs_393_clock = clock; // @[:@139185.4]
  assign regs_393_reset = io_reset; // @[:@139186.4 RegFile.scala 76:16:@139193.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@139192.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@139196.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@139190.4]
  assign regs_394_clock = clock; // @[:@139199.4]
  assign regs_394_reset = io_reset; // @[:@139200.4 RegFile.scala 76:16:@139207.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@139206.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@139210.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@139204.4]
  assign regs_395_clock = clock; // @[:@139213.4]
  assign regs_395_reset = io_reset; // @[:@139214.4 RegFile.scala 76:16:@139221.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@139220.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@139224.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@139218.4]
  assign regs_396_clock = clock; // @[:@139227.4]
  assign regs_396_reset = io_reset; // @[:@139228.4 RegFile.scala 76:16:@139235.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@139234.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@139238.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@139232.4]
  assign regs_397_clock = clock; // @[:@139241.4]
  assign regs_397_reset = io_reset; // @[:@139242.4 RegFile.scala 76:16:@139249.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@139248.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@139252.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@139246.4]
  assign regs_398_clock = clock; // @[:@139255.4]
  assign regs_398_reset = io_reset; // @[:@139256.4 RegFile.scala 76:16:@139263.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@139262.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@139266.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@139260.4]
  assign regs_399_clock = clock; // @[:@139269.4]
  assign regs_399_reset = io_reset; // @[:@139270.4 RegFile.scala 76:16:@139277.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@139276.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@139280.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@139274.4]
  assign regs_400_clock = clock; // @[:@139283.4]
  assign regs_400_reset = io_reset; // @[:@139284.4 RegFile.scala 76:16:@139291.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@139290.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@139294.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@139288.4]
  assign regs_401_clock = clock; // @[:@139297.4]
  assign regs_401_reset = io_reset; // @[:@139298.4 RegFile.scala 76:16:@139305.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@139304.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@139308.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@139302.4]
  assign regs_402_clock = clock; // @[:@139311.4]
  assign regs_402_reset = io_reset; // @[:@139312.4 RegFile.scala 76:16:@139319.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@139318.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@139322.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@139316.4]
  assign regs_403_clock = clock; // @[:@139325.4]
  assign regs_403_reset = io_reset; // @[:@139326.4 RegFile.scala 76:16:@139333.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@139332.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@139336.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@139330.4]
  assign regs_404_clock = clock; // @[:@139339.4]
  assign regs_404_reset = io_reset; // @[:@139340.4 RegFile.scala 76:16:@139347.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@139346.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@139350.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@139344.4]
  assign regs_405_clock = clock; // @[:@139353.4]
  assign regs_405_reset = io_reset; // @[:@139354.4 RegFile.scala 76:16:@139361.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@139360.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@139364.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@139358.4]
  assign regs_406_clock = clock; // @[:@139367.4]
  assign regs_406_reset = io_reset; // @[:@139368.4 RegFile.scala 76:16:@139375.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@139374.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@139378.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@139372.4]
  assign regs_407_clock = clock; // @[:@139381.4]
  assign regs_407_reset = io_reset; // @[:@139382.4 RegFile.scala 76:16:@139389.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@139388.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@139392.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@139386.4]
  assign regs_408_clock = clock; // @[:@139395.4]
  assign regs_408_reset = io_reset; // @[:@139396.4 RegFile.scala 76:16:@139403.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@139402.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@139406.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@139400.4]
  assign regs_409_clock = clock; // @[:@139409.4]
  assign regs_409_reset = io_reset; // @[:@139410.4 RegFile.scala 76:16:@139417.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@139416.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@139420.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@139414.4]
  assign regs_410_clock = clock; // @[:@139423.4]
  assign regs_410_reset = io_reset; // @[:@139424.4 RegFile.scala 76:16:@139431.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@139430.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@139434.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@139428.4]
  assign regs_411_clock = clock; // @[:@139437.4]
  assign regs_411_reset = io_reset; // @[:@139438.4 RegFile.scala 76:16:@139445.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@139444.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@139448.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@139442.4]
  assign regs_412_clock = clock; // @[:@139451.4]
  assign regs_412_reset = io_reset; // @[:@139452.4 RegFile.scala 76:16:@139459.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@139458.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@139462.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@139456.4]
  assign regs_413_clock = clock; // @[:@139465.4]
  assign regs_413_reset = io_reset; // @[:@139466.4 RegFile.scala 76:16:@139473.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@139472.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@139476.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@139470.4]
  assign regs_414_clock = clock; // @[:@139479.4]
  assign regs_414_reset = io_reset; // @[:@139480.4 RegFile.scala 76:16:@139487.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@139486.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@139490.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@139484.4]
  assign regs_415_clock = clock; // @[:@139493.4]
  assign regs_415_reset = io_reset; // @[:@139494.4 RegFile.scala 76:16:@139501.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@139500.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@139504.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@139498.4]
  assign regs_416_clock = clock; // @[:@139507.4]
  assign regs_416_reset = io_reset; // @[:@139508.4 RegFile.scala 76:16:@139515.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@139514.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@139518.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@139512.4]
  assign regs_417_clock = clock; // @[:@139521.4]
  assign regs_417_reset = io_reset; // @[:@139522.4 RegFile.scala 76:16:@139529.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@139528.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@139532.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@139526.4]
  assign regs_418_clock = clock; // @[:@139535.4]
  assign regs_418_reset = io_reset; // @[:@139536.4 RegFile.scala 76:16:@139543.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@139542.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@139546.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@139540.4]
  assign regs_419_clock = clock; // @[:@139549.4]
  assign regs_419_reset = io_reset; // @[:@139550.4 RegFile.scala 76:16:@139557.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@139556.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@139560.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@139554.4]
  assign regs_420_clock = clock; // @[:@139563.4]
  assign regs_420_reset = io_reset; // @[:@139564.4 RegFile.scala 76:16:@139571.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@139570.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@139574.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@139568.4]
  assign regs_421_clock = clock; // @[:@139577.4]
  assign regs_421_reset = io_reset; // @[:@139578.4 RegFile.scala 76:16:@139585.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@139584.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@139588.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@139582.4]
  assign regs_422_clock = clock; // @[:@139591.4]
  assign regs_422_reset = io_reset; // @[:@139592.4 RegFile.scala 76:16:@139599.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@139598.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@139602.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@139596.4]
  assign regs_423_clock = clock; // @[:@139605.4]
  assign regs_423_reset = io_reset; // @[:@139606.4 RegFile.scala 76:16:@139613.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@139612.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@139616.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@139610.4]
  assign regs_424_clock = clock; // @[:@139619.4]
  assign regs_424_reset = io_reset; // @[:@139620.4 RegFile.scala 76:16:@139627.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@139626.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@139630.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@139624.4]
  assign regs_425_clock = clock; // @[:@139633.4]
  assign regs_425_reset = io_reset; // @[:@139634.4 RegFile.scala 76:16:@139641.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@139640.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@139644.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@139638.4]
  assign regs_426_clock = clock; // @[:@139647.4]
  assign regs_426_reset = io_reset; // @[:@139648.4 RegFile.scala 76:16:@139655.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@139654.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@139658.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@139652.4]
  assign regs_427_clock = clock; // @[:@139661.4]
  assign regs_427_reset = io_reset; // @[:@139662.4 RegFile.scala 76:16:@139669.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@139668.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@139672.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@139666.4]
  assign regs_428_clock = clock; // @[:@139675.4]
  assign regs_428_reset = io_reset; // @[:@139676.4 RegFile.scala 76:16:@139683.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@139682.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@139686.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@139680.4]
  assign regs_429_clock = clock; // @[:@139689.4]
  assign regs_429_reset = io_reset; // @[:@139690.4 RegFile.scala 76:16:@139697.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@139696.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@139700.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@139694.4]
  assign regs_430_clock = clock; // @[:@139703.4]
  assign regs_430_reset = io_reset; // @[:@139704.4 RegFile.scala 76:16:@139711.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@139710.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@139714.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@139708.4]
  assign regs_431_clock = clock; // @[:@139717.4]
  assign regs_431_reset = io_reset; // @[:@139718.4 RegFile.scala 76:16:@139725.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@139724.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@139728.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@139722.4]
  assign regs_432_clock = clock; // @[:@139731.4]
  assign regs_432_reset = io_reset; // @[:@139732.4 RegFile.scala 76:16:@139739.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@139738.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@139742.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@139736.4]
  assign regs_433_clock = clock; // @[:@139745.4]
  assign regs_433_reset = io_reset; // @[:@139746.4 RegFile.scala 76:16:@139753.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@139752.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@139756.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@139750.4]
  assign regs_434_clock = clock; // @[:@139759.4]
  assign regs_434_reset = io_reset; // @[:@139760.4 RegFile.scala 76:16:@139767.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@139766.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@139770.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@139764.4]
  assign regs_435_clock = clock; // @[:@139773.4]
  assign regs_435_reset = io_reset; // @[:@139774.4 RegFile.scala 76:16:@139781.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@139780.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@139784.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@139778.4]
  assign regs_436_clock = clock; // @[:@139787.4]
  assign regs_436_reset = io_reset; // @[:@139788.4 RegFile.scala 76:16:@139795.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@139794.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@139798.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@139792.4]
  assign regs_437_clock = clock; // @[:@139801.4]
  assign regs_437_reset = io_reset; // @[:@139802.4 RegFile.scala 76:16:@139809.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@139808.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@139812.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@139806.4]
  assign regs_438_clock = clock; // @[:@139815.4]
  assign regs_438_reset = io_reset; // @[:@139816.4 RegFile.scala 76:16:@139823.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@139822.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@139826.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@139820.4]
  assign regs_439_clock = clock; // @[:@139829.4]
  assign regs_439_reset = io_reset; // @[:@139830.4 RegFile.scala 76:16:@139837.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@139836.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@139840.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@139834.4]
  assign regs_440_clock = clock; // @[:@139843.4]
  assign regs_440_reset = io_reset; // @[:@139844.4 RegFile.scala 76:16:@139851.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@139850.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@139854.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@139848.4]
  assign regs_441_clock = clock; // @[:@139857.4]
  assign regs_441_reset = io_reset; // @[:@139858.4 RegFile.scala 76:16:@139865.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@139864.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@139868.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@139862.4]
  assign regs_442_clock = clock; // @[:@139871.4]
  assign regs_442_reset = io_reset; // @[:@139872.4 RegFile.scala 76:16:@139879.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@139878.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@139882.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@139876.4]
  assign regs_443_clock = clock; // @[:@139885.4]
  assign regs_443_reset = io_reset; // @[:@139886.4 RegFile.scala 76:16:@139893.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@139892.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@139896.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@139890.4]
  assign regs_444_clock = clock; // @[:@139899.4]
  assign regs_444_reset = io_reset; // @[:@139900.4 RegFile.scala 76:16:@139907.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@139906.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@139910.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@139904.4]
  assign regs_445_clock = clock; // @[:@139913.4]
  assign regs_445_reset = io_reset; // @[:@139914.4 RegFile.scala 76:16:@139921.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@139920.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@139924.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@139918.4]
  assign regs_446_clock = clock; // @[:@139927.4]
  assign regs_446_reset = io_reset; // @[:@139928.4 RegFile.scala 76:16:@139935.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@139934.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@139938.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@139932.4]
  assign regs_447_clock = clock; // @[:@139941.4]
  assign regs_447_reset = io_reset; // @[:@139942.4 RegFile.scala 76:16:@139949.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@139948.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@139952.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@139946.4]
  assign regs_448_clock = clock; // @[:@139955.4]
  assign regs_448_reset = io_reset; // @[:@139956.4 RegFile.scala 76:16:@139963.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@139962.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@139966.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@139960.4]
  assign regs_449_clock = clock; // @[:@139969.4]
  assign regs_449_reset = io_reset; // @[:@139970.4 RegFile.scala 76:16:@139977.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@139976.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@139980.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@139974.4]
  assign regs_450_clock = clock; // @[:@139983.4]
  assign regs_450_reset = io_reset; // @[:@139984.4 RegFile.scala 76:16:@139991.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@139990.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@139994.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@139988.4]
  assign regs_451_clock = clock; // @[:@139997.4]
  assign regs_451_reset = io_reset; // @[:@139998.4 RegFile.scala 76:16:@140005.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@140004.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@140008.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@140002.4]
  assign regs_452_clock = clock; // @[:@140011.4]
  assign regs_452_reset = io_reset; // @[:@140012.4 RegFile.scala 76:16:@140019.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@140018.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@140022.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@140016.4]
  assign regs_453_clock = clock; // @[:@140025.4]
  assign regs_453_reset = io_reset; // @[:@140026.4 RegFile.scala 76:16:@140033.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@140032.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@140036.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@140030.4]
  assign regs_454_clock = clock; // @[:@140039.4]
  assign regs_454_reset = io_reset; // @[:@140040.4 RegFile.scala 76:16:@140047.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@140046.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@140050.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@140044.4]
  assign regs_455_clock = clock; // @[:@140053.4]
  assign regs_455_reset = io_reset; // @[:@140054.4 RegFile.scala 76:16:@140061.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@140060.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@140064.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@140058.4]
  assign regs_456_clock = clock; // @[:@140067.4]
  assign regs_456_reset = io_reset; // @[:@140068.4 RegFile.scala 76:16:@140075.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@140074.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@140078.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@140072.4]
  assign regs_457_clock = clock; // @[:@140081.4]
  assign regs_457_reset = io_reset; // @[:@140082.4 RegFile.scala 76:16:@140089.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@140088.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@140092.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@140086.4]
  assign regs_458_clock = clock; // @[:@140095.4]
  assign regs_458_reset = io_reset; // @[:@140096.4 RegFile.scala 76:16:@140103.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@140102.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@140106.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@140100.4]
  assign regs_459_clock = clock; // @[:@140109.4]
  assign regs_459_reset = io_reset; // @[:@140110.4 RegFile.scala 76:16:@140117.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@140116.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@140120.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@140114.4]
  assign regs_460_clock = clock; // @[:@140123.4]
  assign regs_460_reset = io_reset; // @[:@140124.4 RegFile.scala 76:16:@140131.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@140130.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@140134.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@140128.4]
  assign regs_461_clock = clock; // @[:@140137.4]
  assign regs_461_reset = io_reset; // @[:@140138.4 RegFile.scala 76:16:@140145.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@140144.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@140148.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@140142.4]
  assign regs_462_clock = clock; // @[:@140151.4]
  assign regs_462_reset = io_reset; // @[:@140152.4 RegFile.scala 76:16:@140159.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@140158.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@140162.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@140156.4]
  assign regs_463_clock = clock; // @[:@140165.4]
  assign regs_463_reset = io_reset; // @[:@140166.4 RegFile.scala 76:16:@140173.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@140172.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@140176.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@140170.4]
  assign regs_464_clock = clock; // @[:@140179.4]
  assign regs_464_reset = io_reset; // @[:@140180.4 RegFile.scala 76:16:@140187.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@140186.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@140190.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@140184.4]
  assign regs_465_clock = clock; // @[:@140193.4]
  assign regs_465_reset = io_reset; // @[:@140194.4 RegFile.scala 76:16:@140201.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@140200.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@140204.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@140198.4]
  assign regs_466_clock = clock; // @[:@140207.4]
  assign regs_466_reset = io_reset; // @[:@140208.4 RegFile.scala 76:16:@140215.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@140214.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@140218.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@140212.4]
  assign regs_467_clock = clock; // @[:@140221.4]
  assign regs_467_reset = io_reset; // @[:@140222.4 RegFile.scala 76:16:@140229.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@140228.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@140232.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@140226.4]
  assign regs_468_clock = clock; // @[:@140235.4]
  assign regs_468_reset = io_reset; // @[:@140236.4 RegFile.scala 76:16:@140243.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@140242.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@140246.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@140240.4]
  assign regs_469_clock = clock; // @[:@140249.4]
  assign regs_469_reset = io_reset; // @[:@140250.4 RegFile.scala 76:16:@140257.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@140256.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@140260.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@140254.4]
  assign regs_470_clock = clock; // @[:@140263.4]
  assign regs_470_reset = io_reset; // @[:@140264.4 RegFile.scala 76:16:@140271.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@140270.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@140274.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@140268.4]
  assign regs_471_clock = clock; // @[:@140277.4]
  assign regs_471_reset = io_reset; // @[:@140278.4 RegFile.scala 76:16:@140285.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@140284.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@140288.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@140282.4]
  assign regs_472_clock = clock; // @[:@140291.4]
  assign regs_472_reset = io_reset; // @[:@140292.4 RegFile.scala 76:16:@140299.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@140298.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@140302.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@140296.4]
  assign regs_473_clock = clock; // @[:@140305.4]
  assign regs_473_reset = io_reset; // @[:@140306.4 RegFile.scala 76:16:@140313.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@140312.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@140316.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@140310.4]
  assign regs_474_clock = clock; // @[:@140319.4]
  assign regs_474_reset = io_reset; // @[:@140320.4 RegFile.scala 76:16:@140327.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@140326.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@140330.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@140324.4]
  assign regs_475_clock = clock; // @[:@140333.4]
  assign regs_475_reset = io_reset; // @[:@140334.4 RegFile.scala 76:16:@140341.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@140340.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@140344.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@140338.4]
  assign regs_476_clock = clock; // @[:@140347.4]
  assign regs_476_reset = io_reset; // @[:@140348.4 RegFile.scala 76:16:@140355.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@140354.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@140358.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@140352.4]
  assign regs_477_clock = clock; // @[:@140361.4]
  assign regs_477_reset = io_reset; // @[:@140362.4 RegFile.scala 76:16:@140369.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@140368.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@140372.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@140366.4]
  assign regs_478_clock = clock; // @[:@140375.4]
  assign regs_478_reset = io_reset; // @[:@140376.4 RegFile.scala 76:16:@140383.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@140382.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@140386.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@140380.4]
  assign regs_479_clock = clock; // @[:@140389.4]
  assign regs_479_reset = io_reset; // @[:@140390.4 RegFile.scala 76:16:@140397.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@140396.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@140400.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@140394.4]
  assign regs_480_clock = clock; // @[:@140403.4]
  assign regs_480_reset = io_reset; // @[:@140404.4 RegFile.scala 76:16:@140411.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@140410.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@140414.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@140408.4]
  assign regs_481_clock = clock; // @[:@140417.4]
  assign regs_481_reset = io_reset; // @[:@140418.4 RegFile.scala 76:16:@140425.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@140424.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@140428.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@140422.4]
  assign regs_482_clock = clock; // @[:@140431.4]
  assign regs_482_reset = io_reset; // @[:@140432.4 RegFile.scala 76:16:@140439.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@140438.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@140442.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@140436.4]
  assign regs_483_clock = clock; // @[:@140445.4]
  assign regs_483_reset = io_reset; // @[:@140446.4 RegFile.scala 76:16:@140453.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@140452.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@140456.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@140450.4]
  assign regs_484_clock = clock; // @[:@140459.4]
  assign regs_484_reset = io_reset; // @[:@140460.4 RegFile.scala 76:16:@140467.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@140466.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@140470.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@140464.4]
  assign regs_485_clock = clock; // @[:@140473.4]
  assign regs_485_reset = io_reset; // @[:@140474.4 RegFile.scala 76:16:@140481.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@140480.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@140484.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@140478.4]
  assign regs_486_clock = clock; // @[:@140487.4]
  assign regs_486_reset = io_reset; // @[:@140488.4 RegFile.scala 76:16:@140495.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@140494.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@140498.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@140492.4]
  assign regs_487_clock = clock; // @[:@140501.4]
  assign regs_487_reset = io_reset; // @[:@140502.4 RegFile.scala 76:16:@140509.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@140508.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@140512.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@140506.4]
  assign regs_488_clock = clock; // @[:@140515.4]
  assign regs_488_reset = io_reset; // @[:@140516.4 RegFile.scala 76:16:@140523.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@140522.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@140526.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@140520.4]
  assign regs_489_clock = clock; // @[:@140529.4]
  assign regs_489_reset = io_reset; // @[:@140530.4 RegFile.scala 76:16:@140537.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@140536.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@140540.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@140534.4]
  assign regs_490_clock = clock; // @[:@140543.4]
  assign regs_490_reset = io_reset; // @[:@140544.4 RegFile.scala 76:16:@140551.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@140550.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@140554.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@140548.4]
  assign regs_491_clock = clock; // @[:@140557.4]
  assign regs_491_reset = io_reset; // @[:@140558.4 RegFile.scala 76:16:@140565.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@140564.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@140568.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@140562.4]
  assign regs_492_clock = clock; // @[:@140571.4]
  assign regs_492_reset = io_reset; // @[:@140572.4 RegFile.scala 76:16:@140579.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@140578.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@140582.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@140576.4]
  assign regs_493_clock = clock; // @[:@140585.4]
  assign regs_493_reset = io_reset; // @[:@140586.4 RegFile.scala 76:16:@140593.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@140592.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@140596.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@140590.4]
  assign regs_494_clock = clock; // @[:@140599.4]
  assign regs_494_reset = io_reset; // @[:@140600.4 RegFile.scala 76:16:@140607.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@140606.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@140610.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@140604.4]
  assign regs_495_clock = clock; // @[:@140613.4]
  assign regs_495_reset = io_reset; // @[:@140614.4 RegFile.scala 76:16:@140621.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@140620.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@140624.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@140618.4]
  assign regs_496_clock = clock; // @[:@140627.4]
  assign regs_496_reset = io_reset; // @[:@140628.4 RegFile.scala 76:16:@140635.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@140634.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@140638.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@140632.4]
  assign regs_497_clock = clock; // @[:@140641.4]
  assign regs_497_reset = io_reset; // @[:@140642.4 RegFile.scala 76:16:@140649.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@140648.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@140652.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@140646.4]
  assign regs_498_clock = clock; // @[:@140655.4]
  assign regs_498_reset = io_reset; // @[:@140656.4 RegFile.scala 76:16:@140663.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@140662.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@140666.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@140660.4]
  assign regs_499_clock = clock; // @[:@140669.4]
  assign regs_499_reset = io_reset; // @[:@140670.4 RegFile.scala 76:16:@140677.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@140676.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@140680.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@140674.4]
  assign regs_500_clock = clock; // @[:@140683.4]
  assign regs_500_reset = io_reset; // @[:@140684.4 RegFile.scala 76:16:@140691.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@140690.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@140694.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@140688.4]
  assign regs_501_clock = clock; // @[:@140697.4]
  assign regs_501_reset = io_reset; // @[:@140698.4 RegFile.scala 76:16:@140705.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@140704.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@140708.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@140702.4]
  assign regs_502_clock = clock; // @[:@140711.4]
  assign regs_502_reset = io_reset; // @[:@140712.4 RegFile.scala 76:16:@140719.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@140718.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@140722.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@140716.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@141231.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@141232.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@141233.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@141234.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@141235.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@141236.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@141237.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@141238.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@141239.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@141240.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@141241.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@141242.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@141243.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@141244.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@141245.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@141246.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@141247.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@141248.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@141249.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@141250.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@141251.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@141252.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@141253.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@141254.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@141255.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@141256.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@141257.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@141258.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@141259.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@141260.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@141261.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@141262.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@141263.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@141264.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@141265.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@141266.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@141267.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@141268.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@141269.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@141270.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@141271.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@141272.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@141273.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@141274.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@141275.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@141276.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@141277.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@141278.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@141279.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@141280.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@141281.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@141282.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@141283.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@141284.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@141285.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@141286.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@141287.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@141288.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@141289.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@141290.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@141291.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@141292.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@141293.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@141294.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@141295.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@141296.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@141297.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@141298.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@141299.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@141300.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@141301.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@141302.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@141303.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@141304.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@141305.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@141306.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@141307.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@141308.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@141309.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@141310.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@141311.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@141312.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@141313.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@141314.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@141315.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@141316.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@141317.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@141318.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@141319.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@141320.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@141321.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@141322.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@141323.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@141324.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@141325.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@141326.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@141327.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@141328.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@141329.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@141330.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@141331.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@141332.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@141333.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@141334.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@141335.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@141336.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@141337.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@141338.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@141339.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@141340.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@141341.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@141342.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@141343.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@141344.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@141345.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@141346.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@141347.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@141348.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@141349.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@141350.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@141351.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@141352.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@141353.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@141354.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@141355.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@141356.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@141357.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@141358.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@141359.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@141360.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@141361.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@141362.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@141363.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@141364.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@141365.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@141366.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@141367.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@141368.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@141369.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@141370.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@141371.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@141372.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@141373.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@141374.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@141375.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@141376.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@141377.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@141378.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@141379.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@141380.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@141381.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@141382.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@141383.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@141384.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@141385.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@141386.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@141387.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@141388.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@141389.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@141390.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@141391.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@141392.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@141393.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@141394.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@141395.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@141396.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@141397.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@141398.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@141399.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@141400.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@141401.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@141402.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@141403.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@141404.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@141405.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@141406.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@141407.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@141408.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@141409.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@141410.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@141411.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@141412.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@141413.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@141414.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@141415.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@141416.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@141417.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@141418.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@141419.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@141420.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@141421.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@141422.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@141423.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@141424.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@141425.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@141426.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@141427.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@141428.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@141429.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@141430.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@141431.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@141432.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@141433.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@141434.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@141435.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@141436.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@141437.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@141438.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@141439.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@141440.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@141441.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@141442.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@141443.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@141444.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@141445.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@141446.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@141447.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@141448.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@141449.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@141450.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@141451.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@141452.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@141453.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@141454.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@141455.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@141456.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@141457.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@141458.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@141459.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@141460.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@141461.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@141462.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@141463.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@141464.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@141465.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@141466.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@141467.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@141468.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@141469.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@141470.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@141471.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@141472.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@141473.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@141474.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@141475.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@141476.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@141477.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@141478.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@141479.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@141480.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@141481.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@141482.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@141483.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@141484.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@141485.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@141486.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@141487.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@141488.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@141489.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@141490.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@141491.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@141492.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@141493.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@141494.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@141495.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@141496.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@141497.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@141498.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@141499.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@141500.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@141501.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@141502.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@141503.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@141504.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@141505.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@141506.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@141507.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@141508.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@141509.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@141510.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@141511.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@141512.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@141513.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@141514.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@141515.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@141516.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@141517.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@141518.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@141519.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@141520.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@141521.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@141522.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@141523.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@141524.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@141525.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@141526.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@141527.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@141528.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@141529.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@141530.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@141531.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@141532.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@141533.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@141534.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@141535.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@141536.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@141537.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@141538.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@141539.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@141540.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@141541.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@141542.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@141543.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@141544.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@141545.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@141546.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@141547.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@141548.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@141549.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@141550.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@141551.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@141552.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@141553.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@141554.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@141555.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@141556.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@141557.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@141558.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@141559.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@141560.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@141561.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@141562.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@141563.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@141564.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@141565.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@141566.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@141567.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@141568.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@141569.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@141570.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@141571.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@141572.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@141573.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@141574.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@141575.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@141576.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@141577.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@141578.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@141579.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@141580.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@141581.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@141582.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@141583.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@141584.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@141585.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@141586.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@141587.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@141588.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@141589.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@141590.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@141591.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@141592.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@141593.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@141594.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@141595.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@141596.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@141597.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@141598.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@141599.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@141600.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@141601.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@141602.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@141603.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@141604.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@141605.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@141606.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@141607.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@141608.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@141609.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@141610.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@141611.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@141612.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@141613.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@141614.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@141615.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@141616.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@141617.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@141618.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@141619.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@141620.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@141621.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@141622.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@141623.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@141624.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@141625.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@141626.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@141627.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@141628.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@141629.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@141630.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@141631.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@141632.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@141633.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@141634.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@141635.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@141636.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@141637.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@141638.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@141639.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@141640.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@141641.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@141642.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@141643.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@141644.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@141645.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@141646.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@141647.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@141648.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@141649.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@141650.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@141651.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@141652.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@141653.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@141654.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@141655.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@141656.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@141657.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@141658.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@141659.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@141660.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@141661.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@141662.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@141663.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@141664.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@141665.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@141666.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@141667.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@141668.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@141669.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@141670.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@141671.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@141672.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@141673.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@141674.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@141675.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@141676.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@141677.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@141678.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@141679.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@141680.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@141681.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@141682.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@141683.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@141684.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@141685.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@141686.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@141687.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@141688.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@141689.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@141690.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@141691.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@141692.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@141693.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@141694.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@141695.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@141696.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@141697.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@141698.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@141699.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@141700.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@141701.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@141702.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@141703.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@141704.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@141705.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@141706.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@141707.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@141708.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@141709.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@141710.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@141711.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@141712.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@141713.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@141714.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@141715.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@141716.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@141717.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@141718.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@141719.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@141720.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@141721.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@141722.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@141723.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@141724.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@141725.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@141726.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@141727.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@141728.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@141729.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@141730.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@141731.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@141732.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@141733.4]
  assign rport_io_sel = io_raddr[8:0]; // @[RegFile.scala 106:18:@141734.4]
endmodule
module RetimeWrapper_914( // @[:@141758.2]
  input         clock, // @[:@141759.4]
  input         reset, // @[:@141760.4]
  input  [39:0] io_in, // @[:@141761.4]
  output [39:0] io_out // @[:@141761.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@141763.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@141763.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@141763.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@141763.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@141763.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@141763.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@141763.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@141776.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@141775.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@141774.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@141773.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@141772.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@141770.4]
endmodule
module FringeFF_503( // @[:@141778.2]
  input         clock, // @[:@141779.4]
  input         reset, // @[:@141780.4]
  input  [39:0] io_in, // @[:@141781.4]
  output [39:0] io_out, // @[:@141781.4]
  input         io_enable // @[:@141781.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@141784.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@141784.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@141784.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@141784.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@141789.4 package.scala 96:25:@141790.4]
  RetimeWrapper_914 RetimeWrapper ( // @[package.scala 93:22:@141784.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@141789.4 package.scala 96:25:@141790.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@141801.4]
  assign RetimeWrapper_clock = clock; // @[:@141785.4]
  assign RetimeWrapper_reset = reset; // @[:@141786.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@141787.4]
endmodule
module FringeCounter( // @[:@141803.2]
  input   clock, // @[:@141804.4]
  input   reset, // @[:@141805.4]
  input   io_enable, // @[:@141806.4]
  output  io_done // @[:@141806.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@141808.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@141808.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@141808.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@141808.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@141808.4]
  wire [40:0] count; // @[Cat.scala 30:58:@141815.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@141816.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@141817.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@141818.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@141820.4]
  FringeFF_503 reg$ ( // @[FringeCounter.scala 24:19:@141808.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@141815.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@141816.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@141817.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@141818.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@141820.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@141831.4]
  assign reg$_clock = clock; // @[:@141809.4]
  assign reg$_reset = reset; // @[:@141810.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@141822.6 FringeCounter.scala 37:15:@141825.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@141813.4]
endmodule
module FringeFF_504( // @[:@141865.2]
  input   clock, // @[:@141866.4]
  input   reset, // @[:@141867.4]
  input   io_in, // @[:@141868.4]
  input   io_reset, // @[:@141868.4]
  output  io_out, // @[:@141868.4]
  input   io_enable // @[:@141868.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@141871.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@141871.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@141871.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@141871.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@141871.4]
  wire  _T_18; // @[package.scala 96:25:@141876.4 package.scala 96:25:@141877.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@141882.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@141871.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@141876.4 package.scala 96:25:@141877.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@141882.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@141888.4]
  assign RetimeWrapper_clock = clock; // @[:@141872.4]
  assign RetimeWrapper_reset = reset; // @[:@141873.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@141875.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@141874.4]
endmodule
module Depulser( // @[:@141890.2]
  input   clock, // @[:@141891.4]
  input   reset, // @[:@141892.4]
  input   io_in, // @[:@141893.4]
  input   io_rst, // @[:@141893.4]
  output  io_out // @[:@141893.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@141895.4]
  wire  r_reset; // @[Depulser.scala 14:17:@141895.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@141895.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@141895.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@141895.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@141895.4]
  FringeFF_504 r ( // @[Depulser.scala 14:17:@141895.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@141904.4]
  assign r_clock = clock; // @[:@141896.4]
  assign r_reset = reset; // @[:@141897.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@141899.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@141903.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@141902.4]
endmodule
module Fringe( // @[:@141906.2]
  input         clock, // @[:@141907.4]
  input         reset, // @[:@141908.4]
  input  [31:0] io_raddr, // @[:@141909.4]
  input         io_wen, // @[:@141909.4]
  input  [31:0] io_waddr, // @[:@141909.4]
  input  [63:0] io_wdata, // @[:@141909.4]
  output [63:0] io_rdata, // @[:@141909.4]
  output        io_enable, // @[:@141909.4]
  input         io_done, // @[:@141909.4]
  output        io_reset, // @[:@141909.4]
  output [63:0] io_argIns_0, // @[:@141909.4]
  output [63:0] io_argIns_1, // @[:@141909.4]
  input         io_argOuts_0_valid, // @[:@141909.4]
  input  [63:0] io_argOuts_0_bits, // @[:@141909.4]
  output        io_memStreams_stores_0_cmd_ready, // @[:@141909.4]
  input         io_memStreams_stores_0_cmd_valid, // @[:@141909.4]
  input  [63:0] io_memStreams_stores_0_cmd_bits_addr, // @[:@141909.4]
  input  [31:0] io_memStreams_stores_0_cmd_bits_size, // @[:@141909.4]
  output        io_memStreams_stores_0_data_ready, // @[:@141909.4]
  input         io_memStreams_stores_0_data_valid, // @[:@141909.4]
  input  [31:0] io_memStreams_stores_0_data_bits_wdata_0, // @[:@141909.4]
  input         io_memStreams_stores_0_data_bits_wstrb, // @[:@141909.4]
  input         io_memStreams_stores_0_wresp_ready, // @[:@141909.4]
  output        io_memStreams_stores_0_wresp_valid, // @[:@141909.4]
  output        io_memStreams_stores_0_wresp_bits, // @[:@141909.4]
  input         io_dram_0_cmd_ready, // @[:@141909.4]
  output        io_dram_0_cmd_valid, // @[:@141909.4]
  output [63:0] io_dram_0_cmd_bits_addr, // @[:@141909.4]
  output [31:0] io_dram_0_cmd_bits_size, // @[:@141909.4]
  output        io_dram_0_cmd_bits_isWr, // @[:@141909.4]
  output [31:0] io_dram_0_cmd_bits_tag, // @[:@141909.4]
  input         io_dram_0_wdata_ready, // @[:@141909.4]
  output        io_dram_0_wdata_valid, // @[:@141909.4]
  output [31:0] io_dram_0_wdata_bits_wdata_0, // @[:@141909.4]
  output [31:0] io_dram_0_wdata_bits_wdata_1, // @[:@141909.4]
  output [31:0] io_dram_0_wdata_bits_wdata_2, // @[:@141909.4]
  output [31:0] io_dram_0_wdata_bits_wdata_3, // @[:@141909.4]
  output [31:0] io_dram_0_wdata_bits_wdata_4, // @[:@141909.4]
  output [31:0] io_dram_0_wdata_bits_wdata_5, // @[:@141909.4]
  output [31:0] io_dram_0_wdata_bits_wdata_6, // @[:@141909.4]
  output [31:0] io_dram_0_wdata_bits_wdata_7, // @[:@141909.4]
  output [31:0] io_dram_0_wdata_bits_wdata_8, // @[:@141909.4]
  output [31:0] io_dram_0_wdata_bits_wdata_9, // @[:@141909.4]
  output [31:0] io_dram_0_wdata_bits_wdata_10, // @[:@141909.4]
  output [31:0] io_dram_0_wdata_bits_wdata_11, // @[:@141909.4]
  output [31:0] io_dram_0_wdata_bits_wdata_12, // @[:@141909.4]
  output [31:0] io_dram_0_wdata_bits_wdata_13, // @[:@141909.4]
  output [31:0] io_dram_0_wdata_bits_wdata_14, // @[:@141909.4]
  output [31:0] io_dram_0_wdata_bits_wdata_15, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_0, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_1, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_2, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_3, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_4, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_5, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_6, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_7, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_8, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_9, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_10, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_11, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_12, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_13, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_14, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_15, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_16, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_17, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_18, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_19, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_20, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_21, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_22, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_23, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_24, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_25, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_26, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_27, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_28, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_29, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_30, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_31, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_32, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_33, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_34, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_35, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_36, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_37, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_38, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_39, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_40, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_41, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_42, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_43, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_44, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_45, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_46, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_47, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_48, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_49, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_50, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_51, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_52, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_53, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_54, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_55, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_56, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_57, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_58, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_59, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_60, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_61, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_62, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wstrb_63, // @[:@141909.4]
  output        io_dram_0_wdata_bits_wlast, // @[:@141909.4]
  output        io_dram_0_rresp_ready, // @[:@141909.4]
  output        io_dram_0_wresp_ready, // @[:@141909.4]
  input         io_dram_0_wresp_valid, // @[:@141909.4]
  input  [31:0] io_dram_0_wresp_bits_tag, // @[:@141909.4]
  input         io_dram_1_cmd_ready, // @[:@141909.4]
  output        io_dram_1_cmd_valid, // @[:@141909.4]
  output [63:0] io_dram_1_cmd_bits_addr, // @[:@141909.4]
  output [31:0] io_dram_1_cmd_bits_size, // @[:@141909.4]
  output        io_dram_1_cmd_bits_isWr, // @[:@141909.4]
  output [31:0] io_dram_1_cmd_bits_tag, // @[:@141909.4]
  input         io_dram_1_wdata_ready, // @[:@141909.4]
  output        io_dram_1_wdata_valid, // @[:@141909.4]
  output [31:0] io_dram_1_wdata_bits_wdata_0, // @[:@141909.4]
  output [31:0] io_dram_1_wdata_bits_wdata_1, // @[:@141909.4]
  output [31:0] io_dram_1_wdata_bits_wdata_2, // @[:@141909.4]
  output [31:0] io_dram_1_wdata_bits_wdata_3, // @[:@141909.4]
  output [31:0] io_dram_1_wdata_bits_wdata_4, // @[:@141909.4]
  output [31:0] io_dram_1_wdata_bits_wdata_5, // @[:@141909.4]
  output [31:0] io_dram_1_wdata_bits_wdata_6, // @[:@141909.4]
  output [31:0] io_dram_1_wdata_bits_wdata_7, // @[:@141909.4]
  output [31:0] io_dram_1_wdata_bits_wdata_8, // @[:@141909.4]
  output [31:0] io_dram_1_wdata_bits_wdata_9, // @[:@141909.4]
  output [31:0] io_dram_1_wdata_bits_wdata_10, // @[:@141909.4]
  output [31:0] io_dram_1_wdata_bits_wdata_11, // @[:@141909.4]
  output [31:0] io_dram_1_wdata_bits_wdata_12, // @[:@141909.4]
  output [31:0] io_dram_1_wdata_bits_wdata_13, // @[:@141909.4]
  output [31:0] io_dram_1_wdata_bits_wdata_14, // @[:@141909.4]
  output [31:0] io_dram_1_wdata_bits_wdata_15, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_0, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_1, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_2, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_3, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_4, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_5, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_6, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_7, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_8, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_9, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_10, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_11, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_12, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_13, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_14, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_15, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_16, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_17, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_18, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_19, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_20, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_21, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_22, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_23, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_24, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_25, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_26, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_27, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_28, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_29, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_30, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_31, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_32, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_33, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_34, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_35, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_36, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_37, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_38, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_39, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_40, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_41, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_42, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_43, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_44, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_45, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_46, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_47, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_48, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_49, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_50, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_51, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_52, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_53, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_54, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_55, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_56, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_57, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_58, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_59, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_60, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_61, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_62, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wstrb_63, // @[:@141909.4]
  output        io_dram_1_wdata_bits_wlast, // @[:@141909.4]
  output        io_dram_1_rresp_ready, // @[:@141909.4]
  output        io_dram_1_wresp_ready, // @[:@141909.4]
  input         io_dram_1_wresp_valid, // @[:@141909.4]
  input  [31:0] io_dram_1_wresp_bits_tag, // @[:@141909.4]
  input         io_dram_2_cmd_ready, // @[:@141909.4]
  output        io_dram_2_cmd_valid, // @[:@141909.4]
  output [63:0] io_dram_2_cmd_bits_addr, // @[:@141909.4]
  output [31:0] io_dram_2_cmd_bits_size, // @[:@141909.4]
  output        io_dram_2_cmd_bits_isWr, // @[:@141909.4]
  output [31:0] io_dram_2_cmd_bits_tag, // @[:@141909.4]
  input         io_dram_2_wdata_ready, // @[:@141909.4]
  output        io_dram_2_wdata_valid, // @[:@141909.4]
  output [31:0] io_dram_2_wdata_bits_wdata_0, // @[:@141909.4]
  output [31:0] io_dram_2_wdata_bits_wdata_1, // @[:@141909.4]
  output [31:0] io_dram_2_wdata_bits_wdata_2, // @[:@141909.4]
  output [31:0] io_dram_2_wdata_bits_wdata_3, // @[:@141909.4]
  output [31:0] io_dram_2_wdata_bits_wdata_4, // @[:@141909.4]
  output [31:0] io_dram_2_wdata_bits_wdata_5, // @[:@141909.4]
  output [31:0] io_dram_2_wdata_bits_wdata_6, // @[:@141909.4]
  output [31:0] io_dram_2_wdata_bits_wdata_7, // @[:@141909.4]
  output [31:0] io_dram_2_wdata_bits_wdata_8, // @[:@141909.4]
  output [31:0] io_dram_2_wdata_bits_wdata_9, // @[:@141909.4]
  output [31:0] io_dram_2_wdata_bits_wdata_10, // @[:@141909.4]
  output [31:0] io_dram_2_wdata_bits_wdata_11, // @[:@141909.4]
  output [31:0] io_dram_2_wdata_bits_wdata_12, // @[:@141909.4]
  output [31:0] io_dram_2_wdata_bits_wdata_13, // @[:@141909.4]
  output [31:0] io_dram_2_wdata_bits_wdata_14, // @[:@141909.4]
  output [31:0] io_dram_2_wdata_bits_wdata_15, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_0, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_1, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_2, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_3, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_4, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_5, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_6, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_7, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_8, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_9, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_10, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_11, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_12, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_13, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_14, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_15, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_16, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_17, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_18, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_19, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_20, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_21, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_22, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_23, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_24, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_25, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_26, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_27, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_28, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_29, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_30, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_31, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_32, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_33, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_34, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_35, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_36, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_37, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_38, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_39, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_40, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_41, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_42, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_43, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_44, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_45, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_46, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_47, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_48, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_49, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_50, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_51, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_52, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_53, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_54, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_55, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_56, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_57, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_58, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_59, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_60, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_61, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_62, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wstrb_63, // @[:@141909.4]
  output        io_dram_2_wdata_bits_wlast, // @[:@141909.4]
  output        io_dram_2_rresp_ready, // @[:@141909.4]
  output        io_dram_2_wresp_ready, // @[:@141909.4]
  input         io_dram_2_wresp_valid, // @[:@141909.4]
  input  [31:0] io_dram_2_wresp_bits_tag, // @[:@141909.4]
  input         io_dram_3_cmd_ready, // @[:@141909.4]
  output        io_dram_3_cmd_valid, // @[:@141909.4]
  output [63:0] io_dram_3_cmd_bits_addr, // @[:@141909.4]
  output [31:0] io_dram_3_cmd_bits_size, // @[:@141909.4]
  output        io_dram_3_cmd_bits_isWr, // @[:@141909.4]
  output [31:0] io_dram_3_cmd_bits_tag, // @[:@141909.4]
  input         io_dram_3_wdata_ready, // @[:@141909.4]
  output        io_dram_3_wdata_valid, // @[:@141909.4]
  output [31:0] io_dram_3_wdata_bits_wdata_0, // @[:@141909.4]
  output [31:0] io_dram_3_wdata_bits_wdata_1, // @[:@141909.4]
  output [31:0] io_dram_3_wdata_bits_wdata_2, // @[:@141909.4]
  output [31:0] io_dram_3_wdata_bits_wdata_3, // @[:@141909.4]
  output [31:0] io_dram_3_wdata_bits_wdata_4, // @[:@141909.4]
  output [31:0] io_dram_3_wdata_bits_wdata_5, // @[:@141909.4]
  output [31:0] io_dram_3_wdata_bits_wdata_6, // @[:@141909.4]
  output [31:0] io_dram_3_wdata_bits_wdata_7, // @[:@141909.4]
  output [31:0] io_dram_3_wdata_bits_wdata_8, // @[:@141909.4]
  output [31:0] io_dram_3_wdata_bits_wdata_9, // @[:@141909.4]
  output [31:0] io_dram_3_wdata_bits_wdata_10, // @[:@141909.4]
  output [31:0] io_dram_3_wdata_bits_wdata_11, // @[:@141909.4]
  output [31:0] io_dram_3_wdata_bits_wdata_12, // @[:@141909.4]
  output [31:0] io_dram_3_wdata_bits_wdata_13, // @[:@141909.4]
  output [31:0] io_dram_3_wdata_bits_wdata_14, // @[:@141909.4]
  output [31:0] io_dram_3_wdata_bits_wdata_15, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_0, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_1, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_2, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_3, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_4, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_5, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_6, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_7, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_8, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_9, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_10, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_11, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_12, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_13, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_14, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_15, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_16, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_17, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_18, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_19, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_20, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_21, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_22, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_23, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_24, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_25, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_26, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_27, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_28, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_29, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_30, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_31, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_32, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_33, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_34, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_35, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_36, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_37, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_38, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_39, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_40, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_41, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_42, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_43, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_44, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_45, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_46, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_47, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_48, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_49, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_50, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_51, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_52, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_53, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_54, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_55, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_56, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_57, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_58, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_59, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_60, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_61, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_62, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wstrb_63, // @[:@141909.4]
  output        io_dram_3_wdata_bits_wlast, // @[:@141909.4]
  output        io_dram_3_rresp_ready, // @[:@141909.4]
  output        io_dram_3_wresp_ready, // @[:@141909.4]
  input         io_dram_3_wresp_valid, // @[:@141909.4]
  input  [31:0] io_dram_3_wresp_bits_tag, // @[:@141909.4]
  input         io_heap_0_req_valid, // @[:@141909.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@141909.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@141909.4]
  output        io_heap_0_resp_valid, // @[:@141909.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@141909.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@141909.4]
);
  wire  dramArbs_0_clock; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_reset; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_enable; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_app_stores_0_cmd_valid; // @[Fringe.scala 91:25:@141915.4]
  wire [63:0] dramArbs_0_io_app_stores_0_cmd_bits_addr; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_app_stores_0_cmd_bits_size; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_app_stores_0_data_valid; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_app_stores_0_data_bits_wdata_0; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_app_stores_0_data_bits_wstrb; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_app_stores_0_wresp_ready; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_cmd_ready; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 91:25:@141915.4]
  wire [63:0] dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_ready; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_0_io_dram_wresp_valid; // @[Fringe.scala 91:25:@141915.4]
  wire [31:0] dramArbs_0_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@141915.4]
  wire  dramArbs_1_clock; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_reset; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_enable; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_cmd_ready; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 91:25:@142908.4]
  wire [63:0] dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_ready; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_1_io_dram_wresp_valid; // @[Fringe.scala 91:25:@142908.4]
  wire [31:0] dramArbs_1_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@142908.4]
  wire  dramArbs_2_clock; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_reset; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_enable; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_cmd_ready; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 91:25:@143868.4]
  wire [63:0] dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_ready; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_2_io_dram_wresp_valid; // @[Fringe.scala 91:25:@143868.4]
  wire [31:0] dramArbs_2_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@143868.4]
  wire  dramArbs_3_clock; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_reset; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_enable; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_cmd_ready; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 91:25:@144828.4]
  wire [63:0] dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_ready; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 91:25:@144828.4]
  wire  dramArbs_3_io_dram_wresp_valid; // @[Fringe.scala 91:25:@144828.4]
  wire [31:0] dramArbs_3_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@144828.4]
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@145788.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@145788.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@145788.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@145788.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@145788.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@145788.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@145788.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@145788.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@145788.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@145788.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@145788.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@145788.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@145797.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@145797.4]
  wire [31:0] regs_io_raddr; // @[Fringe.scala 116:20:@145797.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@145797.4]
  wire [31:0] regs_io_waddr; // @[Fringe.scala 116:20:@145797.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@145797.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@145797.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@145797.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@145797.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@145797.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@145797.4]
  wire [63:0] regs_io_argIns_3; // @[Fringe.scala 116:20:@145797.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@145797.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@145797.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@145797.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@145797.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@147847.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@147847.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@147847.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@147847.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@147866.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@147866.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@147866.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@147866.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@147866.4]
  wire [63:0] _T_1020; // @[:@147824.4 :@147825.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@147826.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@147828.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@147830.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@147832.4]
  wire  _T_1025; // @[Fringe.scala 134:28:@147834.4]
  wire  _T_1029; // @[Fringe.scala 134:42:@147836.4]
  wire  _T_1030; // @[Fringe.scala 135:27:@147838.4]
  wire [63:0] _T_1040; // @[Fringe.scala 156:22:@147874.4]
  reg  _T_1047; // @[package.scala 152:20:@147877.4]
  reg [31:0] _RAND_0;
  wire  _T_1048; // @[package.scala 153:13:@147879.4]
  wire  _T_1049; // @[package.scala 153:8:@147880.4]
  wire  _T_1052; // @[Fringe.scala 160:55:@147884.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@147885.4]
  wire  _T_1055; // @[Fringe.scala 161:58:@147888.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@147889.4]
  wire [1:0] _T_1059; // @[Fringe.scala 162:57:@147891.4]
  wire [1:0] _T_1061; // @[Fringe.scala 162:34:@147892.4]
  wire [63:0] _T_1063; // @[Fringe.scala 163:30:@147894.4]
  wire [1:0] _T_1064; // @[Fringe.scala 171:37:@147897.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@147876.4 Fringe.scala 163:24:@147895.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@147876.4 Fringe.scala 162:28:@147893.4]
  wire [61:0] _T_1065; // @[Fringe.scala 171:37:@147898.4]
  wire  alloc; // @[Fringe.scala 202:38:@149528.4]
  wire  dealloc; // @[Fringe.scala 203:40:@149529.4]
  wire  _T_1569; // @[Fringe.scala 204:37:@149530.4]
  reg  _T_1572; // @[package.scala 152:20:@149531.4]
  reg [31:0] _RAND_1;
  wire  _T_1573; // @[package.scala 153:13:@149533.4]
  DRAMArbiter dramArbs_0 ( // @[Fringe.scala 91:25:@141915.4]
    .clock(dramArbs_0_clock),
    .reset(dramArbs_0_reset),
    .io_enable(dramArbs_0_io_enable),
    .io_app_stores_0_cmd_ready(dramArbs_0_io_app_stores_0_cmd_ready),
    .io_app_stores_0_cmd_valid(dramArbs_0_io_app_stores_0_cmd_valid),
    .io_app_stores_0_cmd_bits_addr(dramArbs_0_io_app_stores_0_cmd_bits_addr),
    .io_app_stores_0_cmd_bits_size(dramArbs_0_io_app_stores_0_cmd_bits_size),
    .io_app_stores_0_data_ready(dramArbs_0_io_app_stores_0_data_ready),
    .io_app_stores_0_data_valid(dramArbs_0_io_app_stores_0_data_valid),
    .io_app_stores_0_data_bits_wdata_0(dramArbs_0_io_app_stores_0_data_bits_wdata_0),
    .io_app_stores_0_data_bits_wstrb(dramArbs_0_io_app_stores_0_data_bits_wstrb),
    .io_app_stores_0_wresp_ready(dramArbs_0_io_app_stores_0_wresp_ready),
    .io_app_stores_0_wresp_valid(dramArbs_0_io_app_stores_0_wresp_valid),
    .io_app_stores_0_wresp_bits(dramArbs_0_io_app_stores_0_wresp_bits),
    .io_dram_cmd_ready(dramArbs_0_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_0_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_0_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_0_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_0_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_0_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_0_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_0_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_0_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_0_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_0_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_0_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_0_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_0_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_0_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_0_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_0_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_0_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_0_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_0_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_0_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_0_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_0_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_0_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_0_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_0_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_0_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_0_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_0_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_0_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_0_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_0_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_0_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_0_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_0_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_0_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_0_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_0_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_0_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_0_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_0_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_0_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_0_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_0_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_0_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_0_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_0_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_0_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_0_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_0_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_0_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_0_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_0_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_0_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_0_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_0_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_0_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_0_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_0_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_0_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_0_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_0_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_0_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_0_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_0_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_0_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_0_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_0_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_0_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_0_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_0_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_0_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_0_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_0_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_0_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_0_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_0_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_0_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_0_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_0_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_0_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_0_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_0_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_0_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_0_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_0_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_0_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_0_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_0_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_0_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_0_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_0_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_0_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_1 ( // @[Fringe.scala 91:25:@142908.4]
    .clock(dramArbs_1_clock),
    .reset(dramArbs_1_reset),
    .io_enable(dramArbs_1_io_enable),
    .io_dram_cmd_ready(dramArbs_1_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_1_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_1_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_1_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_1_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_1_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_1_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_1_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_1_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_1_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_1_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_1_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_1_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_1_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_1_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_1_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_1_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_1_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_1_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_1_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_1_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_1_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_1_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_1_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_1_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_1_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_1_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_1_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_1_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_1_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_1_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_1_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_1_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_1_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_1_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_1_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_1_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_1_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_1_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_1_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_1_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_1_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_1_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_1_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_1_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_1_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_1_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_1_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_1_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_1_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_1_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_1_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_1_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_1_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_1_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_1_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_1_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_1_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_1_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_1_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_1_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_1_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_1_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_1_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_1_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_1_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_1_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_1_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_1_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_1_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_1_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_1_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_1_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_1_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_1_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_1_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_1_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_1_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_1_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_1_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_1_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_1_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_1_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_1_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_1_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_1_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_1_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_1_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_1_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_1_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_1_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_1_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_1_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_2 ( // @[Fringe.scala 91:25:@143868.4]
    .clock(dramArbs_2_clock),
    .reset(dramArbs_2_reset),
    .io_enable(dramArbs_2_io_enable),
    .io_dram_cmd_ready(dramArbs_2_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_2_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_2_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_2_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_2_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_2_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_2_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_2_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_2_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_2_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_2_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_2_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_2_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_2_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_2_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_2_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_2_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_2_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_2_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_2_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_2_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_2_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_2_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_2_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_2_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_2_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_2_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_2_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_2_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_2_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_2_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_2_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_2_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_2_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_2_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_2_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_2_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_2_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_2_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_2_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_2_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_2_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_2_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_2_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_2_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_2_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_2_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_2_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_2_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_2_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_2_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_2_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_2_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_2_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_2_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_2_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_2_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_2_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_2_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_2_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_2_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_2_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_2_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_2_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_2_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_2_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_2_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_2_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_2_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_2_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_2_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_2_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_2_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_2_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_2_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_2_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_2_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_2_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_2_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_2_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_2_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_2_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_2_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_2_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_2_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_2_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_2_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_2_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_2_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_2_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_2_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_2_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_2_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_3 ( // @[Fringe.scala 91:25:@144828.4]
    .clock(dramArbs_3_clock),
    .reset(dramArbs_3_reset),
    .io_enable(dramArbs_3_io_enable),
    .io_dram_cmd_ready(dramArbs_3_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_3_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_3_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_3_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_3_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_3_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_3_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_3_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_3_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_3_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_3_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_3_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_3_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_3_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_3_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_3_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_3_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_3_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_3_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_3_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_3_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_3_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_3_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_3_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_3_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_3_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_3_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_3_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_3_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_3_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_3_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_3_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_3_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_3_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_3_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_3_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_3_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_3_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_3_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_3_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_3_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_3_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_3_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_3_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_3_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_3_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_3_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_3_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_3_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_3_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_3_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_3_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_3_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_3_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_3_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_3_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_3_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_3_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_3_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_3_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_3_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_3_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_3_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_3_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_3_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_3_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_3_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_3_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_3_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_3_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_3_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_3_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_3_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_3_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_3_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_3_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_3_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_3_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_3_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_3_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_3_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_3_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_3_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_3_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_3_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_3_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_3_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_3_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_3_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_3_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_3_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_3_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_3_io_dram_wresp_bits_tag)
  );
  DRAMHeap heap ( // @[Fringe.scala 107:20:@145788.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@145797.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argIns_3(regs_io_argIns_3),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@147847.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@147866.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_1020 = regs_io_argIns_1; // @[:@147824.4 :@147825.4]
  assign curStatus_done = _T_1020[0]; // @[Fringe.scala 133:45:@147826.4]
  assign curStatus_timeout = _T_1020[1]; // @[Fringe.scala 133:45:@147828.4]
  assign curStatus_allocDealloc = _T_1020[4:2]; // @[Fringe.scala 133:45:@147830.4]
  assign curStatus_sizeAddr = _T_1020[63:5]; // @[Fringe.scala 133:45:@147832.4]
  assign _T_1025 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@147834.4]
  assign _T_1029 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@147836.4]
  assign _T_1030 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@147838.4]
  assign _T_1040 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@147874.4]
  assign _T_1048 = _T_1047 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@147879.4]
  assign _T_1049 = heap_io_host_0_req_valid & _T_1048; // @[package.scala 153:8:@147880.4]
  assign _T_1052 = _T_1025 & depulser_io_out; // @[Fringe.scala 160:55:@147884.4]
  assign status_bits_done = depulser_io_out ? _T_1052 : curStatus_done; // @[Fringe.scala 160:26:@147885.4]
  assign _T_1055 = _T_1025 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@147888.4]
  assign status_bits_timeout = depulser_io_out ? _T_1055 : curStatus_timeout; // @[Fringe.scala 161:29:@147889.4]
  assign _T_1059 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@147891.4]
  assign _T_1061 = heap_io_host_0_req_valid ? _T_1059 : 2'h0; // @[Fringe.scala 162:34:@147892.4]
  assign _T_1063 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@147894.4]
  assign _T_1064 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@147897.4]
  assign status_bits_sizeAddr = _T_1063[58:0]; // @[Fringe.scala 158:20:@147876.4 Fringe.scala 163:24:@147895.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_1061}; // @[Fringe.scala 158:20:@147876.4 Fringe.scala 162:28:@147893.4]
  assign _T_1065 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@147898.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@149528.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@149529.4]
  assign _T_1569 = alloc | dealloc; // @[Fringe.scala 204:37:@149530.4]
  assign _T_1573 = _T_1572 ^ _T_1569; // @[package.scala 153:13:@149533.4]
  assign io_rdata = regs_io_rdata; // @[Fringe.scala 125:14:@147822.4]
  assign io_enable = _T_1025 & _T_1029; // @[Fringe.scala 136:13:@147842.4]
  assign io_reset = _T_1030 | reset; // @[Fringe.scala 137:12:@147843.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@147864.4]
  assign io_argIns_1 = regs_io_argIns_3; // @[Fringe.scala 151:51:@147865.4]
  assign io_memStreams_stores_0_cmd_ready = dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 101:72:@142834.4]
  assign io_memStreams_stores_0_data_ready = dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 101:72:@142830.4]
  assign io_memStreams_stores_0_wresp_valid = dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 101:72:@142825.4]
  assign io_memStreams_stores_0_wresp_bits = dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 101:72:@142824.4]
  assign io_dram_0_cmd_valid = dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 195:72:@149026.4]
  assign io_dram_0_cmd_bits_addr = dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@149025.4]
  assign io_dram_0_cmd_bits_size = dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@149024.4]
  assign io_dram_0_cmd_bits_isWr = dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@149022.4]
  assign io_dram_0_cmd_bits_tag = dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@149021.4]
  assign io_dram_0_wdata_valid = dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 195:72:@149019.4]
  assign io_dram_0_wdata_bits_wdata_0 = dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@149003.4]
  assign io_dram_0_wdata_bits_wdata_1 = dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@149004.4]
  assign io_dram_0_wdata_bits_wdata_2 = dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@149005.4]
  assign io_dram_0_wdata_bits_wdata_3 = dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@149006.4]
  assign io_dram_0_wdata_bits_wdata_4 = dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@149007.4]
  assign io_dram_0_wdata_bits_wdata_5 = dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@149008.4]
  assign io_dram_0_wdata_bits_wdata_6 = dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@149009.4]
  assign io_dram_0_wdata_bits_wdata_7 = dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@149010.4]
  assign io_dram_0_wdata_bits_wdata_8 = dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@149011.4]
  assign io_dram_0_wdata_bits_wdata_9 = dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@149012.4]
  assign io_dram_0_wdata_bits_wdata_10 = dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@149013.4]
  assign io_dram_0_wdata_bits_wdata_11 = dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@149014.4]
  assign io_dram_0_wdata_bits_wdata_12 = dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@149015.4]
  assign io_dram_0_wdata_bits_wdata_13 = dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@149016.4]
  assign io_dram_0_wdata_bits_wdata_14 = dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@149017.4]
  assign io_dram_0_wdata_bits_wdata_15 = dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@149018.4]
  assign io_dram_0_wdata_bits_wstrb_0 = dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@148939.4]
  assign io_dram_0_wdata_bits_wstrb_1 = dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@148940.4]
  assign io_dram_0_wdata_bits_wstrb_2 = dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@148941.4]
  assign io_dram_0_wdata_bits_wstrb_3 = dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@148942.4]
  assign io_dram_0_wdata_bits_wstrb_4 = dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@148943.4]
  assign io_dram_0_wdata_bits_wstrb_5 = dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@148944.4]
  assign io_dram_0_wdata_bits_wstrb_6 = dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@148945.4]
  assign io_dram_0_wdata_bits_wstrb_7 = dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@148946.4]
  assign io_dram_0_wdata_bits_wstrb_8 = dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@148947.4]
  assign io_dram_0_wdata_bits_wstrb_9 = dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@148948.4]
  assign io_dram_0_wdata_bits_wstrb_10 = dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@148949.4]
  assign io_dram_0_wdata_bits_wstrb_11 = dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@148950.4]
  assign io_dram_0_wdata_bits_wstrb_12 = dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@148951.4]
  assign io_dram_0_wdata_bits_wstrb_13 = dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@148952.4]
  assign io_dram_0_wdata_bits_wstrb_14 = dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@148953.4]
  assign io_dram_0_wdata_bits_wstrb_15 = dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@148954.4]
  assign io_dram_0_wdata_bits_wstrb_16 = dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@148955.4]
  assign io_dram_0_wdata_bits_wstrb_17 = dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@148956.4]
  assign io_dram_0_wdata_bits_wstrb_18 = dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@148957.4]
  assign io_dram_0_wdata_bits_wstrb_19 = dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@148958.4]
  assign io_dram_0_wdata_bits_wstrb_20 = dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@148959.4]
  assign io_dram_0_wdata_bits_wstrb_21 = dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@148960.4]
  assign io_dram_0_wdata_bits_wstrb_22 = dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@148961.4]
  assign io_dram_0_wdata_bits_wstrb_23 = dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@148962.4]
  assign io_dram_0_wdata_bits_wstrb_24 = dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@148963.4]
  assign io_dram_0_wdata_bits_wstrb_25 = dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@148964.4]
  assign io_dram_0_wdata_bits_wstrb_26 = dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@148965.4]
  assign io_dram_0_wdata_bits_wstrb_27 = dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@148966.4]
  assign io_dram_0_wdata_bits_wstrb_28 = dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@148967.4]
  assign io_dram_0_wdata_bits_wstrb_29 = dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@148968.4]
  assign io_dram_0_wdata_bits_wstrb_30 = dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@148969.4]
  assign io_dram_0_wdata_bits_wstrb_31 = dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@148970.4]
  assign io_dram_0_wdata_bits_wstrb_32 = dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@148971.4]
  assign io_dram_0_wdata_bits_wstrb_33 = dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@148972.4]
  assign io_dram_0_wdata_bits_wstrb_34 = dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@148973.4]
  assign io_dram_0_wdata_bits_wstrb_35 = dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@148974.4]
  assign io_dram_0_wdata_bits_wstrb_36 = dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@148975.4]
  assign io_dram_0_wdata_bits_wstrb_37 = dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@148976.4]
  assign io_dram_0_wdata_bits_wstrb_38 = dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@148977.4]
  assign io_dram_0_wdata_bits_wstrb_39 = dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@148978.4]
  assign io_dram_0_wdata_bits_wstrb_40 = dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@148979.4]
  assign io_dram_0_wdata_bits_wstrb_41 = dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@148980.4]
  assign io_dram_0_wdata_bits_wstrb_42 = dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@148981.4]
  assign io_dram_0_wdata_bits_wstrb_43 = dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@148982.4]
  assign io_dram_0_wdata_bits_wstrb_44 = dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@148983.4]
  assign io_dram_0_wdata_bits_wstrb_45 = dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@148984.4]
  assign io_dram_0_wdata_bits_wstrb_46 = dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@148985.4]
  assign io_dram_0_wdata_bits_wstrb_47 = dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@148986.4]
  assign io_dram_0_wdata_bits_wstrb_48 = dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@148987.4]
  assign io_dram_0_wdata_bits_wstrb_49 = dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@148988.4]
  assign io_dram_0_wdata_bits_wstrb_50 = dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@148989.4]
  assign io_dram_0_wdata_bits_wstrb_51 = dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@148990.4]
  assign io_dram_0_wdata_bits_wstrb_52 = dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@148991.4]
  assign io_dram_0_wdata_bits_wstrb_53 = dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@148992.4]
  assign io_dram_0_wdata_bits_wstrb_54 = dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@148993.4]
  assign io_dram_0_wdata_bits_wstrb_55 = dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@148994.4]
  assign io_dram_0_wdata_bits_wstrb_56 = dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@148995.4]
  assign io_dram_0_wdata_bits_wstrb_57 = dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@148996.4]
  assign io_dram_0_wdata_bits_wstrb_58 = dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@148997.4]
  assign io_dram_0_wdata_bits_wstrb_59 = dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@148998.4]
  assign io_dram_0_wdata_bits_wstrb_60 = dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@148999.4]
  assign io_dram_0_wdata_bits_wstrb_61 = dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@149000.4]
  assign io_dram_0_wdata_bits_wstrb_62 = dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@149001.4]
  assign io_dram_0_wdata_bits_wstrb_63 = dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@149002.4]
  assign io_dram_0_wdata_bits_wlast = dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@148938.4]
  assign io_dram_0_rresp_ready = dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 195:72:@148937.4]
  assign io_dram_0_wresp_ready = dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 195:72:@148918.4]
  assign io_dram_1_cmd_valid = dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 195:72:@149138.4]
  assign io_dram_1_cmd_bits_addr = dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@149137.4]
  assign io_dram_1_cmd_bits_size = dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@149136.4]
  assign io_dram_1_cmd_bits_isWr = dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@149134.4]
  assign io_dram_1_cmd_bits_tag = dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@149133.4]
  assign io_dram_1_wdata_valid = dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 195:72:@149131.4]
  assign io_dram_1_wdata_bits_wdata_0 = dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@149115.4]
  assign io_dram_1_wdata_bits_wdata_1 = dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@149116.4]
  assign io_dram_1_wdata_bits_wdata_2 = dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@149117.4]
  assign io_dram_1_wdata_bits_wdata_3 = dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@149118.4]
  assign io_dram_1_wdata_bits_wdata_4 = dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@149119.4]
  assign io_dram_1_wdata_bits_wdata_5 = dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@149120.4]
  assign io_dram_1_wdata_bits_wdata_6 = dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@149121.4]
  assign io_dram_1_wdata_bits_wdata_7 = dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@149122.4]
  assign io_dram_1_wdata_bits_wdata_8 = dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@149123.4]
  assign io_dram_1_wdata_bits_wdata_9 = dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@149124.4]
  assign io_dram_1_wdata_bits_wdata_10 = dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@149125.4]
  assign io_dram_1_wdata_bits_wdata_11 = dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@149126.4]
  assign io_dram_1_wdata_bits_wdata_12 = dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@149127.4]
  assign io_dram_1_wdata_bits_wdata_13 = dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@149128.4]
  assign io_dram_1_wdata_bits_wdata_14 = dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@149129.4]
  assign io_dram_1_wdata_bits_wdata_15 = dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@149130.4]
  assign io_dram_1_wdata_bits_wstrb_0 = dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@149051.4]
  assign io_dram_1_wdata_bits_wstrb_1 = dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@149052.4]
  assign io_dram_1_wdata_bits_wstrb_2 = dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@149053.4]
  assign io_dram_1_wdata_bits_wstrb_3 = dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@149054.4]
  assign io_dram_1_wdata_bits_wstrb_4 = dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@149055.4]
  assign io_dram_1_wdata_bits_wstrb_5 = dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@149056.4]
  assign io_dram_1_wdata_bits_wstrb_6 = dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@149057.4]
  assign io_dram_1_wdata_bits_wstrb_7 = dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@149058.4]
  assign io_dram_1_wdata_bits_wstrb_8 = dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@149059.4]
  assign io_dram_1_wdata_bits_wstrb_9 = dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@149060.4]
  assign io_dram_1_wdata_bits_wstrb_10 = dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@149061.4]
  assign io_dram_1_wdata_bits_wstrb_11 = dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@149062.4]
  assign io_dram_1_wdata_bits_wstrb_12 = dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@149063.4]
  assign io_dram_1_wdata_bits_wstrb_13 = dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@149064.4]
  assign io_dram_1_wdata_bits_wstrb_14 = dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@149065.4]
  assign io_dram_1_wdata_bits_wstrb_15 = dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@149066.4]
  assign io_dram_1_wdata_bits_wstrb_16 = dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@149067.4]
  assign io_dram_1_wdata_bits_wstrb_17 = dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@149068.4]
  assign io_dram_1_wdata_bits_wstrb_18 = dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@149069.4]
  assign io_dram_1_wdata_bits_wstrb_19 = dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@149070.4]
  assign io_dram_1_wdata_bits_wstrb_20 = dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@149071.4]
  assign io_dram_1_wdata_bits_wstrb_21 = dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@149072.4]
  assign io_dram_1_wdata_bits_wstrb_22 = dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@149073.4]
  assign io_dram_1_wdata_bits_wstrb_23 = dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@149074.4]
  assign io_dram_1_wdata_bits_wstrb_24 = dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@149075.4]
  assign io_dram_1_wdata_bits_wstrb_25 = dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@149076.4]
  assign io_dram_1_wdata_bits_wstrb_26 = dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@149077.4]
  assign io_dram_1_wdata_bits_wstrb_27 = dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@149078.4]
  assign io_dram_1_wdata_bits_wstrb_28 = dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@149079.4]
  assign io_dram_1_wdata_bits_wstrb_29 = dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@149080.4]
  assign io_dram_1_wdata_bits_wstrb_30 = dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@149081.4]
  assign io_dram_1_wdata_bits_wstrb_31 = dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@149082.4]
  assign io_dram_1_wdata_bits_wstrb_32 = dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@149083.4]
  assign io_dram_1_wdata_bits_wstrb_33 = dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@149084.4]
  assign io_dram_1_wdata_bits_wstrb_34 = dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@149085.4]
  assign io_dram_1_wdata_bits_wstrb_35 = dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@149086.4]
  assign io_dram_1_wdata_bits_wstrb_36 = dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@149087.4]
  assign io_dram_1_wdata_bits_wstrb_37 = dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@149088.4]
  assign io_dram_1_wdata_bits_wstrb_38 = dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@149089.4]
  assign io_dram_1_wdata_bits_wstrb_39 = dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@149090.4]
  assign io_dram_1_wdata_bits_wstrb_40 = dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@149091.4]
  assign io_dram_1_wdata_bits_wstrb_41 = dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@149092.4]
  assign io_dram_1_wdata_bits_wstrb_42 = dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@149093.4]
  assign io_dram_1_wdata_bits_wstrb_43 = dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@149094.4]
  assign io_dram_1_wdata_bits_wstrb_44 = dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@149095.4]
  assign io_dram_1_wdata_bits_wstrb_45 = dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@149096.4]
  assign io_dram_1_wdata_bits_wstrb_46 = dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@149097.4]
  assign io_dram_1_wdata_bits_wstrb_47 = dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@149098.4]
  assign io_dram_1_wdata_bits_wstrb_48 = dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@149099.4]
  assign io_dram_1_wdata_bits_wstrb_49 = dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@149100.4]
  assign io_dram_1_wdata_bits_wstrb_50 = dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@149101.4]
  assign io_dram_1_wdata_bits_wstrb_51 = dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@149102.4]
  assign io_dram_1_wdata_bits_wstrb_52 = dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@149103.4]
  assign io_dram_1_wdata_bits_wstrb_53 = dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@149104.4]
  assign io_dram_1_wdata_bits_wstrb_54 = dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@149105.4]
  assign io_dram_1_wdata_bits_wstrb_55 = dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@149106.4]
  assign io_dram_1_wdata_bits_wstrb_56 = dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@149107.4]
  assign io_dram_1_wdata_bits_wstrb_57 = dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@149108.4]
  assign io_dram_1_wdata_bits_wstrb_58 = dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@149109.4]
  assign io_dram_1_wdata_bits_wstrb_59 = dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@149110.4]
  assign io_dram_1_wdata_bits_wstrb_60 = dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@149111.4]
  assign io_dram_1_wdata_bits_wstrb_61 = dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@149112.4]
  assign io_dram_1_wdata_bits_wstrb_62 = dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@149113.4]
  assign io_dram_1_wdata_bits_wstrb_63 = dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@149114.4]
  assign io_dram_1_wdata_bits_wlast = dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@149050.4]
  assign io_dram_1_rresp_ready = dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 195:72:@149049.4]
  assign io_dram_1_wresp_ready = dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 195:72:@149030.4]
  assign io_dram_2_cmd_valid = dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 195:72:@149250.4]
  assign io_dram_2_cmd_bits_addr = dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@149249.4]
  assign io_dram_2_cmd_bits_size = dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@149248.4]
  assign io_dram_2_cmd_bits_isWr = dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@149246.4]
  assign io_dram_2_cmd_bits_tag = dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@149245.4]
  assign io_dram_2_wdata_valid = dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 195:72:@149243.4]
  assign io_dram_2_wdata_bits_wdata_0 = dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@149227.4]
  assign io_dram_2_wdata_bits_wdata_1 = dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@149228.4]
  assign io_dram_2_wdata_bits_wdata_2 = dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@149229.4]
  assign io_dram_2_wdata_bits_wdata_3 = dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@149230.4]
  assign io_dram_2_wdata_bits_wdata_4 = dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@149231.4]
  assign io_dram_2_wdata_bits_wdata_5 = dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@149232.4]
  assign io_dram_2_wdata_bits_wdata_6 = dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@149233.4]
  assign io_dram_2_wdata_bits_wdata_7 = dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@149234.4]
  assign io_dram_2_wdata_bits_wdata_8 = dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@149235.4]
  assign io_dram_2_wdata_bits_wdata_9 = dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@149236.4]
  assign io_dram_2_wdata_bits_wdata_10 = dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@149237.4]
  assign io_dram_2_wdata_bits_wdata_11 = dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@149238.4]
  assign io_dram_2_wdata_bits_wdata_12 = dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@149239.4]
  assign io_dram_2_wdata_bits_wdata_13 = dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@149240.4]
  assign io_dram_2_wdata_bits_wdata_14 = dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@149241.4]
  assign io_dram_2_wdata_bits_wdata_15 = dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@149242.4]
  assign io_dram_2_wdata_bits_wstrb_0 = dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@149163.4]
  assign io_dram_2_wdata_bits_wstrb_1 = dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@149164.4]
  assign io_dram_2_wdata_bits_wstrb_2 = dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@149165.4]
  assign io_dram_2_wdata_bits_wstrb_3 = dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@149166.4]
  assign io_dram_2_wdata_bits_wstrb_4 = dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@149167.4]
  assign io_dram_2_wdata_bits_wstrb_5 = dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@149168.4]
  assign io_dram_2_wdata_bits_wstrb_6 = dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@149169.4]
  assign io_dram_2_wdata_bits_wstrb_7 = dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@149170.4]
  assign io_dram_2_wdata_bits_wstrb_8 = dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@149171.4]
  assign io_dram_2_wdata_bits_wstrb_9 = dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@149172.4]
  assign io_dram_2_wdata_bits_wstrb_10 = dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@149173.4]
  assign io_dram_2_wdata_bits_wstrb_11 = dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@149174.4]
  assign io_dram_2_wdata_bits_wstrb_12 = dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@149175.4]
  assign io_dram_2_wdata_bits_wstrb_13 = dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@149176.4]
  assign io_dram_2_wdata_bits_wstrb_14 = dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@149177.4]
  assign io_dram_2_wdata_bits_wstrb_15 = dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@149178.4]
  assign io_dram_2_wdata_bits_wstrb_16 = dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@149179.4]
  assign io_dram_2_wdata_bits_wstrb_17 = dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@149180.4]
  assign io_dram_2_wdata_bits_wstrb_18 = dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@149181.4]
  assign io_dram_2_wdata_bits_wstrb_19 = dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@149182.4]
  assign io_dram_2_wdata_bits_wstrb_20 = dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@149183.4]
  assign io_dram_2_wdata_bits_wstrb_21 = dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@149184.4]
  assign io_dram_2_wdata_bits_wstrb_22 = dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@149185.4]
  assign io_dram_2_wdata_bits_wstrb_23 = dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@149186.4]
  assign io_dram_2_wdata_bits_wstrb_24 = dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@149187.4]
  assign io_dram_2_wdata_bits_wstrb_25 = dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@149188.4]
  assign io_dram_2_wdata_bits_wstrb_26 = dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@149189.4]
  assign io_dram_2_wdata_bits_wstrb_27 = dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@149190.4]
  assign io_dram_2_wdata_bits_wstrb_28 = dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@149191.4]
  assign io_dram_2_wdata_bits_wstrb_29 = dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@149192.4]
  assign io_dram_2_wdata_bits_wstrb_30 = dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@149193.4]
  assign io_dram_2_wdata_bits_wstrb_31 = dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@149194.4]
  assign io_dram_2_wdata_bits_wstrb_32 = dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@149195.4]
  assign io_dram_2_wdata_bits_wstrb_33 = dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@149196.4]
  assign io_dram_2_wdata_bits_wstrb_34 = dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@149197.4]
  assign io_dram_2_wdata_bits_wstrb_35 = dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@149198.4]
  assign io_dram_2_wdata_bits_wstrb_36 = dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@149199.4]
  assign io_dram_2_wdata_bits_wstrb_37 = dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@149200.4]
  assign io_dram_2_wdata_bits_wstrb_38 = dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@149201.4]
  assign io_dram_2_wdata_bits_wstrb_39 = dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@149202.4]
  assign io_dram_2_wdata_bits_wstrb_40 = dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@149203.4]
  assign io_dram_2_wdata_bits_wstrb_41 = dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@149204.4]
  assign io_dram_2_wdata_bits_wstrb_42 = dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@149205.4]
  assign io_dram_2_wdata_bits_wstrb_43 = dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@149206.4]
  assign io_dram_2_wdata_bits_wstrb_44 = dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@149207.4]
  assign io_dram_2_wdata_bits_wstrb_45 = dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@149208.4]
  assign io_dram_2_wdata_bits_wstrb_46 = dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@149209.4]
  assign io_dram_2_wdata_bits_wstrb_47 = dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@149210.4]
  assign io_dram_2_wdata_bits_wstrb_48 = dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@149211.4]
  assign io_dram_2_wdata_bits_wstrb_49 = dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@149212.4]
  assign io_dram_2_wdata_bits_wstrb_50 = dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@149213.4]
  assign io_dram_2_wdata_bits_wstrb_51 = dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@149214.4]
  assign io_dram_2_wdata_bits_wstrb_52 = dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@149215.4]
  assign io_dram_2_wdata_bits_wstrb_53 = dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@149216.4]
  assign io_dram_2_wdata_bits_wstrb_54 = dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@149217.4]
  assign io_dram_2_wdata_bits_wstrb_55 = dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@149218.4]
  assign io_dram_2_wdata_bits_wstrb_56 = dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@149219.4]
  assign io_dram_2_wdata_bits_wstrb_57 = dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@149220.4]
  assign io_dram_2_wdata_bits_wstrb_58 = dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@149221.4]
  assign io_dram_2_wdata_bits_wstrb_59 = dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@149222.4]
  assign io_dram_2_wdata_bits_wstrb_60 = dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@149223.4]
  assign io_dram_2_wdata_bits_wstrb_61 = dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@149224.4]
  assign io_dram_2_wdata_bits_wstrb_62 = dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@149225.4]
  assign io_dram_2_wdata_bits_wstrb_63 = dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@149226.4]
  assign io_dram_2_wdata_bits_wlast = dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@149162.4]
  assign io_dram_2_rresp_ready = dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 195:72:@149161.4]
  assign io_dram_2_wresp_ready = dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 195:72:@149142.4]
  assign io_dram_3_cmd_valid = dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 195:72:@149362.4]
  assign io_dram_3_cmd_bits_addr = dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@149361.4]
  assign io_dram_3_cmd_bits_size = dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@149360.4]
  assign io_dram_3_cmd_bits_isWr = dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@149358.4]
  assign io_dram_3_cmd_bits_tag = dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@149357.4]
  assign io_dram_3_wdata_valid = dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 195:72:@149355.4]
  assign io_dram_3_wdata_bits_wdata_0 = dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@149339.4]
  assign io_dram_3_wdata_bits_wdata_1 = dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@149340.4]
  assign io_dram_3_wdata_bits_wdata_2 = dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@149341.4]
  assign io_dram_3_wdata_bits_wdata_3 = dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@149342.4]
  assign io_dram_3_wdata_bits_wdata_4 = dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@149343.4]
  assign io_dram_3_wdata_bits_wdata_5 = dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@149344.4]
  assign io_dram_3_wdata_bits_wdata_6 = dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@149345.4]
  assign io_dram_3_wdata_bits_wdata_7 = dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@149346.4]
  assign io_dram_3_wdata_bits_wdata_8 = dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@149347.4]
  assign io_dram_3_wdata_bits_wdata_9 = dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@149348.4]
  assign io_dram_3_wdata_bits_wdata_10 = dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@149349.4]
  assign io_dram_3_wdata_bits_wdata_11 = dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@149350.4]
  assign io_dram_3_wdata_bits_wdata_12 = dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@149351.4]
  assign io_dram_3_wdata_bits_wdata_13 = dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@149352.4]
  assign io_dram_3_wdata_bits_wdata_14 = dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@149353.4]
  assign io_dram_3_wdata_bits_wdata_15 = dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@149354.4]
  assign io_dram_3_wdata_bits_wstrb_0 = dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@149275.4]
  assign io_dram_3_wdata_bits_wstrb_1 = dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@149276.4]
  assign io_dram_3_wdata_bits_wstrb_2 = dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@149277.4]
  assign io_dram_3_wdata_bits_wstrb_3 = dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@149278.4]
  assign io_dram_3_wdata_bits_wstrb_4 = dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@149279.4]
  assign io_dram_3_wdata_bits_wstrb_5 = dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@149280.4]
  assign io_dram_3_wdata_bits_wstrb_6 = dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@149281.4]
  assign io_dram_3_wdata_bits_wstrb_7 = dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@149282.4]
  assign io_dram_3_wdata_bits_wstrb_8 = dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@149283.4]
  assign io_dram_3_wdata_bits_wstrb_9 = dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@149284.4]
  assign io_dram_3_wdata_bits_wstrb_10 = dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@149285.4]
  assign io_dram_3_wdata_bits_wstrb_11 = dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@149286.4]
  assign io_dram_3_wdata_bits_wstrb_12 = dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@149287.4]
  assign io_dram_3_wdata_bits_wstrb_13 = dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@149288.4]
  assign io_dram_3_wdata_bits_wstrb_14 = dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@149289.4]
  assign io_dram_3_wdata_bits_wstrb_15 = dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@149290.4]
  assign io_dram_3_wdata_bits_wstrb_16 = dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@149291.4]
  assign io_dram_3_wdata_bits_wstrb_17 = dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@149292.4]
  assign io_dram_3_wdata_bits_wstrb_18 = dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@149293.4]
  assign io_dram_3_wdata_bits_wstrb_19 = dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@149294.4]
  assign io_dram_3_wdata_bits_wstrb_20 = dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@149295.4]
  assign io_dram_3_wdata_bits_wstrb_21 = dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@149296.4]
  assign io_dram_3_wdata_bits_wstrb_22 = dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@149297.4]
  assign io_dram_3_wdata_bits_wstrb_23 = dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@149298.4]
  assign io_dram_3_wdata_bits_wstrb_24 = dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@149299.4]
  assign io_dram_3_wdata_bits_wstrb_25 = dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@149300.4]
  assign io_dram_3_wdata_bits_wstrb_26 = dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@149301.4]
  assign io_dram_3_wdata_bits_wstrb_27 = dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@149302.4]
  assign io_dram_3_wdata_bits_wstrb_28 = dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@149303.4]
  assign io_dram_3_wdata_bits_wstrb_29 = dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@149304.4]
  assign io_dram_3_wdata_bits_wstrb_30 = dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@149305.4]
  assign io_dram_3_wdata_bits_wstrb_31 = dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@149306.4]
  assign io_dram_3_wdata_bits_wstrb_32 = dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@149307.4]
  assign io_dram_3_wdata_bits_wstrb_33 = dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@149308.4]
  assign io_dram_3_wdata_bits_wstrb_34 = dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@149309.4]
  assign io_dram_3_wdata_bits_wstrb_35 = dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@149310.4]
  assign io_dram_3_wdata_bits_wstrb_36 = dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@149311.4]
  assign io_dram_3_wdata_bits_wstrb_37 = dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@149312.4]
  assign io_dram_3_wdata_bits_wstrb_38 = dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@149313.4]
  assign io_dram_3_wdata_bits_wstrb_39 = dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@149314.4]
  assign io_dram_3_wdata_bits_wstrb_40 = dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@149315.4]
  assign io_dram_3_wdata_bits_wstrb_41 = dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@149316.4]
  assign io_dram_3_wdata_bits_wstrb_42 = dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@149317.4]
  assign io_dram_3_wdata_bits_wstrb_43 = dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@149318.4]
  assign io_dram_3_wdata_bits_wstrb_44 = dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@149319.4]
  assign io_dram_3_wdata_bits_wstrb_45 = dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@149320.4]
  assign io_dram_3_wdata_bits_wstrb_46 = dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@149321.4]
  assign io_dram_3_wdata_bits_wstrb_47 = dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@149322.4]
  assign io_dram_3_wdata_bits_wstrb_48 = dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@149323.4]
  assign io_dram_3_wdata_bits_wstrb_49 = dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@149324.4]
  assign io_dram_3_wdata_bits_wstrb_50 = dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@149325.4]
  assign io_dram_3_wdata_bits_wstrb_51 = dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@149326.4]
  assign io_dram_3_wdata_bits_wstrb_52 = dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@149327.4]
  assign io_dram_3_wdata_bits_wstrb_53 = dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@149328.4]
  assign io_dram_3_wdata_bits_wstrb_54 = dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@149329.4]
  assign io_dram_3_wdata_bits_wstrb_55 = dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@149330.4]
  assign io_dram_3_wdata_bits_wstrb_56 = dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@149331.4]
  assign io_dram_3_wdata_bits_wstrb_57 = dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@149332.4]
  assign io_dram_3_wdata_bits_wstrb_58 = dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@149333.4]
  assign io_dram_3_wdata_bits_wstrb_59 = dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@149334.4]
  assign io_dram_3_wdata_bits_wstrb_60 = dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@149335.4]
  assign io_dram_3_wdata_bits_wstrb_61 = dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@149336.4]
  assign io_dram_3_wdata_bits_wstrb_62 = dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@149337.4]
  assign io_dram_3_wdata_bits_wstrb_63 = dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@149338.4]
  assign io_dram_3_wdata_bits_wlast = dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@149274.4]
  assign io_dram_3_rresp_ready = dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 195:72:@149273.4]
  assign io_dram_3_wresp_ready = dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 195:72:@149254.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@145793.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@145792.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@145791.4]
  assign dramArbs_0_clock = clock; // @[:@141916.4]
  assign dramArbs_0_reset = _T_1030 | reset; // @[:@141917.4 Fringe.scala 187:30:@148908.4]
  assign dramArbs_0_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@148912.4]
  assign dramArbs_0_io_app_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[Fringe.scala 101:72:@142833.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[Fringe.scala 101:72:@142832.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[Fringe.scala 101:72:@142831.4]
  assign dramArbs_0_io_app_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[Fringe.scala 101:72:@142829.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[Fringe.scala 101:72:@142828.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[Fringe.scala 101:72:@142827.4]
  assign dramArbs_0_io_app_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[Fringe.scala 101:72:@142826.4]
  assign dramArbs_0_io_dram_cmd_ready = io_dram_0_cmd_ready; // @[Fringe.scala 195:72:@149027.4]
  assign dramArbs_0_io_dram_wdata_ready = io_dram_0_wdata_ready; // @[Fringe.scala 195:72:@149020.4]
  assign dramArbs_0_io_dram_wresp_valid = io_dram_0_wresp_valid; // @[Fringe.scala 195:72:@148917.4]
  assign dramArbs_0_io_dram_wresp_bits_tag = io_dram_0_wresp_bits_tag; // @[Fringe.scala 195:72:@148916.4]
  assign dramArbs_1_clock = clock; // @[:@142909.4]
  assign dramArbs_1_reset = _T_1030 | reset; // @[:@142910.4 Fringe.scala 187:30:@148909.4]
  assign dramArbs_1_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@148913.4]
  assign dramArbs_1_io_dram_cmd_ready = io_dram_1_cmd_ready; // @[Fringe.scala 195:72:@149139.4]
  assign dramArbs_1_io_dram_wdata_ready = io_dram_1_wdata_ready; // @[Fringe.scala 195:72:@149132.4]
  assign dramArbs_1_io_dram_wresp_valid = io_dram_1_wresp_valid; // @[Fringe.scala 195:72:@149029.4]
  assign dramArbs_1_io_dram_wresp_bits_tag = io_dram_1_wresp_bits_tag; // @[Fringe.scala 195:72:@149028.4]
  assign dramArbs_2_clock = clock; // @[:@143869.4]
  assign dramArbs_2_reset = _T_1030 | reset; // @[:@143870.4 Fringe.scala 187:30:@148910.4]
  assign dramArbs_2_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@148914.4]
  assign dramArbs_2_io_dram_cmd_ready = io_dram_2_cmd_ready; // @[Fringe.scala 195:72:@149251.4]
  assign dramArbs_2_io_dram_wdata_ready = io_dram_2_wdata_ready; // @[Fringe.scala 195:72:@149244.4]
  assign dramArbs_2_io_dram_wresp_valid = io_dram_2_wresp_valid; // @[Fringe.scala 195:72:@149141.4]
  assign dramArbs_2_io_dram_wresp_bits_tag = io_dram_2_wresp_bits_tag; // @[Fringe.scala 195:72:@149140.4]
  assign dramArbs_3_clock = clock; // @[:@144829.4]
  assign dramArbs_3_reset = _T_1030 | reset; // @[:@144830.4 Fringe.scala 187:30:@148911.4]
  assign dramArbs_3_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@148915.4]
  assign dramArbs_3_io_dram_cmd_ready = io_dram_3_cmd_ready; // @[Fringe.scala 195:72:@149363.4]
  assign dramArbs_3_io_dram_wdata_ready = io_dram_3_wdata_ready; // @[Fringe.scala 195:72:@149356.4]
  assign dramArbs_3_io_dram_wresp_valid = io_dram_3_wresp_valid; // @[Fringe.scala 195:72:@149253.4]
  assign dramArbs_3_io_dram_wresp_bits_tag = io_dram_3_wresp_bits_tag; // @[Fringe.scala 195:72:@149252.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@145796.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@145795.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@145794.4]
  assign heap_io_host_0_resp_valid = _T_1569 & _T_1573; // @[Fringe.scala 204:22:@149535.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@149536.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@149537.4]
  assign regs_clock = clock; // @[:@145798.4]
  assign regs_reset = reset; // @[:@145799.4 Fringe.scala 139:14:@147846.4]
  assign regs_io_raddr = io_raddr; // @[Fringe.scala 118:17:@147818.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@147820.4]
  assign regs_io_waddr = io_waddr; // @[Fringe.scala 119:17:@147819.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@147821.4]
  assign regs_io_reset = _T_1030 | reset; // @[Fringe.scala 138:17:@147844.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_1049; // @[Fringe.scala 170:23:@147896.4]
  assign regs_io_argOuts_0_bits = {_T_1065,_T_1064}; // @[Fringe.scala 171:22:@147900.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@147903.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@147902.4]
  assign timeoutCtr_clock = clock; // @[:@147848.4]
  assign timeoutCtr_reset = reset; // @[:@147849.4]
  assign timeoutCtr_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 149:24:@147863.4]
  assign depulser_clock = clock; // @[:@147867.4]
  assign depulser_reset = reset; // @[:@147868.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@147873.4]
  assign depulser_io_rst = _T_1040[0]; // @[Fringe.scala 156:19:@147875.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1047 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1572 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1047 <= 1'h0;
    end else begin
      _T_1047 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1572 <= 1'h0;
    end else begin
      _T_1572 <= _T_1569;
    end
  end
endmodule
module AXI4LiteToRFBridge( // @[:@149552.2]
  input         clock, // @[:@149553.4]
  input         reset, // @[:@149554.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@149555.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@149555.4]
  input         io_S_AXI_AWVALID, // @[:@149555.4]
  output        io_S_AXI_AWREADY, // @[:@149555.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@149555.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@149555.4]
  input         io_S_AXI_ARVALID, // @[:@149555.4]
  output        io_S_AXI_ARREADY, // @[:@149555.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@149555.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@149555.4]
  input         io_S_AXI_WVALID, // @[:@149555.4]
  output        io_S_AXI_WREADY, // @[:@149555.4]
  output [31:0] io_S_AXI_RDATA, // @[:@149555.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@149555.4]
  output        io_S_AXI_RVALID, // @[:@149555.4]
  input         io_S_AXI_RREADY, // @[:@149555.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@149555.4]
  output        io_S_AXI_BVALID, // @[:@149555.4]
  input         io_S_AXI_BREADY, // @[:@149555.4]
  output [31:0] io_raddr, // @[:@149555.4]
  output        io_wen, // @[:@149555.4]
  output [31:0] io_waddr, // @[:@149555.4]
  output [31:0] io_wdata, // @[:@149555.4]
  input  [31:0] io_rdata // @[:@149555.4]
);
  wire [31:0] d_rf_rdata; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire [31:0] d_rf_wdata; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire [31:0] d_rf_waddr; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire  d_rf_wen; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire [31:0] d_rf_raddr; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire  d_S_AXI_ARESETN; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire  d_S_AXI_ACLK; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire [31:0] d_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire [2:0] d_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire  d_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire  d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire [31:0] d_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire [2:0] d_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire  d_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire  d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire [31:0] d_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire [3:0] d_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire  d_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire  d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire [31:0] d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire [1:0] d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire  d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire  d_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire [1:0] d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire  d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  wire  d_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
  AXI4LiteToRFBridgeVerilog d ( // @[AXI4LiteToRFBridge.scala 36:17:@149557.4]
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 38:14:@149581.4]
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 38:14:@149577.4]
  assign io_S_AXI_WREADY = d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 38:14:@149573.4]
  assign io_S_AXI_RDATA = d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 38:14:@149572.4]
  assign io_S_AXI_RRESP = d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 38:14:@149571.4]
  assign io_S_AXI_RVALID = d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 38:14:@149570.4]
  assign io_S_AXI_BRESP = d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 38:14:@149568.4]
  assign io_S_AXI_BVALID = d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 38:14:@149567.4]
  assign io_raddr = d_rf_raddr; // @[AXI4LiteToRFBridge.scala 42:12:@149589.4]
  assign io_wen = d_rf_wen; // @[AXI4LiteToRFBridge.scala 45:12:@149592.4]
  assign io_waddr = d_rf_waddr; // @[AXI4LiteToRFBridge.scala 43:12:@149590.4]
  assign io_wdata = d_rf_wdata; // @[AXI4LiteToRFBridge.scala 44:12:@149591.4]
  assign d_rf_rdata = io_rdata; // @[AXI4LiteToRFBridge.scala 46:17:@149593.4]
  assign d_S_AXI_ARESETN = ~ reset; // @[AXI4LiteToRFBridge.scala 40:22:@149588.4]
  assign d_S_AXI_ACLK = clock; // @[AXI4LiteToRFBridge.scala 39:19:@149585.4]
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 38:14:@149584.4]
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 38:14:@149583.4]
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 38:14:@149582.4]
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 38:14:@149580.4]
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 38:14:@149579.4]
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 38:14:@149578.4]
  assign d_S_AXI_WDATA = io_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 38:14:@149576.4]
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 38:14:@149575.4]
  assign d_S_AXI_WVALID = io_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 38:14:@149574.4]
  assign d_S_AXI_RREADY = io_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 38:14:@149569.4]
  assign d_S_AXI_BREADY = io_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 38:14:@149566.4]
endmodule
module MAGToAXI4Bridge( // @[:@149595.2]
  output         io_in_cmd_ready, // @[:@149598.4]
  input          io_in_cmd_valid, // @[:@149598.4]
  input  [63:0]  io_in_cmd_bits_addr, // @[:@149598.4]
  input  [31:0]  io_in_cmd_bits_size, // @[:@149598.4]
  input          io_in_cmd_bits_isWr, // @[:@149598.4]
  input  [31:0]  io_in_cmd_bits_tag, // @[:@149598.4]
  output         io_in_wdata_ready, // @[:@149598.4]
  input          io_in_wdata_valid, // @[:@149598.4]
  input  [31:0]  io_in_wdata_bits_wdata_0, // @[:@149598.4]
  input  [31:0]  io_in_wdata_bits_wdata_1, // @[:@149598.4]
  input  [31:0]  io_in_wdata_bits_wdata_2, // @[:@149598.4]
  input  [31:0]  io_in_wdata_bits_wdata_3, // @[:@149598.4]
  input  [31:0]  io_in_wdata_bits_wdata_4, // @[:@149598.4]
  input  [31:0]  io_in_wdata_bits_wdata_5, // @[:@149598.4]
  input  [31:0]  io_in_wdata_bits_wdata_6, // @[:@149598.4]
  input  [31:0]  io_in_wdata_bits_wdata_7, // @[:@149598.4]
  input  [31:0]  io_in_wdata_bits_wdata_8, // @[:@149598.4]
  input  [31:0]  io_in_wdata_bits_wdata_9, // @[:@149598.4]
  input  [31:0]  io_in_wdata_bits_wdata_10, // @[:@149598.4]
  input  [31:0]  io_in_wdata_bits_wdata_11, // @[:@149598.4]
  input  [31:0]  io_in_wdata_bits_wdata_12, // @[:@149598.4]
  input  [31:0]  io_in_wdata_bits_wdata_13, // @[:@149598.4]
  input  [31:0]  io_in_wdata_bits_wdata_14, // @[:@149598.4]
  input  [31:0]  io_in_wdata_bits_wdata_15, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_0, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_1, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_2, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_3, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_4, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_5, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_6, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_7, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_8, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_9, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_10, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_11, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_12, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_13, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_14, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_15, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_16, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_17, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_18, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_19, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_20, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_21, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_22, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_23, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_24, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_25, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_26, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_27, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_28, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_29, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_30, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_31, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_32, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_33, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_34, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_35, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_36, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_37, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_38, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_39, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_40, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_41, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_42, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_43, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_44, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_45, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_46, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_47, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_48, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_49, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_50, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_51, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_52, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_53, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_54, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_55, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_56, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_57, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_58, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_59, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_60, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_61, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_62, // @[:@149598.4]
  input          io_in_wdata_bits_wstrb_63, // @[:@149598.4]
  input          io_in_wdata_bits_wlast, // @[:@149598.4]
  input          io_in_rresp_ready, // @[:@149598.4]
  input          io_in_wresp_ready, // @[:@149598.4]
  output         io_in_wresp_valid, // @[:@149598.4]
  output [31:0]  io_in_wresp_bits_tag, // @[:@149598.4]
  output [31:0]  io_M_AXI_AWID, // @[:@149598.4]
  output [31:0]  io_M_AXI_AWADDR, // @[:@149598.4]
  output [7:0]   io_M_AXI_AWLEN, // @[:@149598.4]
  output         io_M_AXI_AWVALID, // @[:@149598.4]
  input          io_M_AXI_AWREADY, // @[:@149598.4]
  output [31:0]  io_M_AXI_ARID, // @[:@149598.4]
  output [31:0]  io_M_AXI_ARADDR, // @[:@149598.4]
  output [7:0]   io_M_AXI_ARLEN, // @[:@149598.4]
  output         io_M_AXI_ARVALID, // @[:@149598.4]
  input          io_M_AXI_ARREADY, // @[:@149598.4]
  output [511:0] io_M_AXI_WDATA, // @[:@149598.4]
  output [63:0]  io_M_AXI_WSTRB, // @[:@149598.4]
  output         io_M_AXI_WLAST, // @[:@149598.4]
  output         io_M_AXI_WVALID, // @[:@149598.4]
  input          io_M_AXI_WREADY, // @[:@149598.4]
  output         io_M_AXI_RREADY, // @[:@149598.4]
  input  [31:0]  io_M_AXI_BID, // @[:@149598.4]
  input          io_M_AXI_BVALID, // @[:@149598.4]
  output         io_M_AXI_BREADY // @[:@149598.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@149755.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@149756.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@149757.4]
  wire  _T_228; // @[MAGToAXI4Bridge.scala 35:42:@149765.4]
  wire [319:0] _T_250; // @[Cat.scala 30:58:@149792.4]
  wire [479:0] _T_255; // @[Cat.scala 30:58:@149797.4]
  wire [9:0] _T_265; // @[Cat.scala 30:58:@149808.4]
  wire [18:0] _T_274; // @[Cat.scala 30:58:@149817.4]
  wire [27:0] _T_283; // @[Cat.scala 30:58:@149826.4]
  wire [36:0] _T_292; // @[Cat.scala 30:58:@149835.4]
  wire [45:0] _T_301; // @[Cat.scala 30:58:@149844.4]
  wire [54:0] _T_310; // @[Cat.scala 30:58:@149853.4]
  wire [62:0] _T_318; // @[Cat.scala 30:58:@149861.4]
  assign _T_218 = io_in_cmd_bits_size - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@149755.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@149756.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@149757.4]
  assign _T_228 = io_in_cmd_bits_isWr == 1'h0; // @[MAGToAXI4Bridge.scala 35:42:@149765.4]
  assign _T_250 = {io_in_wdata_bits_wdata_15,io_in_wdata_bits_wdata_14,io_in_wdata_bits_wdata_13,io_in_wdata_bits_wdata_12,io_in_wdata_bits_wdata_11,io_in_wdata_bits_wdata_10,io_in_wdata_bits_wdata_9,io_in_wdata_bits_wdata_8,io_in_wdata_bits_wdata_7,io_in_wdata_bits_wdata_6}; // @[Cat.scala 30:58:@149792.4]
  assign _T_255 = {_T_250,io_in_wdata_bits_wdata_5,io_in_wdata_bits_wdata_4,io_in_wdata_bits_wdata_3,io_in_wdata_bits_wdata_2,io_in_wdata_bits_wdata_1}; // @[Cat.scala 30:58:@149797.4]
  assign _T_265 = {io_in_wdata_bits_wstrb_63,io_in_wdata_bits_wstrb_62,io_in_wdata_bits_wstrb_61,io_in_wdata_bits_wstrb_60,io_in_wdata_bits_wstrb_59,io_in_wdata_bits_wstrb_58,io_in_wdata_bits_wstrb_57,io_in_wdata_bits_wstrb_56,io_in_wdata_bits_wstrb_55,io_in_wdata_bits_wstrb_54}; // @[Cat.scala 30:58:@149808.4]
  assign _T_274 = {_T_265,io_in_wdata_bits_wstrb_53,io_in_wdata_bits_wstrb_52,io_in_wdata_bits_wstrb_51,io_in_wdata_bits_wstrb_50,io_in_wdata_bits_wstrb_49,io_in_wdata_bits_wstrb_48,io_in_wdata_bits_wstrb_47,io_in_wdata_bits_wstrb_46,io_in_wdata_bits_wstrb_45}; // @[Cat.scala 30:58:@149817.4]
  assign _T_283 = {_T_274,io_in_wdata_bits_wstrb_44,io_in_wdata_bits_wstrb_43,io_in_wdata_bits_wstrb_42,io_in_wdata_bits_wstrb_41,io_in_wdata_bits_wstrb_40,io_in_wdata_bits_wstrb_39,io_in_wdata_bits_wstrb_38,io_in_wdata_bits_wstrb_37,io_in_wdata_bits_wstrb_36}; // @[Cat.scala 30:58:@149826.4]
  assign _T_292 = {_T_283,io_in_wdata_bits_wstrb_35,io_in_wdata_bits_wstrb_34,io_in_wdata_bits_wstrb_33,io_in_wdata_bits_wstrb_32,io_in_wdata_bits_wstrb_31,io_in_wdata_bits_wstrb_30,io_in_wdata_bits_wstrb_29,io_in_wdata_bits_wstrb_28,io_in_wdata_bits_wstrb_27}; // @[Cat.scala 30:58:@149835.4]
  assign _T_301 = {_T_292,io_in_wdata_bits_wstrb_26,io_in_wdata_bits_wstrb_25,io_in_wdata_bits_wstrb_24,io_in_wdata_bits_wstrb_23,io_in_wdata_bits_wstrb_22,io_in_wdata_bits_wstrb_21,io_in_wdata_bits_wstrb_20,io_in_wdata_bits_wstrb_19,io_in_wdata_bits_wstrb_18}; // @[Cat.scala 30:58:@149844.4]
  assign _T_310 = {_T_301,io_in_wdata_bits_wstrb_17,io_in_wdata_bits_wstrb_16,io_in_wdata_bits_wstrb_15,io_in_wdata_bits_wstrb_14,io_in_wdata_bits_wstrb_13,io_in_wdata_bits_wstrb_12,io_in_wdata_bits_wstrb_11,io_in_wdata_bits_wstrb_10,io_in_wdata_bits_wstrb_9}; // @[Cat.scala 30:58:@149853.4]
  assign _T_318 = {_T_310,io_in_wdata_bits_wstrb_8,io_in_wdata_bits_wstrb_7,io_in_wdata_bits_wstrb_6,io_in_wdata_bits_wstrb_5,io_in_wdata_bits_wstrb_4,io_in_wdata_bits_wstrb_3,io_in_wdata_bits_wstrb_2,io_in_wdata_bits_wstrb_1}; // @[Cat.scala 30:58:@149861.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? io_M_AXI_AWREADY : io_M_AXI_ARREADY; // @[MAGToAXI4Bridge.scala 36:21:@149769.4]
  assign io_in_wdata_ready = io_M_AXI_WREADY; // @[MAGToAXI4Bridge.scala 56:21:@149866.4]
  assign io_in_wresp_valid = io_M_AXI_BVALID; // @[MAGToAXI4Bridge.scala 71:21:@149919.4]
  assign io_in_wresp_bits_tag = io_M_AXI_BID; // @[MAGToAXI4Bridge.scala 74:24:@149921.4]
  assign io_M_AXI_AWID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 39:21:@149770.4]
  assign io_M_AXI_AWADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 40:21:@149771.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@149775.4]
  assign io_M_AXI_AWVALID = io_in_cmd_valid & io_in_cmd_bits_isWr; // @[MAGToAXI4Bridge.scala 49:21:@149783.4]
  assign io_M_AXI_ARID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 25:21:@149753.4]
  assign io_M_AXI_ARADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 26:21:@149754.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@149758.4]
  assign io_M_AXI_ARVALID = io_in_cmd_valid & _T_228; // @[MAGToAXI4Bridge.scala 35:21:@149767.4]
  assign io_M_AXI_WDATA = {_T_255,io_in_wdata_bits_wdata_0}; // @[MAGToAXI4Bridge.scala 52:21:@149799.4]
  assign io_M_AXI_WSTRB = {_T_318,io_in_wdata_bits_wstrb_0}; // @[MAGToAXI4Bridge.scala 53:21:@149863.4]
  assign io_M_AXI_WLAST = io_in_wdata_bits_wlast; // @[MAGToAXI4Bridge.scala 54:21:@149864.4]
  assign io_M_AXI_WVALID = io_in_wdata_valid; // @[MAGToAXI4Bridge.scala 55:21:@149865.4]
  assign io_M_AXI_RREADY = io_in_rresp_ready; // @[MAGToAXI4Bridge.scala 64:19:@149916.4]
  assign io_M_AXI_BREADY = io_in_wresp_ready; // @[MAGToAXI4Bridge.scala 67:19:@149917.4]
endmodule
module FringeZynq( // @[:@150907.2]
  input          clock, // @[:@150908.4]
  input          reset, // @[:@150909.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@150910.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@150910.4]
  input          io_S_AXI_AWVALID, // @[:@150910.4]
  output         io_S_AXI_AWREADY, // @[:@150910.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@150910.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@150910.4]
  input          io_S_AXI_ARVALID, // @[:@150910.4]
  output         io_S_AXI_ARREADY, // @[:@150910.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@150910.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@150910.4]
  input          io_S_AXI_WVALID, // @[:@150910.4]
  output         io_S_AXI_WREADY, // @[:@150910.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@150910.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@150910.4]
  output         io_S_AXI_RVALID, // @[:@150910.4]
  input          io_S_AXI_RREADY, // @[:@150910.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@150910.4]
  output         io_S_AXI_BVALID, // @[:@150910.4]
  input          io_S_AXI_BREADY, // @[:@150910.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@150910.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@150910.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@150910.4]
  output         io_M_AXI_0_AWVALID, // @[:@150910.4]
  input          io_M_AXI_0_AWREADY, // @[:@150910.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@150910.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@150910.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@150910.4]
  output         io_M_AXI_0_ARVALID, // @[:@150910.4]
  input          io_M_AXI_0_ARREADY, // @[:@150910.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@150910.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@150910.4]
  output         io_M_AXI_0_WLAST, // @[:@150910.4]
  output         io_M_AXI_0_WVALID, // @[:@150910.4]
  input          io_M_AXI_0_WREADY, // @[:@150910.4]
  output         io_M_AXI_0_RREADY, // @[:@150910.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@150910.4]
  input          io_M_AXI_0_BVALID, // @[:@150910.4]
  output         io_M_AXI_0_BREADY, // @[:@150910.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@150910.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@150910.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@150910.4]
  output         io_M_AXI_1_AWVALID, // @[:@150910.4]
  input          io_M_AXI_1_AWREADY, // @[:@150910.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@150910.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@150910.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@150910.4]
  output         io_M_AXI_1_ARVALID, // @[:@150910.4]
  input          io_M_AXI_1_ARREADY, // @[:@150910.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@150910.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@150910.4]
  output         io_M_AXI_1_WLAST, // @[:@150910.4]
  output         io_M_AXI_1_WVALID, // @[:@150910.4]
  input          io_M_AXI_1_WREADY, // @[:@150910.4]
  output         io_M_AXI_1_RREADY, // @[:@150910.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@150910.4]
  input          io_M_AXI_1_BVALID, // @[:@150910.4]
  output         io_M_AXI_1_BREADY, // @[:@150910.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@150910.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@150910.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@150910.4]
  output         io_M_AXI_2_AWVALID, // @[:@150910.4]
  input          io_M_AXI_2_AWREADY, // @[:@150910.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@150910.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@150910.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@150910.4]
  output         io_M_AXI_2_ARVALID, // @[:@150910.4]
  input          io_M_AXI_2_ARREADY, // @[:@150910.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@150910.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@150910.4]
  output         io_M_AXI_2_WLAST, // @[:@150910.4]
  output         io_M_AXI_2_WVALID, // @[:@150910.4]
  input          io_M_AXI_2_WREADY, // @[:@150910.4]
  output         io_M_AXI_2_RREADY, // @[:@150910.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@150910.4]
  input          io_M_AXI_2_BVALID, // @[:@150910.4]
  output         io_M_AXI_2_BREADY, // @[:@150910.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@150910.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@150910.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@150910.4]
  output         io_M_AXI_3_AWVALID, // @[:@150910.4]
  input          io_M_AXI_3_AWREADY, // @[:@150910.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@150910.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@150910.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@150910.4]
  output         io_M_AXI_3_ARVALID, // @[:@150910.4]
  input          io_M_AXI_3_ARREADY, // @[:@150910.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@150910.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@150910.4]
  output         io_M_AXI_3_WLAST, // @[:@150910.4]
  output         io_M_AXI_3_WVALID, // @[:@150910.4]
  input          io_M_AXI_3_WREADY, // @[:@150910.4]
  output         io_M_AXI_3_RREADY, // @[:@150910.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@150910.4]
  input          io_M_AXI_3_BVALID, // @[:@150910.4]
  output         io_M_AXI_3_BREADY, // @[:@150910.4]
  output         io_enable, // @[:@150910.4]
  input          io_done, // @[:@150910.4]
  output         io_reset, // @[:@150910.4]
  output [63:0]  io_argIns_0, // @[:@150910.4]
  output [63:0]  io_argIns_1, // @[:@150910.4]
  input          io_argOuts_0_valid, // @[:@150910.4]
  input  [63:0]  io_argOuts_0_bits, // @[:@150910.4]
  output         io_memStreams_stores_0_cmd_ready, // @[:@150910.4]
  input          io_memStreams_stores_0_cmd_valid, // @[:@150910.4]
  input  [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@150910.4]
  input  [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@150910.4]
  output         io_memStreams_stores_0_data_ready, // @[:@150910.4]
  input          io_memStreams_stores_0_data_valid, // @[:@150910.4]
  input  [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@150910.4]
  input          io_memStreams_stores_0_data_bits_wstrb, // @[:@150910.4]
  input          io_memStreams_stores_0_wresp_ready, // @[:@150910.4]
  output         io_memStreams_stores_0_wresp_valid, // @[:@150910.4]
  output         io_memStreams_stores_0_wresp_bits, // @[:@150910.4]
  input          io_heap_0_req_valid, // @[:@150910.4]
  input          io_heap_0_req_bits_allocDealloc, // @[:@150910.4]
  input  [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@150910.4]
  output         io_heap_0_resp_valid, // @[:@150910.4]
  output         io_heap_0_resp_bits_allocDealloc, // @[:@150910.4]
  output [63:0]  io_heap_0_resp_bits_sizeAddr // @[:@150910.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_raddr; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_wen; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_waddr; // @[FringeZynq.scala 69:28:@151381.4]
  wire [63:0] fringeCommon_io_wdata; // @[FringeZynq.scala 69:28:@151381.4]
  wire [63:0] fringeCommon_io_rdata; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 69:28:@151381.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 69:28:@151381.4]
  wire [63:0] fringeCommon_io_argIns_1; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 69:28:@151381.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 69:28:@151381.4]
  wire [63:0] fringeCommon_io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_cmd_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 69:28:@151381.4]
  wire [63:0] fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_0_wresp_valid; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_0_wresp_bits_tag; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_cmd_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 69:28:@151381.4]
  wire [63:0] fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_1_wresp_valid; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_1_wresp_bits_tag; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_cmd_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 69:28:@151381.4]
  wire [63:0] fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_2_wresp_valid; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_2_wresp_bits_tag; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_cmd_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 69:28:@151381.4]
  wire [63:0] fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_dram_3_wresp_valid; // @[FringeZynq.scala 69:28:@151381.4]
  wire [31:0] fringeCommon_io_dram_3_wresp_bits_tag; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_heap_0_req_valid; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 69:28:@151381.4]
  wire [63:0] fringeCommon_io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 69:28:@151381.4]
  wire  fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 69:28:@151381.4]
  wire [63:0] fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 69:28:@151381.4]
  wire  AXI4LiteToRFBridge_clock; // @[FringeZynq.scala 90:31:@152287.4]
  wire  AXI4LiteToRFBridge_reset; // @[FringeZynq.scala 90:31:@152287.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_AWADDR; // @[FringeZynq.scala 90:31:@152287.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_AWPROT; // @[FringeZynq.scala 90:31:@152287.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWVALID; // @[FringeZynq.scala 90:31:@152287.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 90:31:@152287.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_ARADDR; // @[FringeZynq.scala 90:31:@152287.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_ARPROT; // @[FringeZynq.scala 90:31:@152287.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARVALID; // @[FringeZynq.scala 90:31:@152287.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 90:31:@152287.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_WDATA; // @[FringeZynq.scala 90:31:@152287.4]
  wire [3:0] AXI4LiteToRFBridge_io_S_AXI_WSTRB; // @[FringeZynq.scala 90:31:@152287.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WVALID; // @[FringeZynq.scala 90:31:@152287.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 90:31:@152287.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 90:31:@152287.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 90:31:@152287.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 90:31:@152287.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RREADY; // @[FringeZynq.scala 90:31:@152287.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 90:31:@152287.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 90:31:@152287.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BREADY; // @[FringeZynq.scala 90:31:@152287.4]
  wire [31:0] AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 90:31:@152287.4]
  wire  AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 90:31:@152287.4]
  wire [31:0] AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 90:31:@152287.4]
  wire [31:0] AXI4LiteToRFBridge_io_wdata; // @[FringeZynq.scala 90:31:@152287.4]
  wire [31:0] AXI4LiteToRFBridge_io_rdata; // @[FringeZynq.scala 90:31:@152287.4]
  wire  MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@152437.4]
  wire [63:0] MAGToAXI4Bridge_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@152437.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@152437.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@152437.4]
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@152437.4]
  wire [63:0] MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@152437.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@152437.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@152593.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@152593.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@152593.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@152593.4]
  wire [511:0] MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@152593.4]
  wire [63:0] MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@152593.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@152593.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@152749.4]
  wire [63:0] MAGToAXI4Bridge_2_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@152749.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@152749.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@152749.4]
  wire [511:0] MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@152749.4]
  wire [63:0] MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@152749.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@152749.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@152905.4]
  wire [63:0] MAGToAXI4Bridge_3_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@152905.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@152905.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@152905.4]
  wire [511:0] MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@152905.4]
  wire [63:0] MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@152905.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@152905.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@152905.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 69:28:@151381.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argIns_1(fringeCommon_io_argIns_1),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(fringeCommon_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(fringeCommon_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(fringeCommon_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(fringeCommon_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(fringeCommon_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(fringeCommon_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(fringeCommon_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(fringeCommon_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(fringeCommon_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(fringeCommon_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(fringeCommon_io_memStreams_stores_0_wresp_bits),
    .io_dram_0_cmd_ready(fringeCommon_io_dram_0_cmd_ready),
    .io_dram_0_cmd_valid(fringeCommon_io_dram_0_cmd_valid),
    .io_dram_0_cmd_bits_addr(fringeCommon_io_dram_0_cmd_bits_addr),
    .io_dram_0_cmd_bits_size(fringeCommon_io_dram_0_cmd_bits_size),
    .io_dram_0_cmd_bits_isWr(fringeCommon_io_dram_0_cmd_bits_isWr),
    .io_dram_0_cmd_bits_tag(fringeCommon_io_dram_0_cmd_bits_tag),
    .io_dram_0_wdata_ready(fringeCommon_io_dram_0_wdata_ready),
    .io_dram_0_wdata_valid(fringeCommon_io_dram_0_wdata_valid),
    .io_dram_0_wdata_bits_wdata_0(fringeCommon_io_dram_0_wdata_bits_wdata_0),
    .io_dram_0_wdata_bits_wdata_1(fringeCommon_io_dram_0_wdata_bits_wdata_1),
    .io_dram_0_wdata_bits_wdata_2(fringeCommon_io_dram_0_wdata_bits_wdata_2),
    .io_dram_0_wdata_bits_wdata_3(fringeCommon_io_dram_0_wdata_bits_wdata_3),
    .io_dram_0_wdata_bits_wdata_4(fringeCommon_io_dram_0_wdata_bits_wdata_4),
    .io_dram_0_wdata_bits_wdata_5(fringeCommon_io_dram_0_wdata_bits_wdata_5),
    .io_dram_0_wdata_bits_wdata_6(fringeCommon_io_dram_0_wdata_bits_wdata_6),
    .io_dram_0_wdata_bits_wdata_7(fringeCommon_io_dram_0_wdata_bits_wdata_7),
    .io_dram_0_wdata_bits_wdata_8(fringeCommon_io_dram_0_wdata_bits_wdata_8),
    .io_dram_0_wdata_bits_wdata_9(fringeCommon_io_dram_0_wdata_bits_wdata_9),
    .io_dram_0_wdata_bits_wdata_10(fringeCommon_io_dram_0_wdata_bits_wdata_10),
    .io_dram_0_wdata_bits_wdata_11(fringeCommon_io_dram_0_wdata_bits_wdata_11),
    .io_dram_0_wdata_bits_wdata_12(fringeCommon_io_dram_0_wdata_bits_wdata_12),
    .io_dram_0_wdata_bits_wdata_13(fringeCommon_io_dram_0_wdata_bits_wdata_13),
    .io_dram_0_wdata_bits_wdata_14(fringeCommon_io_dram_0_wdata_bits_wdata_14),
    .io_dram_0_wdata_bits_wdata_15(fringeCommon_io_dram_0_wdata_bits_wdata_15),
    .io_dram_0_wdata_bits_wstrb_0(fringeCommon_io_dram_0_wdata_bits_wstrb_0),
    .io_dram_0_wdata_bits_wstrb_1(fringeCommon_io_dram_0_wdata_bits_wstrb_1),
    .io_dram_0_wdata_bits_wstrb_2(fringeCommon_io_dram_0_wdata_bits_wstrb_2),
    .io_dram_0_wdata_bits_wstrb_3(fringeCommon_io_dram_0_wdata_bits_wstrb_3),
    .io_dram_0_wdata_bits_wstrb_4(fringeCommon_io_dram_0_wdata_bits_wstrb_4),
    .io_dram_0_wdata_bits_wstrb_5(fringeCommon_io_dram_0_wdata_bits_wstrb_5),
    .io_dram_0_wdata_bits_wstrb_6(fringeCommon_io_dram_0_wdata_bits_wstrb_6),
    .io_dram_0_wdata_bits_wstrb_7(fringeCommon_io_dram_0_wdata_bits_wstrb_7),
    .io_dram_0_wdata_bits_wstrb_8(fringeCommon_io_dram_0_wdata_bits_wstrb_8),
    .io_dram_0_wdata_bits_wstrb_9(fringeCommon_io_dram_0_wdata_bits_wstrb_9),
    .io_dram_0_wdata_bits_wstrb_10(fringeCommon_io_dram_0_wdata_bits_wstrb_10),
    .io_dram_0_wdata_bits_wstrb_11(fringeCommon_io_dram_0_wdata_bits_wstrb_11),
    .io_dram_0_wdata_bits_wstrb_12(fringeCommon_io_dram_0_wdata_bits_wstrb_12),
    .io_dram_0_wdata_bits_wstrb_13(fringeCommon_io_dram_0_wdata_bits_wstrb_13),
    .io_dram_0_wdata_bits_wstrb_14(fringeCommon_io_dram_0_wdata_bits_wstrb_14),
    .io_dram_0_wdata_bits_wstrb_15(fringeCommon_io_dram_0_wdata_bits_wstrb_15),
    .io_dram_0_wdata_bits_wstrb_16(fringeCommon_io_dram_0_wdata_bits_wstrb_16),
    .io_dram_0_wdata_bits_wstrb_17(fringeCommon_io_dram_0_wdata_bits_wstrb_17),
    .io_dram_0_wdata_bits_wstrb_18(fringeCommon_io_dram_0_wdata_bits_wstrb_18),
    .io_dram_0_wdata_bits_wstrb_19(fringeCommon_io_dram_0_wdata_bits_wstrb_19),
    .io_dram_0_wdata_bits_wstrb_20(fringeCommon_io_dram_0_wdata_bits_wstrb_20),
    .io_dram_0_wdata_bits_wstrb_21(fringeCommon_io_dram_0_wdata_bits_wstrb_21),
    .io_dram_0_wdata_bits_wstrb_22(fringeCommon_io_dram_0_wdata_bits_wstrb_22),
    .io_dram_0_wdata_bits_wstrb_23(fringeCommon_io_dram_0_wdata_bits_wstrb_23),
    .io_dram_0_wdata_bits_wstrb_24(fringeCommon_io_dram_0_wdata_bits_wstrb_24),
    .io_dram_0_wdata_bits_wstrb_25(fringeCommon_io_dram_0_wdata_bits_wstrb_25),
    .io_dram_0_wdata_bits_wstrb_26(fringeCommon_io_dram_0_wdata_bits_wstrb_26),
    .io_dram_0_wdata_bits_wstrb_27(fringeCommon_io_dram_0_wdata_bits_wstrb_27),
    .io_dram_0_wdata_bits_wstrb_28(fringeCommon_io_dram_0_wdata_bits_wstrb_28),
    .io_dram_0_wdata_bits_wstrb_29(fringeCommon_io_dram_0_wdata_bits_wstrb_29),
    .io_dram_0_wdata_bits_wstrb_30(fringeCommon_io_dram_0_wdata_bits_wstrb_30),
    .io_dram_0_wdata_bits_wstrb_31(fringeCommon_io_dram_0_wdata_bits_wstrb_31),
    .io_dram_0_wdata_bits_wstrb_32(fringeCommon_io_dram_0_wdata_bits_wstrb_32),
    .io_dram_0_wdata_bits_wstrb_33(fringeCommon_io_dram_0_wdata_bits_wstrb_33),
    .io_dram_0_wdata_bits_wstrb_34(fringeCommon_io_dram_0_wdata_bits_wstrb_34),
    .io_dram_0_wdata_bits_wstrb_35(fringeCommon_io_dram_0_wdata_bits_wstrb_35),
    .io_dram_0_wdata_bits_wstrb_36(fringeCommon_io_dram_0_wdata_bits_wstrb_36),
    .io_dram_0_wdata_bits_wstrb_37(fringeCommon_io_dram_0_wdata_bits_wstrb_37),
    .io_dram_0_wdata_bits_wstrb_38(fringeCommon_io_dram_0_wdata_bits_wstrb_38),
    .io_dram_0_wdata_bits_wstrb_39(fringeCommon_io_dram_0_wdata_bits_wstrb_39),
    .io_dram_0_wdata_bits_wstrb_40(fringeCommon_io_dram_0_wdata_bits_wstrb_40),
    .io_dram_0_wdata_bits_wstrb_41(fringeCommon_io_dram_0_wdata_bits_wstrb_41),
    .io_dram_0_wdata_bits_wstrb_42(fringeCommon_io_dram_0_wdata_bits_wstrb_42),
    .io_dram_0_wdata_bits_wstrb_43(fringeCommon_io_dram_0_wdata_bits_wstrb_43),
    .io_dram_0_wdata_bits_wstrb_44(fringeCommon_io_dram_0_wdata_bits_wstrb_44),
    .io_dram_0_wdata_bits_wstrb_45(fringeCommon_io_dram_0_wdata_bits_wstrb_45),
    .io_dram_0_wdata_bits_wstrb_46(fringeCommon_io_dram_0_wdata_bits_wstrb_46),
    .io_dram_0_wdata_bits_wstrb_47(fringeCommon_io_dram_0_wdata_bits_wstrb_47),
    .io_dram_0_wdata_bits_wstrb_48(fringeCommon_io_dram_0_wdata_bits_wstrb_48),
    .io_dram_0_wdata_bits_wstrb_49(fringeCommon_io_dram_0_wdata_bits_wstrb_49),
    .io_dram_0_wdata_bits_wstrb_50(fringeCommon_io_dram_0_wdata_bits_wstrb_50),
    .io_dram_0_wdata_bits_wstrb_51(fringeCommon_io_dram_0_wdata_bits_wstrb_51),
    .io_dram_0_wdata_bits_wstrb_52(fringeCommon_io_dram_0_wdata_bits_wstrb_52),
    .io_dram_0_wdata_bits_wstrb_53(fringeCommon_io_dram_0_wdata_bits_wstrb_53),
    .io_dram_0_wdata_bits_wstrb_54(fringeCommon_io_dram_0_wdata_bits_wstrb_54),
    .io_dram_0_wdata_bits_wstrb_55(fringeCommon_io_dram_0_wdata_bits_wstrb_55),
    .io_dram_0_wdata_bits_wstrb_56(fringeCommon_io_dram_0_wdata_bits_wstrb_56),
    .io_dram_0_wdata_bits_wstrb_57(fringeCommon_io_dram_0_wdata_bits_wstrb_57),
    .io_dram_0_wdata_bits_wstrb_58(fringeCommon_io_dram_0_wdata_bits_wstrb_58),
    .io_dram_0_wdata_bits_wstrb_59(fringeCommon_io_dram_0_wdata_bits_wstrb_59),
    .io_dram_0_wdata_bits_wstrb_60(fringeCommon_io_dram_0_wdata_bits_wstrb_60),
    .io_dram_0_wdata_bits_wstrb_61(fringeCommon_io_dram_0_wdata_bits_wstrb_61),
    .io_dram_0_wdata_bits_wstrb_62(fringeCommon_io_dram_0_wdata_bits_wstrb_62),
    .io_dram_0_wdata_bits_wstrb_63(fringeCommon_io_dram_0_wdata_bits_wstrb_63),
    .io_dram_0_wdata_bits_wlast(fringeCommon_io_dram_0_wdata_bits_wlast),
    .io_dram_0_rresp_ready(fringeCommon_io_dram_0_rresp_ready),
    .io_dram_0_wresp_ready(fringeCommon_io_dram_0_wresp_ready),
    .io_dram_0_wresp_valid(fringeCommon_io_dram_0_wresp_valid),
    .io_dram_0_wresp_bits_tag(fringeCommon_io_dram_0_wresp_bits_tag),
    .io_dram_1_cmd_ready(fringeCommon_io_dram_1_cmd_ready),
    .io_dram_1_cmd_valid(fringeCommon_io_dram_1_cmd_valid),
    .io_dram_1_cmd_bits_addr(fringeCommon_io_dram_1_cmd_bits_addr),
    .io_dram_1_cmd_bits_size(fringeCommon_io_dram_1_cmd_bits_size),
    .io_dram_1_cmd_bits_isWr(fringeCommon_io_dram_1_cmd_bits_isWr),
    .io_dram_1_cmd_bits_tag(fringeCommon_io_dram_1_cmd_bits_tag),
    .io_dram_1_wdata_ready(fringeCommon_io_dram_1_wdata_ready),
    .io_dram_1_wdata_valid(fringeCommon_io_dram_1_wdata_valid),
    .io_dram_1_wdata_bits_wdata_0(fringeCommon_io_dram_1_wdata_bits_wdata_0),
    .io_dram_1_wdata_bits_wdata_1(fringeCommon_io_dram_1_wdata_bits_wdata_1),
    .io_dram_1_wdata_bits_wdata_2(fringeCommon_io_dram_1_wdata_bits_wdata_2),
    .io_dram_1_wdata_bits_wdata_3(fringeCommon_io_dram_1_wdata_bits_wdata_3),
    .io_dram_1_wdata_bits_wdata_4(fringeCommon_io_dram_1_wdata_bits_wdata_4),
    .io_dram_1_wdata_bits_wdata_5(fringeCommon_io_dram_1_wdata_bits_wdata_5),
    .io_dram_1_wdata_bits_wdata_6(fringeCommon_io_dram_1_wdata_bits_wdata_6),
    .io_dram_1_wdata_bits_wdata_7(fringeCommon_io_dram_1_wdata_bits_wdata_7),
    .io_dram_1_wdata_bits_wdata_8(fringeCommon_io_dram_1_wdata_bits_wdata_8),
    .io_dram_1_wdata_bits_wdata_9(fringeCommon_io_dram_1_wdata_bits_wdata_9),
    .io_dram_1_wdata_bits_wdata_10(fringeCommon_io_dram_1_wdata_bits_wdata_10),
    .io_dram_1_wdata_bits_wdata_11(fringeCommon_io_dram_1_wdata_bits_wdata_11),
    .io_dram_1_wdata_bits_wdata_12(fringeCommon_io_dram_1_wdata_bits_wdata_12),
    .io_dram_1_wdata_bits_wdata_13(fringeCommon_io_dram_1_wdata_bits_wdata_13),
    .io_dram_1_wdata_bits_wdata_14(fringeCommon_io_dram_1_wdata_bits_wdata_14),
    .io_dram_1_wdata_bits_wdata_15(fringeCommon_io_dram_1_wdata_bits_wdata_15),
    .io_dram_1_wdata_bits_wstrb_0(fringeCommon_io_dram_1_wdata_bits_wstrb_0),
    .io_dram_1_wdata_bits_wstrb_1(fringeCommon_io_dram_1_wdata_bits_wstrb_1),
    .io_dram_1_wdata_bits_wstrb_2(fringeCommon_io_dram_1_wdata_bits_wstrb_2),
    .io_dram_1_wdata_bits_wstrb_3(fringeCommon_io_dram_1_wdata_bits_wstrb_3),
    .io_dram_1_wdata_bits_wstrb_4(fringeCommon_io_dram_1_wdata_bits_wstrb_4),
    .io_dram_1_wdata_bits_wstrb_5(fringeCommon_io_dram_1_wdata_bits_wstrb_5),
    .io_dram_1_wdata_bits_wstrb_6(fringeCommon_io_dram_1_wdata_bits_wstrb_6),
    .io_dram_1_wdata_bits_wstrb_7(fringeCommon_io_dram_1_wdata_bits_wstrb_7),
    .io_dram_1_wdata_bits_wstrb_8(fringeCommon_io_dram_1_wdata_bits_wstrb_8),
    .io_dram_1_wdata_bits_wstrb_9(fringeCommon_io_dram_1_wdata_bits_wstrb_9),
    .io_dram_1_wdata_bits_wstrb_10(fringeCommon_io_dram_1_wdata_bits_wstrb_10),
    .io_dram_1_wdata_bits_wstrb_11(fringeCommon_io_dram_1_wdata_bits_wstrb_11),
    .io_dram_1_wdata_bits_wstrb_12(fringeCommon_io_dram_1_wdata_bits_wstrb_12),
    .io_dram_1_wdata_bits_wstrb_13(fringeCommon_io_dram_1_wdata_bits_wstrb_13),
    .io_dram_1_wdata_bits_wstrb_14(fringeCommon_io_dram_1_wdata_bits_wstrb_14),
    .io_dram_1_wdata_bits_wstrb_15(fringeCommon_io_dram_1_wdata_bits_wstrb_15),
    .io_dram_1_wdata_bits_wstrb_16(fringeCommon_io_dram_1_wdata_bits_wstrb_16),
    .io_dram_1_wdata_bits_wstrb_17(fringeCommon_io_dram_1_wdata_bits_wstrb_17),
    .io_dram_1_wdata_bits_wstrb_18(fringeCommon_io_dram_1_wdata_bits_wstrb_18),
    .io_dram_1_wdata_bits_wstrb_19(fringeCommon_io_dram_1_wdata_bits_wstrb_19),
    .io_dram_1_wdata_bits_wstrb_20(fringeCommon_io_dram_1_wdata_bits_wstrb_20),
    .io_dram_1_wdata_bits_wstrb_21(fringeCommon_io_dram_1_wdata_bits_wstrb_21),
    .io_dram_1_wdata_bits_wstrb_22(fringeCommon_io_dram_1_wdata_bits_wstrb_22),
    .io_dram_1_wdata_bits_wstrb_23(fringeCommon_io_dram_1_wdata_bits_wstrb_23),
    .io_dram_1_wdata_bits_wstrb_24(fringeCommon_io_dram_1_wdata_bits_wstrb_24),
    .io_dram_1_wdata_bits_wstrb_25(fringeCommon_io_dram_1_wdata_bits_wstrb_25),
    .io_dram_1_wdata_bits_wstrb_26(fringeCommon_io_dram_1_wdata_bits_wstrb_26),
    .io_dram_1_wdata_bits_wstrb_27(fringeCommon_io_dram_1_wdata_bits_wstrb_27),
    .io_dram_1_wdata_bits_wstrb_28(fringeCommon_io_dram_1_wdata_bits_wstrb_28),
    .io_dram_1_wdata_bits_wstrb_29(fringeCommon_io_dram_1_wdata_bits_wstrb_29),
    .io_dram_1_wdata_bits_wstrb_30(fringeCommon_io_dram_1_wdata_bits_wstrb_30),
    .io_dram_1_wdata_bits_wstrb_31(fringeCommon_io_dram_1_wdata_bits_wstrb_31),
    .io_dram_1_wdata_bits_wstrb_32(fringeCommon_io_dram_1_wdata_bits_wstrb_32),
    .io_dram_1_wdata_bits_wstrb_33(fringeCommon_io_dram_1_wdata_bits_wstrb_33),
    .io_dram_1_wdata_bits_wstrb_34(fringeCommon_io_dram_1_wdata_bits_wstrb_34),
    .io_dram_1_wdata_bits_wstrb_35(fringeCommon_io_dram_1_wdata_bits_wstrb_35),
    .io_dram_1_wdata_bits_wstrb_36(fringeCommon_io_dram_1_wdata_bits_wstrb_36),
    .io_dram_1_wdata_bits_wstrb_37(fringeCommon_io_dram_1_wdata_bits_wstrb_37),
    .io_dram_1_wdata_bits_wstrb_38(fringeCommon_io_dram_1_wdata_bits_wstrb_38),
    .io_dram_1_wdata_bits_wstrb_39(fringeCommon_io_dram_1_wdata_bits_wstrb_39),
    .io_dram_1_wdata_bits_wstrb_40(fringeCommon_io_dram_1_wdata_bits_wstrb_40),
    .io_dram_1_wdata_bits_wstrb_41(fringeCommon_io_dram_1_wdata_bits_wstrb_41),
    .io_dram_1_wdata_bits_wstrb_42(fringeCommon_io_dram_1_wdata_bits_wstrb_42),
    .io_dram_1_wdata_bits_wstrb_43(fringeCommon_io_dram_1_wdata_bits_wstrb_43),
    .io_dram_1_wdata_bits_wstrb_44(fringeCommon_io_dram_1_wdata_bits_wstrb_44),
    .io_dram_1_wdata_bits_wstrb_45(fringeCommon_io_dram_1_wdata_bits_wstrb_45),
    .io_dram_1_wdata_bits_wstrb_46(fringeCommon_io_dram_1_wdata_bits_wstrb_46),
    .io_dram_1_wdata_bits_wstrb_47(fringeCommon_io_dram_1_wdata_bits_wstrb_47),
    .io_dram_1_wdata_bits_wstrb_48(fringeCommon_io_dram_1_wdata_bits_wstrb_48),
    .io_dram_1_wdata_bits_wstrb_49(fringeCommon_io_dram_1_wdata_bits_wstrb_49),
    .io_dram_1_wdata_bits_wstrb_50(fringeCommon_io_dram_1_wdata_bits_wstrb_50),
    .io_dram_1_wdata_bits_wstrb_51(fringeCommon_io_dram_1_wdata_bits_wstrb_51),
    .io_dram_1_wdata_bits_wstrb_52(fringeCommon_io_dram_1_wdata_bits_wstrb_52),
    .io_dram_1_wdata_bits_wstrb_53(fringeCommon_io_dram_1_wdata_bits_wstrb_53),
    .io_dram_1_wdata_bits_wstrb_54(fringeCommon_io_dram_1_wdata_bits_wstrb_54),
    .io_dram_1_wdata_bits_wstrb_55(fringeCommon_io_dram_1_wdata_bits_wstrb_55),
    .io_dram_1_wdata_bits_wstrb_56(fringeCommon_io_dram_1_wdata_bits_wstrb_56),
    .io_dram_1_wdata_bits_wstrb_57(fringeCommon_io_dram_1_wdata_bits_wstrb_57),
    .io_dram_1_wdata_bits_wstrb_58(fringeCommon_io_dram_1_wdata_bits_wstrb_58),
    .io_dram_1_wdata_bits_wstrb_59(fringeCommon_io_dram_1_wdata_bits_wstrb_59),
    .io_dram_1_wdata_bits_wstrb_60(fringeCommon_io_dram_1_wdata_bits_wstrb_60),
    .io_dram_1_wdata_bits_wstrb_61(fringeCommon_io_dram_1_wdata_bits_wstrb_61),
    .io_dram_1_wdata_bits_wstrb_62(fringeCommon_io_dram_1_wdata_bits_wstrb_62),
    .io_dram_1_wdata_bits_wstrb_63(fringeCommon_io_dram_1_wdata_bits_wstrb_63),
    .io_dram_1_wdata_bits_wlast(fringeCommon_io_dram_1_wdata_bits_wlast),
    .io_dram_1_rresp_ready(fringeCommon_io_dram_1_rresp_ready),
    .io_dram_1_wresp_ready(fringeCommon_io_dram_1_wresp_ready),
    .io_dram_1_wresp_valid(fringeCommon_io_dram_1_wresp_valid),
    .io_dram_1_wresp_bits_tag(fringeCommon_io_dram_1_wresp_bits_tag),
    .io_dram_2_cmd_ready(fringeCommon_io_dram_2_cmd_ready),
    .io_dram_2_cmd_valid(fringeCommon_io_dram_2_cmd_valid),
    .io_dram_2_cmd_bits_addr(fringeCommon_io_dram_2_cmd_bits_addr),
    .io_dram_2_cmd_bits_size(fringeCommon_io_dram_2_cmd_bits_size),
    .io_dram_2_cmd_bits_isWr(fringeCommon_io_dram_2_cmd_bits_isWr),
    .io_dram_2_cmd_bits_tag(fringeCommon_io_dram_2_cmd_bits_tag),
    .io_dram_2_wdata_ready(fringeCommon_io_dram_2_wdata_ready),
    .io_dram_2_wdata_valid(fringeCommon_io_dram_2_wdata_valid),
    .io_dram_2_wdata_bits_wdata_0(fringeCommon_io_dram_2_wdata_bits_wdata_0),
    .io_dram_2_wdata_bits_wdata_1(fringeCommon_io_dram_2_wdata_bits_wdata_1),
    .io_dram_2_wdata_bits_wdata_2(fringeCommon_io_dram_2_wdata_bits_wdata_2),
    .io_dram_2_wdata_bits_wdata_3(fringeCommon_io_dram_2_wdata_bits_wdata_3),
    .io_dram_2_wdata_bits_wdata_4(fringeCommon_io_dram_2_wdata_bits_wdata_4),
    .io_dram_2_wdata_bits_wdata_5(fringeCommon_io_dram_2_wdata_bits_wdata_5),
    .io_dram_2_wdata_bits_wdata_6(fringeCommon_io_dram_2_wdata_bits_wdata_6),
    .io_dram_2_wdata_bits_wdata_7(fringeCommon_io_dram_2_wdata_bits_wdata_7),
    .io_dram_2_wdata_bits_wdata_8(fringeCommon_io_dram_2_wdata_bits_wdata_8),
    .io_dram_2_wdata_bits_wdata_9(fringeCommon_io_dram_2_wdata_bits_wdata_9),
    .io_dram_2_wdata_bits_wdata_10(fringeCommon_io_dram_2_wdata_bits_wdata_10),
    .io_dram_2_wdata_bits_wdata_11(fringeCommon_io_dram_2_wdata_bits_wdata_11),
    .io_dram_2_wdata_bits_wdata_12(fringeCommon_io_dram_2_wdata_bits_wdata_12),
    .io_dram_2_wdata_bits_wdata_13(fringeCommon_io_dram_2_wdata_bits_wdata_13),
    .io_dram_2_wdata_bits_wdata_14(fringeCommon_io_dram_2_wdata_bits_wdata_14),
    .io_dram_2_wdata_bits_wdata_15(fringeCommon_io_dram_2_wdata_bits_wdata_15),
    .io_dram_2_wdata_bits_wstrb_0(fringeCommon_io_dram_2_wdata_bits_wstrb_0),
    .io_dram_2_wdata_bits_wstrb_1(fringeCommon_io_dram_2_wdata_bits_wstrb_1),
    .io_dram_2_wdata_bits_wstrb_2(fringeCommon_io_dram_2_wdata_bits_wstrb_2),
    .io_dram_2_wdata_bits_wstrb_3(fringeCommon_io_dram_2_wdata_bits_wstrb_3),
    .io_dram_2_wdata_bits_wstrb_4(fringeCommon_io_dram_2_wdata_bits_wstrb_4),
    .io_dram_2_wdata_bits_wstrb_5(fringeCommon_io_dram_2_wdata_bits_wstrb_5),
    .io_dram_2_wdata_bits_wstrb_6(fringeCommon_io_dram_2_wdata_bits_wstrb_6),
    .io_dram_2_wdata_bits_wstrb_7(fringeCommon_io_dram_2_wdata_bits_wstrb_7),
    .io_dram_2_wdata_bits_wstrb_8(fringeCommon_io_dram_2_wdata_bits_wstrb_8),
    .io_dram_2_wdata_bits_wstrb_9(fringeCommon_io_dram_2_wdata_bits_wstrb_9),
    .io_dram_2_wdata_bits_wstrb_10(fringeCommon_io_dram_2_wdata_bits_wstrb_10),
    .io_dram_2_wdata_bits_wstrb_11(fringeCommon_io_dram_2_wdata_bits_wstrb_11),
    .io_dram_2_wdata_bits_wstrb_12(fringeCommon_io_dram_2_wdata_bits_wstrb_12),
    .io_dram_2_wdata_bits_wstrb_13(fringeCommon_io_dram_2_wdata_bits_wstrb_13),
    .io_dram_2_wdata_bits_wstrb_14(fringeCommon_io_dram_2_wdata_bits_wstrb_14),
    .io_dram_2_wdata_bits_wstrb_15(fringeCommon_io_dram_2_wdata_bits_wstrb_15),
    .io_dram_2_wdata_bits_wstrb_16(fringeCommon_io_dram_2_wdata_bits_wstrb_16),
    .io_dram_2_wdata_bits_wstrb_17(fringeCommon_io_dram_2_wdata_bits_wstrb_17),
    .io_dram_2_wdata_bits_wstrb_18(fringeCommon_io_dram_2_wdata_bits_wstrb_18),
    .io_dram_2_wdata_bits_wstrb_19(fringeCommon_io_dram_2_wdata_bits_wstrb_19),
    .io_dram_2_wdata_bits_wstrb_20(fringeCommon_io_dram_2_wdata_bits_wstrb_20),
    .io_dram_2_wdata_bits_wstrb_21(fringeCommon_io_dram_2_wdata_bits_wstrb_21),
    .io_dram_2_wdata_bits_wstrb_22(fringeCommon_io_dram_2_wdata_bits_wstrb_22),
    .io_dram_2_wdata_bits_wstrb_23(fringeCommon_io_dram_2_wdata_bits_wstrb_23),
    .io_dram_2_wdata_bits_wstrb_24(fringeCommon_io_dram_2_wdata_bits_wstrb_24),
    .io_dram_2_wdata_bits_wstrb_25(fringeCommon_io_dram_2_wdata_bits_wstrb_25),
    .io_dram_2_wdata_bits_wstrb_26(fringeCommon_io_dram_2_wdata_bits_wstrb_26),
    .io_dram_2_wdata_bits_wstrb_27(fringeCommon_io_dram_2_wdata_bits_wstrb_27),
    .io_dram_2_wdata_bits_wstrb_28(fringeCommon_io_dram_2_wdata_bits_wstrb_28),
    .io_dram_2_wdata_bits_wstrb_29(fringeCommon_io_dram_2_wdata_bits_wstrb_29),
    .io_dram_2_wdata_bits_wstrb_30(fringeCommon_io_dram_2_wdata_bits_wstrb_30),
    .io_dram_2_wdata_bits_wstrb_31(fringeCommon_io_dram_2_wdata_bits_wstrb_31),
    .io_dram_2_wdata_bits_wstrb_32(fringeCommon_io_dram_2_wdata_bits_wstrb_32),
    .io_dram_2_wdata_bits_wstrb_33(fringeCommon_io_dram_2_wdata_bits_wstrb_33),
    .io_dram_2_wdata_bits_wstrb_34(fringeCommon_io_dram_2_wdata_bits_wstrb_34),
    .io_dram_2_wdata_bits_wstrb_35(fringeCommon_io_dram_2_wdata_bits_wstrb_35),
    .io_dram_2_wdata_bits_wstrb_36(fringeCommon_io_dram_2_wdata_bits_wstrb_36),
    .io_dram_2_wdata_bits_wstrb_37(fringeCommon_io_dram_2_wdata_bits_wstrb_37),
    .io_dram_2_wdata_bits_wstrb_38(fringeCommon_io_dram_2_wdata_bits_wstrb_38),
    .io_dram_2_wdata_bits_wstrb_39(fringeCommon_io_dram_2_wdata_bits_wstrb_39),
    .io_dram_2_wdata_bits_wstrb_40(fringeCommon_io_dram_2_wdata_bits_wstrb_40),
    .io_dram_2_wdata_bits_wstrb_41(fringeCommon_io_dram_2_wdata_bits_wstrb_41),
    .io_dram_2_wdata_bits_wstrb_42(fringeCommon_io_dram_2_wdata_bits_wstrb_42),
    .io_dram_2_wdata_bits_wstrb_43(fringeCommon_io_dram_2_wdata_bits_wstrb_43),
    .io_dram_2_wdata_bits_wstrb_44(fringeCommon_io_dram_2_wdata_bits_wstrb_44),
    .io_dram_2_wdata_bits_wstrb_45(fringeCommon_io_dram_2_wdata_bits_wstrb_45),
    .io_dram_2_wdata_bits_wstrb_46(fringeCommon_io_dram_2_wdata_bits_wstrb_46),
    .io_dram_2_wdata_bits_wstrb_47(fringeCommon_io_dram_2_wdata_bits_wstrb_47),
    .io_dram_2_wdata_bits_wstrb_48(fringeCommon_io_dram_2_wdata_bits_wstrb_48),
    .io_dram_2_wdata_bits_wstrb_49(fringeCommon_io_dram_2_wdata_bits_wstrb_49),
    .io_dram_2_wdata_bits_wstrb_50(fringeCommon_io_dram_2_wdata_bits_wstrb_50),
    .io_dram_2_wdata_bits_wstrb_51(fringeCommon_io_dram_2_wdata_bits_wstrb_51),
    .io_dram_2_wdata_bits_wstrb_52(fringeCommon_io_dram_2_wdata_bits_wstrb_52),
    .io_dram_2_wdata_bits_wstrb_53(fringeCommon_io_dram_2_wdata_bits_wstrb_53),
    .io_dram_2_wdata_bits_wstrb_54(fringeCommon_io_dram_2_wdata_bits_wstrb_54),
    .io_dram_2_wdata_bits_wstrb_55(fringeCommon_io_dram_2_wdata_bits_wstrb_55),
    .io_dram_2_wdata_bits_wstrb_56(fringeCommon_io_dram_2_wdata_bits_wstrb_56),
    .io_dram_2_wdata_bits_wstrb_57(fringeCommon_io_dram_2_wdata_bits_wstrb_57),
    .io_dram_2_wdata_bits_wstrb_58(fringeCommon_io_dram_2_wdata_bits_wstrb_58),
    .io_dram_2_wdata_bits_wstrb_59(fringeCommon_io_dram_2_wdata_bits_wstrb_59),
    .io_dram_2_wdata_bits_wstrb_60(fringeCommon_io_dram_2_wdata_bits_wstrb_60),
    .io_dram_2_wdata_bits_wstrb_61(fringeCommon_io_dram_2_wdata_bits_wstrb_61),
    .io_dram_2_wdata_bits_wstrb_62(fringeCommon_io_dram_2_wdata_bits_wstrb_62),
    .io_dram_2_wdata_bits_wstrb_63(fringeCommon_io_dram_2_wdata_bits_wstrb_63),
    .io_dram_2_wdata_bits_wlast(fringeCommon_io_dram_2_wdata_bits_wlast),
    .io_dram_2_rresp_ready(fringeCommon_io_dram_2_rresp_ready),
    .io_dram_2_wresp_ready(fringeCommon_io_dram_2_wresp_ready),
    .io_dram_2_wresp_valid(fringeCommon_io_dram_2_wresp_valid),
    .io_dram_2_wresp_bits_tag(fringeCommon_io_dram_2_wresp_bits_tag),
    .io_dram_3_cmd_ready(fringeCommon_io_dram_3_cmd_ready),
    .io_dram_3_cmd_valid(fringeCommon_io_dram_3_cmd_valid),
    .io_dram_3_cmd_bits_addr(fringeCommon_io_dram_3_cmd_bits_addr),
    .io_dram_3_cmd_bits_size(fringeCommon_io_dram_3_cmd_bits_size),
    .io_dram_3_cmd_bits_isWr(fringeCommon_io_dram_3_cmd_bits_isWr),
    .io_dram_3_cmd_bits_tag(fringeCommon_io_dram_3_cmd_bits_tag),
    .io_dram_3_wdata_ready(fringeCommon_io_dram_3_wdata_ready),
    .io_dram_3_wdata_valid(fringeCommon_io_dram_3_wdata_valid),
    .io_dram_3_wdata_bits_wdata_0(fringeCommon_io_dram_3_wdata_bits_wdata_0),
    .io_dram_3_wdata_bits_wdata_1(fringeCommon_io_dram_3_wdata_bits_wdata_1),
    .io_dram_3_wdata_bits_wdata_2(fringeCommon_io_dram_3_wdata_bits_wdata_2),
    .io_dram_3_wdata_bits_wdata_3(fringeCommon_io_dram_3_wdata_bits_wdata_3),
    .io_dram_3_wdata_bits_wdata_4(fringeCommon_io_dram_3_wdata_bits_wdata_4),
    .io_dram_3_wdata_bits_wdata_5(fringeCommon_io_dram_3_wdata_bits_wdata_5),
    .io_dram_3_wdata_bits_wdata_6(fringeCommon_io_dram_3_wdata_bits_wdata_6),
    .io_dram_3_wdata_bits_wdata_7(fringeCommon_io_dram_3_wdata_bits_wdata_7),
    .io_dram_3_wdata_bits_wdata_8(fringeCommon_io_dram_3_wdata_bits_wdata_8),
    .io_dram_3_wdata_bits_wdata_9(fringeCommon_io_dram_3_wdata_bits_wdata_9),
    .io_dram_3_wdata_bits_wdata_10(fringeCommon_io_dram_3_wdata_bits_wdata_10),
    .io_dram_3_wdata_bits_wdata_11(fringeCommon_io_dram_3_wdata_bits_wdata_11),
    .io_dram_3_wdata_bits_wdata_12(fringeCommon_io_dram_3_wdata_bits_wdata_12),
    .io_dram_3_wdata_bits_wdata_13(fringeCommon_io_dram_3_wdata_bits_wdata_13),
    .io_dram_3_wdata_bits_wdata_14(fringeCommon_io_dram_3_wdata_bits_wdata_14),
    .io_dram_3_wdata_bits_wdata_15(fringeCommon_io_dram_3_wdata_bits_wdata_15),
    .io_dram_3_wdata_bits_wstrb_0(fringeCommon_io_dram_3_wdata_bits_wstrb_0),
    .io_dram_3_wdata_bits_wstrb_1(fringeCommon_io_dram_3_wdata_bits_wstrb_1),
    .io_dram_3_wdata_bits_wstrb_2(fringeCommon_io_dram_3_wdata_bits_wstrb_2),
    .io_dram_3_wdata_bits_wstrb_3(fringeCommon_io_dram_3_wdata_bits_wstrb_3),
    .io_dram_3_wdata_bits_wstrb_4(fringeCommon_io_dram_3_wdata_bits_wstrb_4),
    .io_dram_3_wdata_bits_wstrb_5(fringeCommon_io_dram_3_wdata_bits_wstrb_5),
    .io_dram_3_wdata_bits_wstrb_6(fringeCommon_io_dram_3_wdata_bits_wstrb_6),
    .io_dram_3_wdata_bits_wstrb_7(fringeCommon_io_dram_3_wdata_bits_wstrb_7),
    .io_dram_3_wdata_bits_wstrb_8(fringeCommon_io_dram_3_wdata_bits_wstrb_8),
    .io_dram_3_wdata_bits_wstrb_9(fringeCommon_io_dram_3_wdata_bits_wstrb_9),
    .io_dram_3_wdata_bits_wstrb_10(fringeCommon_io_dram_3_wdata_bits_wstrb_10),
    .io_dram_3_wdata_bits_wstrb_11(fringeCommon_io_dram_3_wdata_bits_wstrb_11),
    .io_dram_3_wdata_bits_wstrb_12(fringeCommon_io_dram_3_wdata_bits_wstrb_12),
    .io_dram_3_wdata_bits_wstrb_13(fringeCommon_io_dram_3_wdata_bits_wstrb_13),
    .io_dram_3_wdata_bits_wstrb_14(fringeCommon_io_dram_3_wdata_bits_wstrb_14),
    .io_dram_3_wdata_bits_wstrb_15(fringeCommon_io_dram_3_wdata_bits_wstrb_15),
    .io_dram_3_wdata_bits_wstrb_16(fringeCommon_io_dram_3_wdata_bits_wstrb_16),
    .io_dram_3_wdata_bits_wstrb_17(fringeCommon_io_dram_3_wdata_bits_wstrb_17),
    .io_dram_3_wdata_bits_wstrb_18(fringeCommon_io_dram_3_wdata_bits_wstrb_18),
    .io_dram_3_wdata_bits_wstrb_19(fringeCommon_io_dram_3_wdata_bits_wstrb_19),
    .io_dram_3_wdata_bits_wstrb_20(fringeCommon_io_dram_3_wdata_bits_wstrb_20),
    .io_dram_3_wdata_bits_wstrb_21(fringeCommon_io_dram_3_wdata_bits_wstrb_21),
    .io_dram_3_wdata_bits_wstrb_22(fringeCommon_io_dram_3_wdata_bits_wstrb_22),
    .io_dram_3_wdata_bits_wstrb_23(fringeCommon_io_dram_3_wdata_bits_wstrb_23),
    .io_dram_3_wdata_bits_wstrb_24(fringeCommon_io_dram_3_wdata_bits_wstrb_24),
    .io_dram_3_wdata_bits_wstrb_25(fringeCommon_io_dram_3_wdata_bits_wstrb_25),
    .io_dram_3_wdata_bits_wstrb_26(fringeCommon_io_dram_3_wdata_bits_wstrb_26),
    .io_dram_3_wdata_bits_wstrb_27(fringeCommon_io_dram_3_wdata_bits_wstrb_27),
    .io_dram_3_wdata_bits_wstrb_28(fringeCommon_io_dram_3_wdata_bits_wstrb_28),
    .io_dram_3_wdata_bits_wstrb_29(fringeCommon_io_dram_3_wdata_bits_wstrb_29),
    .io_dram_3_wdata_bits_wstrb_30(fringeCommon_io_dram_3_wdata_bits_wstrb_30),
    .io_dram_3_wdata_bits_wstrb_31(fringeCommon_io_dram_3_wdata_bits_wstrb_31),
    .io_dram_3_wdata_bits_wstrb_32(fringeCommon_io_dram_3_wdata_bits_wstrb_32),
    .io_dram_3_wdata_bits_wstrb_33(fringeCommon_io_dram_3_wdata_bits_wstrb_33),
    .io_dram_3_wdata_bits_wstrb_34(fringeCommon_io_dram_3_wdata_bits_wstrb_34),
    .io_dram_3_wdata_bits_wstrb_35(fringeCommon_io_dram_3_wdata_bits_wstrb_35),
    .io_dram_3_wdata_bits_wstrb_36(fringeCommon_io_dram_3_wdata_bits_wstrb_36),
    .io_dram_3_wdata_bits_wstrb_37(fringeCommon_io_dram_3_wdata_bits_wstrb_37),
    .io_dram_3_wdata_bits_wstrb_38(fringeCommon_io_dram_3_wdata_bits_wstrb_38),
    .io_dram_3_wdata_bits_wstrb_39(fringeCommon_io_dram_3_wdata_bits_wstrb_39),
    .io_dram_3_wdata_bits_wstrb_40(fringeCommon_io_dram_3_wdata_bits_wstrb_40),
    .io_dram_3_wdata_bits_wstrb_41(fringeCommon_io_dram_3_wdata_bits_wstrb_41),
    .io_dram_3_wdata_bits_wstrb_42(fringeCommon_io_dram_3_wdata_bits_wstrb_42),
    .io_dram_3_wdata_bits_wstrb_43(fringeCommon_io_dram_3_wdata_bits_wstrb_43),
    .io_dram_3_wdata_bits_wstrb_44(fringeCommon_io_dram_3_wdata_bits_wstrb_44),
    .io_dram_3_wdata_bits_wstrb_45(fringeCommon_io_dram_3_wdata_bits_wstrb_45),
    .io_dram_3_wdata_bits_wstrb_46(fringeCommon_io_dram_3_wdata_bits_wstrb_46),
    .io_dram_3_wdata_bits_wstrb_47(fringeCommon_io_dram_3_wdata_bits_wstrb_47),
    .io_dram_3_wdata_bits_wstrb_48(fringeCommon_io_dram_3_wdata_bits_wstrb_48),
    .io_dram_3_wdata_bits_wstrb_49(fringeCommon_io_dram_3_wdata_bits_wstrb_49),
    .io_dram_3_wdata_bits_wstrb_50(fringeCommon_io_dram_3_wdata_bits_wstrb_50),
    .io_dram_3_wdata_bits_wstrb_51(fringeCommon_io_dram_3_wdata_bits_wstrb_51),
    .io_dram_3_wdata_bits_wstrb_52(fringeCommon_io_dram_3_wdata_bits_wstrb_52),
    .io_dram_3_wdata_bits_wstrb_53(fringeCommon_io_dram_3_wdata_bits_wstrb_53),
    .io_dram_3_wdata_bits_wstrb_54(fringeCommon_io_dram_3_wdata_bits_wstrb_54),
    .io_dram_3_wdata_bits_wstrb_55(fringeCommon_io_dram_3_wdata_bits_wstrb_55),
    .io_dram_3_wdata_bits_wstrb_56(fringeCommon_io_dram_3_wdata_bits_wstrb_56),
    .io_dram_3_wdata_bits_wstrb_57(fringeCommon_io_dram_3_wdata_bits_wstrb_57),
    .io_dram_3_wdata_bits_wstrb_58(fringeCommon_io_dram_3_wdata_bits_wstrb_58),
    .io_dram_3_wdata_bits_wstrb_59(fringeCommon_io_dram_3_wdata_bits_wstrb_59),
    .io_dram_3_wdata_bits_wstrb_60(fringeCommon_io_dram_3_wdata_bits_wstrb_60),
    .io_dram_3_wdata_bits_wstrb_61(fringeCommon_io_dram_3_wdata_bits_wstrb_61),
    .io_dram_3_wdata_bits_wstrb_62(fringeCommon_io_dram_3_wdata_bits_wstrb_62),
    .io_dram_3_wdata_bits_wstrb_63(fringeCommon_io_dram_3_wdata_bits_wstrb_63),
    .io_dram_3_wdata_bits_wlast(fringeCommon_io_dram_3_wdata_bits_wlast),
    .io_dram_3_rresp_ready(fringeCommon_io_dram_3_rresp_ready),
    .io_dram_3_wresp_ready(fringeCommon_io_dram_3_wresp_ready),
    .io_dram_3_wresp_valid(fringeCommon_io_dram_3_wresp_valid),
    .io_dram_3_wresp_bits_tag(fringeCommon_io_dram_3_wresp_bits_tag),
    .io_heap_0_req_valid(fringeCommon_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(fringeCommon_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(fringeCommon_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(fringeCommon_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(fringeCommon_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(fringeCommon_io_heap_0_resp_bits_sizeAddr)
  );
  AXI4LiteToRFBridge AXI4LiteToRFBridge ( // @[FringeZynq.scala 90:31:@152287.4]
    .clock(AXI4LiteToRFBridge_clock),
    .reset(AXI4LiteToRFBridge_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridge_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridge_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridge_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridge_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridge_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridge_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridge_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridge_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridge_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridge_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridge_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridge_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridge_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridge_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridge_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridge_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridge_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridge_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridge_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridge_io_raddr),
    .io_wen(AXI4LiteToRFBridge_io_wen),
    .io_waddr(AXI4LiteToRFBridge_io_waddr),
    .io_wdata(AXI4LiteToRFBridge_io_wdata),
    .io_rdata(AXI4LiteToRFBridge_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 131:27:@152437.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_1 ( // @[FringeZynq.scala 131:27:@152593.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_1_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_1_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_1_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_1_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_1_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_1_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_1_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_1_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_1_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_1_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_1_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_1_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_1_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_1_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_1_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_1_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_1_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_1_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_1_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_1_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_1_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_1_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_1_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_1_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_1_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_1_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_1_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_1_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_1_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_1_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_1_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_1_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_2 ( // @[FringeZynq.scala 131:27:@152749.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_2_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_2_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_2_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_2_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_2_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_2_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_2_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_2_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_2_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_2_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_2_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_2_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_2_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_2_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_2_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_2_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_2_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_2_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_2_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_2_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_2_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_2_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_2_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_2_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_2_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_2_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_2_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_2_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_2_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_2_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_2_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_2_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_3 ( // @[FringeZynq.scala 131:27:@152905.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_3_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_3_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_3_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_3_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_3_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_3_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_3_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_3_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_3_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_3_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_3_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_3_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_3_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_3_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_3_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_3_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_3_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_3_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_3_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_3_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_3_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_3_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_3_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_3_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_3_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_3_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_3_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_3_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_3_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_3_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_3_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_3_io_M_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 91:28:@152305.4]
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 91:28:@152301.4]
  assign io_S_AXI_WREADY = AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 91:28:@152297.4]
  assign io_S_AXI_RDATA = AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 91:28:@152296.4]
  assign io_S_AXI_RRESP = AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 91:28:@152295.4]
  assign io_S_AXI_RVALID = AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 91:28:@152294.4]
  assign io_S_AXI_BRESP = AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 91:28:@152292.4]
  assign io_S_AXI_BVALID = AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 91:28:@152291.4]
  assign io_M_AXI_0_AWID = MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@152592.4]
  assign io_M_AXI_0_AWADDR = MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@152590.4]
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@152589.4]
  assign io_M_AXI_0_AWVALID = MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@152582.4]
  assign io_M_AXI_0_ARID = MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@152580.4]
  assign io_M_AXI_0_ARADDR = MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@152578.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@152577.4]
  assign io_M_AXI_0_ARVALID = MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@152570.4]
  assign io_M_AXI_0_WDATA = MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@152568.4]
  assign io_M_AXI_0_WSTRB = MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@152567.4]
  assign io_M_AXI_0_WLAST = MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@152566.4]
  assign io_M_AXI_0_WVALID = MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@152565.4]
  assign io_M_AXI_0_RREADY = MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@152557.4]
  assign io_M_AXI_0_BREADY = MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@152552.4]
  assign io_M_AXI_1_AWID = MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@152748.4]
  assign io_M_AXI_1_AWADDR = MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@152746.4]
  assign io_M_AXI_1_AWLEN = MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@152745.4]
  assign io_M_AXI_1_AWVALID = MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@152738.4]
  assign io_M_AXI_1_ARID = MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@152736.4]
  assign io_M_AXI_1_ARADDR = MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@152734.4]
  assign io_M_AXI_1_ARLEN = MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@152733.4]
  assign io_M_AXI_1_ARVALID = MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@152726.4]
  assign io_M_AXI_1_WDATA = MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@152724.4]
  assign io_M_AXI_1_WSTRB = MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@152723.4]
  assign io_M_AXI_1_WLAST = MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@152722.4]
  assign io_M_AXI_1_WVALID = MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@152721.4]
  assign io_M_AXI_1_RREADY = MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@152713.4]
  assign io_M_AXI_1_BREADY = MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@152708.4]
  assign io_M_AXI_2_AWID = MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@152904.4]
  assign io_M_AXI_2_AWADDR = MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@152902.4]
  assign io_M_AXI_2_AWLEN = MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@152901.4]
  assign io_M_AXI_2_AWVALID = MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@152894.4]
  assign io_M_AXI_2_ARID = MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@152892.4]
  assign io_M_AXI_2_ARADDR = MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@152890.4]
  assign io_M_AXI_2_ARLEN = MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@152889.4]
  assign io_M_AXI_2_ARVALID = MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@152882.4]
  assign io_M_AXI_2_WDATA = MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@152880.4]
  assign io_M_AXI_2_WSTRB = MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@152879.4]
  assign io_M_AXI_2_WLAST = MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@152878.4]
  assign io_M_AXI_2_WVALID = MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@152877.4]
  assign io_M_AXI_2_RREADY = MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@152869.4]
  assign io_M_AXI_2_BREADY = MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@152864.4]
  assign io_M_AXI_3_AWID = MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@153060.4]
  assign io_M_AXI_3_AWADDR = MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@153058.4]
  assign io_M_AXI_3_AWLEN = MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@153057.4]
  assign io_M_AXI_3_AWVALID = MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@153050.4]
  assign io_M_AXI_3_ARID = MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@153048.4]
  assign io_M_AXI_3_ARADDR = MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@153046.4]
  assign io_M_AXI_3_ARLEN = MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@153045.4]
  assign io_M_AXI_3_ARVALID = MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@153038.4]
  assign io_M_AXI_3_WDATA = MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@153036.4]
  assign io_M_AXI_3_WSTRB = MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@153035.4]
  assign io_M_AXI_3_WLAST = MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@153034.4]
  assign io_M_AXI_3_WVALID = MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@153033.4]
  assign io_M_AXI_3_RREADY = MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@153025.4]
  assign io_M_AXI_3_BREADY = MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@153020.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 115:13:@152315.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 119:12:@152319.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 121:13:@152320.4]
  assign io_argIns_1 = fringeCommon_io_argIns_1; // @[FringeZynq.scala 121:13:@152321.4]
  assign io_memStreams_stores_0_cmd_ready = fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 126:17:@152408.4]
  assign io_memStreams_stores_0_data_ready = fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 126:17:@152404.4]
  assign io_memStreams_stores_0_wresp_valid = fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 126:17:@152399.4]
  assign io_memStreams_stores_0_wresp_bits = fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 126:17:@152398.4]
  assign io_heap_0_resp_valid = fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 127:11:@152433.4]
  assign io_heap_0_resp_bits_allocDealloc = fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 127:11:@152432.4]
  assign io_heap_0_resp_bits_sizeAddr = fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 127:11:@152431.4]
  assign fringeCommon_clock = clock; // @[:@151382.4]
  assign fringeCommon_reset = reset; // @[:@151383.4 FringeZynq.scala 117:22:@152318.4]
  assign fringeCommon_io_raddr = AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 94:27:@152309.4]
  assign fringeCommon_io_wen = AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 95:27:@152310.4]
  assign fringeCommon_io_waddr = AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 96:27:@152311.4]
  assign fringeCommon_io_wdata = {{32'd0}, AXI4LiteToRFBridge_io_wdata}; // @[FringeZynq.scala 97:27:@152312.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 116:24:@152316.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 122:27:@152323.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 122:27:@152322.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 126:17:@152407.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 126:17:@152406.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 126:17:@152405.4]
  assign fringeCommon_io_memStreams_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 126:17:@152403.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 126:17:@152402.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 126:17:@152401.4]
  assign fringeCommon_io_memStreams_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 126:17:@152400.4]
  assign fringeCommon_io_dram_0_cmd_ready = MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@152551.4]
  assign fringeCommon_io_dram_0_wdata_ready = MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@152544.4]
  assign fringeCommon_io_dram_0_wresp_valid = MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@152441.4]
  assign fringeCommon_io_dram_0_wresp_bits_tag = MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@152440.4]
  assign fringeCommon_io_dram_1_cmd_ready = MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@152707.4]
  assign fringeCommon_io_dram_1_wdata_ready = MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@152700.4]
  assign fringeCommon_io_dram_1_wresp_valid = MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@152597.4]
  assign fringeCommon_io_dram_1_wresp_bits_tag = MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@152596.4]
  assign fringeCommon_io_dram_2_cmd_ready = MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@152863.4]
  assign fringeCommon_io_dram_2_wdata_ready = MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@152856.4]
  assign fringeCommon_io_dram_2_wresp_valid = MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@152753.4]
  assign fringeCommon_io_dram_2_wresp_bits_tag = MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@152752.4]
  assign fringeCommon_io_dram_3_cmd_ready = MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@153019.4]
  assign fringeCommon_io_dram_3_wdata_ready = MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@153012.4]
  assign fringeCommon_io_dram_3_wresp_valid = MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@152909.4]
  assign fringeCommon_io_dram_3_wresp_bits_tag = MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@152908.4]
  assign fringeCommon_io_heap_0_req_valid = io_heap_0_req_valid; // @[FringeZynq.scala 127:11:@152436.4]
  assign fringeCommon_io_heap_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 127:11:@152435.4]
  assign fringeCommon_io_heap_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 127:11:@152434.4]
  assign AXI4LiteToRFBridge_clock = clock; // @[:@152288.4]
  assign AXI4LiteToRFBridge_reset = reset; // @[:@152289.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[FringeZynq.scala 91:28:@152308.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[FringeZynq.scala 91:28:@152307.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[FringeZynq.scala 91:28:@152306.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[FringeZynq.scala 91:28:@152304.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[FringeZynq.scala 91:28:@152303.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[FringeZynq.scala 91:28:@152302.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[FringeZynq.scala 91:28:@152300.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[FringeZynq.scala 91:28:@152299.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[FringeZynq.scala 91:28:@152298.4]
  assign AXI4LiteToRFBridge_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[FringeZynq.scala 91:28:@152293.4]
  assign AXI4LiteToRFBridge_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[FringeZynq.scala 91:28:@152290.4]
  assign AXI4LiteToRFBridge_io_rdata = fringeCommon_io_rdata[31:0]; // @[FringeZynq.scala 98:28:@152313.4]
  assign MAGToAXI4Bridge_io_in_cmd_valid = fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 132:21:@152550.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_addr = fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 132:21:@152549.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_size = fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 132:21:@152548.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_isWr = fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@152546.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_tag = fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 132:21:@152545.4]
  assign MAGToAXI4Bridge_io_in_wdata_valid = fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 132:21:@152543.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@152527.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@152528.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@152529.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@152530.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@152531.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@152532.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@152533.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@152534.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@152535.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@152536.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@152537.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@152538.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@152539.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@152540.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@152541.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@152542.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@152463.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@152464.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@152465.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@152466.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@152467.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@152468.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@152469.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@152470.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@152471.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@152472.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@152473.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@152474.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@152475.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@152476.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@152477.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@152478.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@152479.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@152480.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@152481.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@152482.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@152483.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@152484.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@152485.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@152486.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@152487.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@152488.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@152489.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@152490.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@152491.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@152492.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@152493.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@152494.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@152495.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@152496.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@152497.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@152498.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@152499.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@152500.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@152501.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@152502.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@152503.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@152504.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@152505.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@152506.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@152507.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@152508.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@152509.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@152510.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@152511.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@152512.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@152513.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@152514.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@152515.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@152516.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@152517.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@152518.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@152519.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@152520.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@152521.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@152522.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@152523.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@152524.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@152525.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@152526.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wlast = fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@152462.4]
  assign MAGToAXI4Bridge_io_in_rresp_ready = fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 132:21:@152461.4]
  assign MAGToAXI4Bridge_io_in_wresp_ready = fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 132:21:@152442.4]
  assign MAGToAXI4Bridge_io_M_AXI_AWREADY = io_M_AXI_0_AWREADY; // @[FringeZynq.scala 133:10:@152581.4]
  assign MAGToAXI4Bridge_io_M_AXI_ARREADY = io_M_AXI_0_ARREADY; // @[FringeZynq.scala 133:10:@152569.4]
  assign MAGToAXI4Bridge_io_M_AXI_WREADY = io_M_AXI_0_WREADY; // @[FringeZynq.scala 133:10:@152564.4]
  assign MAGToAXI4Bridge_io_M_AXI_BID = io_M_AXI_0_BID; // @[FringeZynq.scala 133:10:@152556.4]
  assign MAGToAXI4Bridge_io_M_AXI_BVALID = io_M_AXI_0_BVALID; // @[FringeZynq.scala 133:10:@152553.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_valid = fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 132:21:@152706.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_addr = fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 132:21:@152705.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_size = fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 132:21:@152704.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_isWr = fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@152702.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_tag = fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 132:21:@152701.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_valid = fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 132:21:@152699.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@152683.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@152684.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@152685.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@152686.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@152687.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@152688.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@152689.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@152690.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@152691.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@152692.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@152693.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@152694.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@152695.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@152696.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@152697.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@152698.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@152619.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@152620.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@152621.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@152622.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@152623.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@152624.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@152625.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@152626.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@152627.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@152628.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@152629.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@152630.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@152631.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@152632.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@152633.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@152634.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@152635.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@152636.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@152637.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@152638.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@152639.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@152640.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@152641.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@152642.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@152643.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@152644.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@152645.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@152646.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@152647.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@152648.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@152649.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@152650.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@152651.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@152652.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@152653.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@152654.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@152655.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@152656.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@152657.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@152658.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@152659.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@152660.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@152661.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@152662.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@152663.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@152664.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@152665.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@152666.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@152667.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@152668.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@152669.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@152670.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@152671.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@152672.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@152673.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@152674.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@152675.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@152676.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@152677.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@152678.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@152679.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@152680.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@152681.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@152682.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wlast = fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@152618.4]
  assign MAGToAXI4Bridge_1_io_in_rresp_ready = fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 132:21:@152617.4]
  assign MAGToAXI4Bridge_1_io_in_wresp_ready = fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 132:21:@152598.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_AWREADY = io_M_AXI_1_AWREADY; // @[FringeZynq.scala 133:10:@152737.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_ARREADY = io_M_AXI_1_ARREADY; // @[FringeZynq.scala 133:10:@152725.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_WREADY = io_M_AXI_1_WREADY; // @[FringeZynq.scala 133:10:@152720.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BID = io_M_AXI_1_BID; // @[FringeZynq.scala 133:10:@152712.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BVALID = io_M_AXI_1_BVALID; // @[FringeZynq.scala 133:10:@152709.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_valid = fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 132:21:@152862.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_addr = fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 132:21:@152861.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_size = fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 132:21:@152860.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_isWr = fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@152858.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_tag = fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 132:21:@152857.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_valid = fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 132:21:@152855.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@152839.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@152840.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@152841.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@152842.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@152843.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@152844.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@152845.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@152846.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@152847.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@152848.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@152849.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@152850.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@152851.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@152852.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@152853.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@152854.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@152775.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@152776.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@152777.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@152778.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@152779.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@152780.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@152781.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@152782.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@152783.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@152784.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@152785.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@152786.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@152787.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@152788.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@152789.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@152790.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@152791.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@152792.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@152793.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@152794.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@152795.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@152796.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@152797.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@152798.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@152799.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@152800.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@152801.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@152802.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@152803.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@152804.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@152805.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@152806.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@152807.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@152808.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@152809.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@152810.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@152811.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@152812.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@152813.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@152814.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@152815.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@152816.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@152817.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@152818.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@152819.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@152820.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@152821.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@152822.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@152823.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@152824.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@152825.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@152826.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@152827.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@152828.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@152829.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@152830.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@152831.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@152832.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@152833.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@152834.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@152835.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@152836.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@152837.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@152838.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wlast = fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@152774.4]
  assign MAGToAXI4Bridge_2_io_in_rresp_ready = fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 132:21:@152773.4]
  assign MAGToAXI4Bridge_2_io_in_wresp_ready = fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 132:21:@152754.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_AWREADY = io_M_AXI_2_AWREADY; // @[FringeZynq.scala 133:10:@152893.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_ARREADY = io_M_AXI_2_ARREADY; // @[FringeZynq.scala 133:10:@152881.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_WREADY = io_M_AXI_2_WREADY; // @[FringeZynq.scala 133:10:@152876.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BID = io_M_AXI_2_BID; // @[FringeZynq.scala 133:10:@152868.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BVALID = io_M_AXI_2_BVALID; // @[FringeZynq.scala 133:10:@152865.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_valid = fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 132:21:@153018.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_addr = fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 132:21:@153017.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_size = fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 132:21:@153016.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_isWr = fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@153014.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_tag = fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 132:21:@153013.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_valid = fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 132:21:@153011.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@152995.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@152996.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@152997.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@152998.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@152999.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@153000.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@153001.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@153002.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@153003.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@153004.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@153005.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@153006.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@153007.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@153008.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@153009.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@153010.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@152931.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@152932.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@152933.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@152934.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@152935.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@152936.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@152937.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@152938.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@152939.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@152940.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@152941.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@152942.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@152943.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@152944.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@152945.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@152946.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@152947.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@152948.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@152949.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@152950.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@152951.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@152952.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@152953.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@152954.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@152955.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@152956.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@152957.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@152958.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@152959.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@152960.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@152961.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@152962.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@152963.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@152964.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@152965.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@152966.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@152967.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@152968.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@152969.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@152970.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@152971.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@152972.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@152973.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@152974.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@152975.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@152976.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@152977.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@152978.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@152979.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@152980.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@152981.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@152982.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@152983.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@152984.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@152985.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@152986.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@152987.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@152988.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@152989.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@152990.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@152991.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@152992.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@152993.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@152994.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wlast = fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@152930.4]
  assign MAGToAXI4Bridge_3_io_in_rresp_ready = fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 132:21:@152929.4]
  assign MAGToAXI4Bridge_3_io_in_wresp_ready = fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 132:21:@152910.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_AWREADY = io_M_AXI_3_AWREADY; // @[FringeZynq.scala 133:10:@153049.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_ARREADY = io_M_AXI_3_ARREADY; // @[FringeZynq.scala 133:10:@153037.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_WREADY = io_M_AXI_3_WREADY; // @[FringeZynq.scala 133:10:@153032.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BID = io_M_AXI_3_BID; // @[FringeZynq.scala 133:10:@153024.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BVALID = io_M_AXI_3_BVALID; // @[FringeZynq.scala 133:10:@153021.4]
endmodule
module SpatialIP( // @[:@153062.2]
  input          clock, // @[:@153063.4]
  input          reset, // @[:@153064.4]
  input          io_raddr, // @[:@153065.4]
  input          io_wen, // @[:@153065.4]
  input          io_waddr, // @[:@153065.4]
  input          io_wdata, // @[:@153065.4]
  output         io_rdata, // @[:@153065.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@153065.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@153065.4]
  input          io_S_AXI_AWVALID, // @[:@153065.4]
  output         io_S_AXI_AWREADY, // @[:@153065.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@153065.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@153065.4]
  input          io_S_AXI_ARVALID, // @[:@153065.4]
  output         io_S_AXI_ARREADY, // @[:@153065.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@153065.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@153065.4]
  input          io_S_AXI_WVALID, // @[:@153065.4]
  output         io_S_AXI_WREADY, // @[:@153065.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@153065.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@153065.4]
  output         io_S_AXI_RVALID, // @[:@153065.4]
  input          io_S_AXI_RREADY, // @[:@153065.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@153065.4]
  output         io_S_AXI_BVALID, // @[:@153065.4]
  input          io_S_AXI_BREADY, // @[:@153065.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@153065.4]
  output [31:0]  io_M_AXI_0_AWUSER, // @[:@153065.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@153065.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@153065.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@153065.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@153065.4]
  output         io_M_AXI_0_AWLOCK, // @[:@153065.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@153065.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@153065.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@153065.4]
  output         io_M_AXI_0_AWVALID, // @[:@153065.4]
  input          io_M_AXI_0_AWREADY, // @[:@153065.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@153065.4]
  output [31:0]  io_M_AXI_0_ARUSER, // @[:@153065.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@153065.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@153065.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@153065.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@153065.4]
  output         io_M_AXI_0_ARLOCK, // @[:@153065.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@153065.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@153065.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@153065.4]
  output         io_M_AXI_0_ARVALID, // @[:@153065.4]
  input          io_M_AXI_0_ARREADY, // @[:@153065.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@153065.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@153065.4]
  output         io_M_AXI_0_WLAST, // @[:@153065.4]
  output         io_M_AXI_0_WVALID, // @[:@153065.4]
  input          io_M_AXI_0_WREADY, // @[:@153065.4]
  input  [31:0]  io_M_AXI_0_RID, // @[:@153065.4]
  input  [31:0]  io_M_AXI_0_RUSER, // @[:@153065.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@153065.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@153065.4]
  input          io_M_AXI_0_RLAST, // @[:@153065.4]
  input          io_M_AXI_0_RVALID, // @[:@153065.4]
  output         io_M_AXI_0_RREADY, // @[:@153065.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@153065.4]
  input  [31:0]  io_M_AXI_0_BUSER, // @[:@153065.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@153065.4]
  input          io_M_AXI_0_BVALID, // @[:@153065.4]
  output         io_M_AXI_0_BREADY, // @[:@153065.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@153065.4]
  output [31:0]  io_M_AXI_1_AWUSER, // @[:@153065.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@153065.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@153065.4]
  output [2:0]   io_M_AXI_1_AWSIZE, // @[:@153065.4]
  output [1:0]   io_M_AXI_1_AWBURST, // @[:@153065.4]
  output         io_M_AXI_1_AWLOCK, // @[:@153065.4]
  output [3:0]   io_M_AXI_1_AWCACHE, // @[:@153065.4]
  output [2:0]   io_M_AXI_1_AWPROT, // @[:@153065.4]
  output [3:0]   io_M_AXI_1_AWQOS, // @[:@153065.4]
  output         io_M_AXI_1_AWVALID, // @[:@153065.4]
  input          io_M_AXI_1_AWREADY, // @[:@153065.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@153065.4]
  output [31:0]  io_M_AXI_1_ARUSER, // @[:@153065.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@153065.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@153065.4]
  output [2:0]   io_M_AXI_1_ARSIZE, // @[:@153065.4]
  output [1:0]   io_M_AXI_1_ARBURST, // @[:@153065.4]
  output         io_M_AXI_1_ARLOCK, // @[:@153065.4]
  output [3:0]   io_M_AXI_1_ARCACHE, // @[:@153065.4]
  output [2:0]   io_M_AXI_1_ARPROT, // @[:@153065.4]
  output [3:0]   io_M_AXI_1_ARQOS, // @[:@153065.4]
  output         io_M_AXI_1_ARVALID, // @[:@153065.4]
  input          io_M_AXI_1_ARREADY, // @[:@153065.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@153065.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@153065.4]
  output         io_M_AXI_1_WLAST, // @[:@153065.4]
  output         io_M_AXI_1_WVALID, // @[:@153065.4]
  input          io_M_AXI_1_WREADY, // @[:@153065.4]
  input  [31:0]  io_M_AXI_1_RID, // @[:@153065.4]
  input  [31:0]  io_M_AXI_1_RUSER, // @[:@153065.4]
  input  [511:0] io_M_AXI_1_RDATA, // @[:@153065.4]
  input  [1:0]   io_M_AXI_1_RRESP, // @[:@153065.4]
  input          io_M_AXI_1_RLAST, // @[:@153065.4]
  input          io_M_AXI_1_RVALID, // @[:@153065.4]
  output         io_M_AXI_1_RREADY, // @[:@153065.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@153065.4]
  input  [31:0]  io_M_AXI_1_BUSER, // @[:@153065.4]
  input  [1:0]   io_M_AXI_1_BRESP, // @[:@153065.4]
  input          io_M_AXI_1_BVALID, // @[:@153065.4]
  output         io_M_AXI_1_BREADY, // @[:@153065.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@153065.4]
  output [31:0]  io_M_AXI_2_AWUSER, // @[:@153065.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@153065.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@153065.4]
  output [2:0]   io_M_AXI_2_AWSIZE, // @[:@153065.4]
  output [1:0]   io_M_AXI_2_AWBURST, // @[:@153065.4]
  output         io_M_AXI_2_AWLOCK, // @[:@153065.4]
  output [3:0]   io_M_AXI_2_AWCACHE, // @[:@153065.4]
  output [2:0]   io_M_AXI_2_AWPROT, // @[:@153065.4]
  output [3:0]   io_M_AXI_2_AWQOS, // @[:@153065.4]
  output         io_M_AXI_2_AWVALID, // @[:@153065.4]
  input          io_M_AXI_2_AWREADY, // @[:@153065.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@153065.4]
  output [31:0]  io_M_AXI_2_ARUSER, // @[:@153065.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@153065.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@153065.4]
  output [2:0]   io_M_AXI_2_ARSIZE, // @[:@153065.4]
  output [1:0]   io_M_AXI_2_ARBURST, // @[:@153065.4]
  output         io_M_AXI_2_ARLOCK, // @[:@153065.4]
  output [3:0]   io_M_AXI_2_ARCACHE, // @[:@153065.4]
  output [2:0]   io_M_AXI_2_ARPROT, // @[:@153065.4]
  output [3:0]   io_M_AXI_2_ARQOS, // @[:@153065.4]
  output         io_M_AXI_2_ARVALID, // @[:@153065.4]
  input          io_M_AXI_2_ARREADY, // @[:@153065.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@153065.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@153065.4]
  output         io_M_AXI_2_WLAST, // @[:@153065.4]
  output         io_M_AXI_2_WVALID, // @[:@153065.4]
  input          io_M_AXI_2_WREADY, // @[:@153065.4]
  input  [31:0]  io_M_AXI_2_RID, // @[:@153065.4]
  input  [31:0]  io_M_AXI_2_RUSER, // @[:@153065.4]
  input  [511:0] io_M_AXI_2_RDATA, // @[:@153065.4]
  input  [1:0]   io_M_AXI_2_RRESP, // @[:@153065.4]
  input          io_M_AXI_2_RLAST, // @[:@153065.4]
  input          io_M_AXI_2_RVALID, // @[:@153065.4]
  output         io_M_AXI_2_RREADY, // @[:@153065.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@153065.4]
  input  [31:0]  io_M_AXI_2_BUSER, // @[:@153065.4]
  input  [1:0]   io_M_AXI_2_BRESP, // @[:@153065.4]
  input          io_M_AXI_2_BVALID, // @[:@153065.4]
  output         io_M_AXI_2_BREADY, // @[:@153065.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@153065.4]
  output [31:0]  io_M_AXI_3_AWUSER, // @[:@153065.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@153065.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@153065.4]
  output [2:0]   io_M_AXI_3_AWSIZE, // @[:@153065.4]
  output [1:0]   io_M_AXI_3_AWBURST, // @[:@153065.4]
  output         io_M_AXI_3_AWLOCK, // @[:@153065.4]
  output [3:0]   io_M_AXI_3_AWCACHE, // @[:@153065.4]
  output [2:0]   io_M_AXI_3_AWPROT, // @[:@153065.4]
  output [3:0]   io_M_AXI_3_AWQOS, // @[:@153065.4]
  output         io_M_AXI_3_AWVALID, // @[:@153065.4]
  input          io_M_AXI_3_AWREADY, // @[:@153065.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@153065.4]
  output [31:0]  io_M_AXI_3_ARUSER, // @[:@153065.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@153065.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@153065.4]
  output [2:0]   io_M_AXI_3_ARSIZE, // @[:@153065.4]
  output [1:0]   io_M_AXI_3_ARBURST, // @[:@153065.4]
  output         io_M_AXI_3_ARLOCK, // @[:@153065.4]
  output [3:0]   io_M_AXI_3_ARCACHE, // @[:@153065.4]
  output [2:0]   io_M_AXI_3_ARPROT, // @[:@153065.4]
  output [3:0]   io_M_AXI_3_ARQOS, // @[:@153065.4]
  output         io_M_AXI_3_ARVALID, // @[:@153065.4]
  input          io_M_AXI_3_ARREADY, // @[:@153065.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@153065.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@153065.4]
  output         io_M_AXI_3_WLAST, // @[:@153065.4]
  output         io_M_AXI_3_WVALID, // @[:@153065.4]
  input          io_M_AXI_3_WREADY, // @[:@153065.4]
  input  [31:0]  io_M_AXI_3_RID, // @[:@153065.4]
  input  [31:0]  io_M_AXI_3_RUSER, // @[:@153065.4]
  input  [511:0] io_M_AXI_3_RDATA, // @[:@153065.4]
  input  [1:0]   io_M_AXI_3_RRESP, // @[:@153065.4]
  input          io_M_AXI_3_RLAST, // @[:@153065.4]
  input          io_M_AXI_3_RVALID, // @[:@153065.4]
  output         io_M_AXI_3_RREADY, // @[:@153065.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@153065.4]
  input  [31:0]  io_M_AXI_3_BUSER, // @[:@153065.4]
  input  [1:0]   io_M_AXI_3_BRESP, // @[:@153065.4]
  input          io_M_AXI_3_BVALID, // @[:@153065.4]
  output         io_M_AXI_3_BREADY, // @[:@153065.4]
  input          io_TOP_AXI_AWID, // @[:@153065.4]
  input          io_TOP_AXI_AWUSER, // @[:@153065.4]
  input  [31:0]  io_TOP_AXI_AWADDR, // @[:@153065.4]
  input  [7:0]   io_TOP_AXI_AWLEN, // @[:@153065.4]
  input  [2:0]   io_TOP_AXI_AWSIZE, // @[:@153065.4]
  input  [1:0]   io_TOP_AXI_AWBURST, // @[:@153065.4]
  input          io_TOP_AXI_AWLOCK, // @[:@153065.4]
  input  [3:0]   io_TOP_AXI_AWCACHE, // @[:@153065.4]
  input  [2:0]   io_TOP_AXI_AWPROT, // @[:@153065.4]
  input  [3:0]   io_TOP_AXI_AWQOS, // @[:@153065.4]
  input          io_TOP_AXI_AWVALID, // @[:@153065.4]
  input          io_TOP_AXI_AWREADY, // @[:@153065.4]
  input          io_TOP_AXI_ARID, // @[:@153065.4]
  input          io_TOP_AXI_ARUSER, // @[:@153065.4]
  input  [31:0]  io_TOP_AXI_ARADDR, // @[:@153065.4]
  input  [7:0]   io_TOP_AXI_ARLEN, // @[:@153065.4]
  input  [2:0]   io_TOP_AXI_ARSIZE, // @[:@153065.4]
  input  [1:0]   io_TOP_AXI_ARBURST, // @[:@153065.4]
  input          io_TOP_AXI_ARLOCK, // @[:@153065.4]
  input  [3:0]   io_TOP_AXI_ARCACHE, // @[:@153065.4]
  input  [2:0]   io_TOP_AXI_ARPROT, // @[:@153065.4]
  input  [3:0]   io_TOP_AXI_ARQOS, // @[:@153065.4]
  input          io_TOP_AXI_ARVALID, // @[:@153065.4]
  input          io_TOP_AXI_ARREADY, // @[:@153065.4]
  input  [31:0]  io_TOP_AXI_WDATA, // @[:@153065.4]
  input  [63:0]  io_TOP_AXI_WSTRB, // @[:@153065.4]
  input          io_TOP_AXI_WLAST, // @[:@153065.4]
  input          io_TOP_AXI_WVALID, // @[:@153065.4]
  input          io_TOP_AXI_WREADY, // @[:@153065.4]
  input          io_TOP_AXI_RID, // @[:@153065.4]
  input          io_TOP_AXI_RUSER, // @[:@153065.4]
  input  [31:0]  io_TOP_AXI_RDATA, // @[:@153065.4]
  input  [1:0]   io_TOP_AXI_RRESP, // @[:@153065.4]
  input          io_TOP_AXI_RLAST, // @[:@153065.4]
  input          io_TOP_AXI_RVALID, // @[:@153065.4]
  input          io_TOP_AXI_RREADY, // @[:@153065.4]
  input          io_TOP_AXI_BID, // @[:@153065.4]
  input          io_TOP_AXI_BUSER, // @[:@153065.4]
  input  [1:0]   io_TOP_AXI_BRESP, // @[:@153065.4]
  input          io_TOP_AXI_BVALID, // @[:@153065.4]
  input          io_TOP_AXI_BREADY, // @[:@153065.4]
  input          io_DWIDTH_AXI_AWID, // @[:@153065.4]
  input          io_DWIDTH_AXI_AWUSER, // @[:@153065.4]
  input  [31:0]  io_DWIDTH_AXI_AWADDR, // @[:@153065.4]
  input  [7:0]   io_DWIDTH_AXI_AWLEN, // @[:@153065.4]
  input  [2:0]   io_DWIDTH_AXI_AWSIZE, // @[:@153065.4]
  input  [1:0]   io_DWIDTH_AXI_AWBURST, // @[:@153065.4]
  input          io_DWIDTH_AXI_AWLOCK, // @[:@153065.4]
  input  [3:0]   io_DWIDTH_AXI_AWCACHE, // @[:@153065.4]
  input  [2:0]   io_DWIDTH_AXI_AWPROT, // @[:@153065.4]
  input  [3:0]   io_DWIDTH_AXI_AWQOS, // @[:@153065.4]
  input          io_DWIDTH_AXI_AWVALID, // @[:@153065.4]
  input          io_DWIDTH_AXI_AWREADY, // @[:@153065.4]
  input          io_DWIDTH_AXI_ARID, // @[:@153065.4]
  input          io_DWIDTH_AXI_ARUSER, // @[:@153065.4]
  input  [31:0]  io_DWIDTH_AXI_ARADDR, // @[:@153065.4]
  input  [7:0]   io_DWIDTH_AXI_ARLEN, // @[:@153065.4]
  input  [2:0]   io_DWIDTH_AXI_ARSIZE, // @[:@153065.4]
  input  [1:0]   io_DWIDTH_AXI_ARBURST, // @[:@153065.4]
  input          io_DWIDTH_AXI_ARLOCK, // @[:@153065.4]
  input  [3:0]   io_DWIDTH_AXI_ARCACHE, // @[:@153065.4]
  input  [2:0]   io_DWIDTH_AXI_ARPROT, // @[:@153065.4]
  input  [3:0]   io_DWIDTH_AXI_ARQOS, // @[:@153065.4]
  input          io_DWIDTH_AXI_ARVALID, // @[:@153065.4]
  input          io_DWIDTH_AXI_ARREADY, // @[:@153065.4]
  input  [31:0]  io_DWIDTH_AXI_WDATA, // @[:@153065.4]
  input  [63:0]  io_DWIDTH_AXI_WSTRB, // @[:@153065.4]
  input          io_DWIDTH_AXI_WLAST, // @[:@153065.4]
  input          io_DWIDTH_AXI_WVALID, // @[:@153065.4]
  input          io_DWIDTH_AXI_WREADY, // @[:@153065.4]
  input          io_DWIDTH_AXI_RID, // @[:@153065.4]
  input          io_DWIDTH_AXI_RUSER, // @[:@153065.4]
  input  [31:0]  io_DWIDTH_AXI_RDATA, // @[:@153065.4]
  input  [1:0]   io_DWIDTH_AXI_RRESP, // @[:@153065.4]
  input          io_DWIDTH_AXI_RLAST, // @[:@153065.4]
  input          io_DWIDTH_AXI_RVALID, // @[:@153065.4]
  input          io_DWIDTH_AXI_RREADY, // @[:@153065.4]
  input          io_DWIDTH_AXI_BID, // @[:@153065.4]
  input          io_DWIDTH_AXI_BUSER, // @[:@153065.4]
  input  [1:0]   io_DWIDTH_AXI_BRESP, // @[:@153065.4]
  input          io_DWIDTH_AXI_BVALID, // @[:@153065.4]
  input          io_DWIDTH_AXI_BREADY, // @[:@153065.4]
  input          io_PROTOCOL_AXI_AWID, // @[:@153065.4]
  input          io_PROTOCOL_AXI_AWUSER, // @[:@153065.4]
  input  [31:0]  io_PROTOCOL_AXI_AWADDR, // @[:@153065.4]
  input  [7:0]   io_PROTOCOL_AXI_AWLEN, // @[:@153065.4]
  input  [2:0]   io_PROTOCOL_AXI_AWSIZE, // @[:@153065.4]
  input  [1:0]   io_PROTOCOL_AXI_AWBURST, // @[:@153065.4]
  input          io_PROTOCOL_AXI_AWLOCK, // @[:@153065.4]
  input  [3:0]   io_PROTOCOL_AXI_AWCACHE, // @[:@153065.4]
  input  [2:0]   io_PROTOCOL_AXI_AWPROT, // @[:@153065.4]
  input  [3:0]   io_PROTOCOL_AXI_AWQOS, // @[:@153065.4]
  input          io_PROTOCOL_AXI_AWVALID, // @[:@153065.4]
  input          io_PROTOCOL_AXI_AWREADY, // @[:@153065.4]
  input          io_PROTOCOL_AXI_ARID, // @[:@153065.4]
  input          io_PROTOCOL_AXI_ARUSER, // @[:@153065.4]
  input  [31:0]  io_PROTOCOL_AXI_ARADDR, // @[:@153065.4]
  input  [7:0]   io_PROTOCOL_AXI_ARLEN, // @[:@153065.4]
  input  [2:0]   io_PROTOCOL_AXI_ARSIZE, // @[:@153065.4]
  input  [1:0]   io_PROTOCOL_AXI_ARBURST, // @[:@153065.4]
  input          io_PROTOCOL_AXI_ARLOCK, // @[:@153065.4]
  input  [3:0]   io_PROTOCOL_AXI_ARCACHE, // @[:@153065.4]
  input  [2:0]   io_PROTOCOL_AXI_ARPROT, // @[:@153065.4]
  input  [3:0]   io_PROTOCOL_AXI_ARQOS, // @[:@153065.4]
  input          io_PROTOCOL_AXI_ARVALID, // @[:@153065.4]
  input          io_PROTOCOL_AXI_ARREADY, // @[:@153065.4]
  input  [31:0]  io_PROTOCOL_AXI_WDATA, // @[:@153065.4]
  input  [63:0]  io_PROTOCOL_AXI_WSTRB, // @[:@153065.4]
  input          io_PROTOCOL_AXI_WLAST, // @[:@153065.4]
  input          io_PROTOCOL_AXI_WVALID, // @[:@153065.4]
  input          io_PROTOCOL_AXI_WREADY, // @[:@153065.4]
  input          io_PROTOCOL_AXI_RID, // @[:@153065.4]
  input          io_PROTOCOL_AXI_RUSER, // @[:@153065.4]
  input  [31:0]  io_PROTOCOL_AXI_RDATA, // @[:@153065.4]
  input  [1:0]   io_PROTOCOL_AXI_RRESP, // @[:@153065.4]
  input          io_PROTOCOL_AXI_RLAST, // @[:@153065.4]
  input          io_PROTOCOL_AXI_RVALID, // @[:@153065.4]
  input          io_PROTOCOL_AXI_RREADY, // @[:@153065.4]
  input          io_PROTOCOL_AXI_BID, // @[:@153065.4]
  input          io_PROTOCOL_AXI_BUSER, // @[:@153065.4]
  input  [1:0]   io_PROTOCOL_AXI_BRESP, // @[:@153065.4]
  input          io_PROTOCOL_AXI_BVALID, // @[:@153065.4]
  input          io_PROTOCOL_AXI_BREADY, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_AWID, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_AWUSER, // @[:@153065.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_AWADDR, // @[:@153065.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_AWLEN, // @[:@153065.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWSIZE, // @[:@153065.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_AWBURST, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_AWLOCK, // @[:@153065.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWCACHE, // @[:@153065.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWPROT, // @[:@153065.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWQOS, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_AWVALID, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_AWREADY, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_ARID, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_ARUSER, // @[:@153065.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_ARADDR, // @[:@153065.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_ARLEN, // @[:@153065.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARSIZE, // @[:@153065.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_ARBURST, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_ARLOCK, // @[:@153065.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARCACHE, // @[:@153065.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARPROT, // @[:@153065.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARQOS, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_ARVALID, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_ARREADY, // @[:@153065.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_WDATA, // @[:@153065.4]
  input  [63:0]  io_CLOCKCONVERT_AXI_WSTRB, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_WLAST, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_WVALID, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_WREADY, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_RID, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_RUSER, // @[:@153065.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_RDATA, // @[:@153065.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_RRESP, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_RLAST, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_RVALID, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_RREADY, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_BID, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_BUSER, // @[:@153065.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_BRESP, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_BVALID, // @[:@153065.4]
  input          io_CLOCKCONVERT_AXI_BREADY // @[:@153065.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@153067.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@153067.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@153067.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@153067.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@153067.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@153067.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@153067.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@153067.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@153067.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@153067.4]
  wire  FringeZynq_clock; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_reset; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_S_AXI_AWADDR; // @[Zynq.scala 18:24:@153209.4]
  wire [2:0] FringeZynq_io_S_AXI_AWPROT; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_S_AXI_AWVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_S_AXI_ARADDR; // @[Zynq.scala 18:24:@153209.4]
  wire [2:0] FringeZynq_io_S_AXI_ARPROT; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_S_AXI_ARVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_S_AXI_WDATA; // @[Zynq.scala 18:24:@153209.4]
  wire [3:0] FringeZynq_io_S_AXI_WSTRB; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_S_AXI_WVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 18:24:@153209.4]
  wire [1:0] FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_S_AXI_RREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [1:0] FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_S_AXI_BREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 18:24:@153209.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_0_AWREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 18:24:@153209.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_0_ARREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [511:0] FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 18:24:@153209.4]
  wire [63:0] FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_0_WREADY; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_0_BID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_0_BVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 18:24:@153209.4]
  wire [7:0] FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_1_AWREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 18:24:@153209.4]
  wire [7:0] FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_1_ARREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [511:0] FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 18:24:@153209.4]
  wire [63:0] FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_1_WREADY; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_1_BID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_1_BVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 18:24:@153209.4]
  wire [7:0] FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_2_AWREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 18:24:@153209.4]
  wire [7:0] FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_2_ARREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [511:0] FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 18:24:@153209.4]
  wire [63:0] FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_2_WREADY; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_2_BID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_2_BVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 18:24:@153209.4]
  wire [7:0] FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_3_AWREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 18:24:@153209.4]
  wire [7:0] FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_3_ARREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [511:0] FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 18:24:@153209.4]
  wire [63:0] FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_3_WREADY; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_M_AXI_3_BID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_3_BVALID; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_enable; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_done; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_reset; // @[Zynq.scala 18:24:@153209.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[Zynq.scala 18:24:@153209.4]
  wire [63:0] FringeZynq_io_argIns_1; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[Zynq.scala 18:24:@153209.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 18:24:@153209.4]
  wire [63:0] FringeZynq_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_memStreams_stores_0_data_valid; // @[Zynq.scala 18:24:@153209.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_heap_0_req_valid; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 18:24:@153209.4]
  wire [63:0] FringeZynq_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 18:24:@153209.4]
  wire  FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 18:24:@153209.4]
  wire [63:0] FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 18:24:@153209.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@153067.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  FringeZynq FringeZynq ( // @[Zynq.scala 18:24:@153209.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWID(FringeZynq_io_M_AXI_0_AWID),
    .io_M_AXI_0_AWADDR(FringeZynq_io_M_AXI_0_AWADDR),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_AWVALID(FringeZynq_io_M_AXI_0_AWVALID),
    .io_M_AXI_0_AWREADY(FringeZynq_io_M_AXI_0_AWREADY),
    .io_M_AXI_0_ARID(FringeZynq_io_M_AXI_0_ARID),
    .io_M_AXI_0_ARADDR(FringeZynq_io_M_AXI_0_ARADDR),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_M_AXI_0_ARVALID(FringeZynq_io_M_AXI_0_ARVALID),
    .io_M_AXI_0_ARREADY(FringeZynq_io_M_AXI_0_ARREADY),
    .io_M_AXI_0_WDATA(FringeZynq_io_M_AXI_0_WDATA),
    .io_M_AXI_0_WSTRB(FringeZynq_io_M_AXI_0_WSTRB),
    .io_M_AXI_0_WLAST(FringeZynq_io_M_AXI_0_WLAST),
    .io_M_AXI_0_WVALID(FringeZynq_io_M_AXI_0_WVALID),
    .io_M_AXI_0_WREADY(FringeZynq_io_M_AXI_0_WREADY),
    .io_M_AXI_0_RREADY(FringeZynq_io_M_AXI_0_RREADY),
    .io_M_AXI_0_BID(FringeZynq_io_M_AXI_0_BID),
    .io_M_AXI_0_BVALID(FringeZynq_io_M_AXI_0_BVALID),
    .io_M_AXI_0_BREADY(FringeZynq_io_M_AXI_0_BREADY),
    .io_M_AXI_1_AWID(FringeZynq_io_M_AXI_1_AWID),
    .io_M_AXI_1_AWADDR(FringeZynq_io_M_AXI_1_AWADDR),
    .io_M_AXI_1_AWLEN(FringeZynq_io_M_AXI_1_AWLEN),
    .io_M_AXI_1_AWVALID(FringeZynq_io_M_AXI_1_AWVALID),
    .io_M_AXI_1_AWREADY(FringeZynq_io_M_AXI_1_AWREADY),
    .io_M_AXI_1_ARID(FringeZynq_io_M_AXI_1_ARID),
    .io_M_AXI_1_ARADDR(FringeZynq_io_M_AXI_1_ARADDR),
    .io_M_AXI_1_ARLEN(FringeZynq_io_M_AXI_1_ARLEN),
    .io_M_AXI_1_ARVALID(FringeZynq_io_M_AXI_1_ARVALID),
    .io_M_AXI_1_ARREADY(FringeZynq_io_M_AXI_1_ARREADY),
    .io_M_AXI_1_WDATA(FringeZynq_io_M_AXI_1_WDATA),
    .io_M_AXI_1_WSTRB(FringeZynq_io_M_AXI_1_WSTRB),
    .io_M_AXI_1_WLAST(FringeZynq_io_M_AXI_1_WLAST),
    .io_M_AXI_1_WVALID(FringeZynq_io_M_AXI_1_WVALID),
    .io_M_AXI_1_WREADY(FringeZynq_io_M_AXI_1_WREADY),
    .io_M_AXI_1_RREADY(FringeZynq_io_M_AXI_1_RREADY),
    .io_M_AXI_1_BID(FringeZynq_io_M_AXI_1_BID),
    .io_M_AXI_1_BVALID(FringeZynq_io_M_AXI_1_BVALID),
    .io_M_AXI_1_BREADY(FringeZynq_io_M_AXI_1_BREADY),
    .io_M_AXI_2_AWID(FringeZynq_io_M_AXI_2_AWID),
    .io_M_AXI_2_AWADDR(FringeZynq_io_M_AXI_2_AWADDR),
    .io_M_AXI_2_AWLEN(FringeZynq_io_M_AXI_2_AWLEN),
    .io_M_AXI_2_AWVALID(FringeZynq_io_M_AXI_2_AWVALID),
    .io_M_AXI_2_AWREADY(FringeZynq_io_M_AXI_2_AWREADY),
    .io_M_AXI_2_ARID(FringeZynq_io_M_AXI_2_ARID),
    .io_M_AXI_2_ARADDR(FringeZynq_io_M_AXI_2_ARADDR),
    .io_M_AXI_2_ARLEN(FringeZynq_io_M_AXI_2_ARLEN),
    .io_M_AXI_2_ARVALID(FringeZynq_io_M_AXI_2_ARVALID),
    .io_M_AXI_2_ARREADY(FringeZynq_io_M_AXI_2_ARREADY),
    .io_M_AXI_2_WDATA(FringeZynq_io_M_AXI_2_WDATA),
    .io_M_AXI_2_WSTRB(FringeZynq_io_M_AXI_2_WSTRB),
    .io_M_AXI_2_WLAST(FringeZynq_io_M_AXI_2_WLAST),
    .io_M_AXI_2_WVALID(FringeZynq_io_M_AXI_2_WVALID),
    .io_M_AXI_2_WREADY(FringeZynq_io_M_AXI_2_WREADY),
    .io_M_AXI_2_RREADY(FringeZynq_io_M_AXI_2_RREADY),
    .io_M_AXI_2_BID(FringeZynq_io_M_AXI_2_BID),
    .io_M_AXI_2_BVALID(FringeZynq_io_M_AXI_2_BVALID),
    .io_M_AXI_2_BREADY(FringeZynq_io_M_AXI_2_BREADY),
    .io_M_AXI_3_AWID(FringeZynq_io_M_AXI_3_AWID),
    .io_M_AXI_3_AWADDR(FringeZynq_io_M_AXI_3_AWADDR),
    .io_M_AXI_3_AWLEN(FringeZynq_io_M_AXI_3_AWLEN),
    .io_M_AXI_3_AWVALID(FringeZynq_io_M_AXI_3_AWVALID),
    .io_M_AXI_3_AWREADY(FringeZynq_io_M_AXI_3_AWREADY),
    .io_M_AXI_3_ARID(FringeZynq_io_M_AXI_3_ARID),
    .io_M_AXI_3_ARADDR(FringeZynq_io_M_AXI_3_ARADDR),
    .io_M_AXI_3_ARLEN(FringeZynq_io_M_AXI_3_ARLEN),
    .io_M_AXI_3_ARVALID(FringeZynq_io_M_AXI_3_ARVALID),
    .io_M_AXI_3_ARREADY(FringeZynq_io_M_AXI_3_ARREADY),
    .io_M_AXI_3_WDATA(FringeZynq_io_M_AXI_3_WDATA),
    .io_M_AXI_3_WSTRB(FringeZynq_io_M_AXI_3_WSTRB),
    .io_M_AXI_3_WLAST(FringeZynq_io_M_AXI_3_WLAST),
    .io_M_AXI_3_WVALID(FringeZynq_io_M_AXI_3_WVALID),
    .io_M_AXI_3_WREADY(FringeZynq_io_M_AXI_3_WREADY),
    .io_M_AXI_3_RREADY(FringeZynq_io_M_AXI_3_RREADY),
    .io_M_AXI_3_BID(FringeZynq_io_M_AXI_3_BID),
    .io_M_AXI_3_BVALID(FringeZynq_io_M_AXI_3_BVALID),
    .io_M_AXI_3_BREADY(FringeZynq_io_M_AXI_3_BREADY),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argIns_1(FringeZynq_io_argIns_1),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(FringeZynq_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(FringeZynq_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(FringeZynq_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(FringeZynq_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(FringeZynq_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(FringeZynq_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(FringeZynq_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(FringeZynq_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(FringeZynq_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(FringeZynq_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(FringeZynq_io_memStreams_stores_0_wresp_bits),
    .io_heap_0_req_valid(FringeZynq_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(FringeZynq_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(FringeZynq_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(FringeZynq_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(FringeZynq_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(FringeZynq_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 21:21:@153227.4]
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 21:21:@153223.4]
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 21:21:@153219.4]
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 21:21:@153218.4]
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 21:21:@153217.4]
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 21:21:@153216.4]
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 21:21:@153214.4]
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 21:21:@153213.4]
  assign io_M_AXI_0_AWID = FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 24:14:@153271.4]
  assign io_M_AXI_0_AWUSER = 32'h0; // @[Zynq.scala 24:14:@153270.4]
  assign io_M_AXI_0_AWADDR = FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 24:14:@153269.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 24:14:@153268.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@153267.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[Zynq.scala 24:14:@153266.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@153265.4]
  assign io_M_AXI_0_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@153264.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[Zynq.scala 24:14:@153263.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[Zynq.scala 24:14:@153262.4]
  assign io_M_AXI_0_AWVALID = FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 24:14:@153261.4]
  assign io_M_AXI_0_ARID = FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 24:14:@153259.4]
  assign io_M_AXI_0_ARUSER = 32'h0; // @[Zynq.scala 24:14:@153258.4]
  assign io_M_AXI_0_ARADDR = FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 24:14:@153257.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 24:14:@153256.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@153255.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[Zynq.scala 24:14:@153254.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@153253.4]
  assign io_M_AXI_0_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@153252.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[Zynq.scala 24:14:@153251.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[Zynq.scala 24:14:@153250.4]
  assign io_M_AXI_0_ARVALID = FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 24:14:@153249.4]
  assign io_M_AXI_0_WDATA = FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 24:14:@153247.4]
  assign io_M_AXI_0_WSTRB = FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 24:14:@153246.4]
  assign io_M_AXI_0_WLAST = FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 24:14:@153245.4]
  assign io_M_AXI_0_WVALID = FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 24:14:@153244.4]
  assign io_M_AXI_0_RREADY = FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 24:14:@153236.4]
  assign io_M_AXI_0_BREADY = FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 24:14:@153231.4]
  assign io_M_AXI_1_AWID = FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 24:14:@153312.4]
  assign io_M_AXI_1_AWUSER = 32'h0; // @[Zynq.scala 24:14:@153311.4]
  assign io_M_AXI_1_AWADDR = FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 24:14:@153310.4]
  assign io_M_AXI_1_AWLEN = FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 24:14:@153309.4]
  assign io_M_AXI_1_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@153308.4]
  assign io_M_AXI_1_AWBURST = 2'h1; // @[Zynq.scala 24:14:@153307.4]
  assign io_M_AXI_1_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@153306.4]
  assign io_M_AXI_1_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@153305.4]
  assign io_M_AXI_1_AWPROT = 3'h0; // @[Zynq.scala 24:14:@153304.4]
  assign io_M_AXI_1_AWQOS = 4'h0; // @[Zynq.scala 24:14:@153303.4]
  assign io_M_AXI_1_AWVALID = FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 24:14:@153302.4]
  assign io_M_AXI_1_ARID = FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 24:14:@153300.4]
  assign io_M_AXI_1_ARUSER = 32'h0; // @[Zynq.scala 24:14:@153299.4]
  assign io_M_AXI_1_ARADDR = FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 24:14:@153298.4]
  assign io_M_AXI_1_ARLEN = FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 24:14:@153297.4]
  assign io_M_AXI_1_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@153296.4]
  assign io_M_AXI_1_ARBURST = 2'h1; // @[Zynq.scala 24:14:@153295.4]
  assign io_M_AXI_1_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@153294.4]
  assign io_M_AXI_1_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@153293.4]
  assign io_M_AXI_1_ARPROT = 3'h0; // @[Zynq.scala 24:14:@153292.4]
  assign io_M_AXI_1_ARQOS = 4'h0; // @[Zynq.scala 24:14:@153291.4]
  assign io_M_AXI_1_ARVALID = FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 24:14:@153290.4]
  assign io_M_AXI_1_WDATA = FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 24:14:@153288.4]
  assign io_M_AXI_1_WSTRB = FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 24:14:@153287.4]
  assign io_M_AXI_1_WLAST = FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 24:14:@153286.4]
  assign io_M_AXI_1_WVALID = FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 24:14:@153285.4]
  assign io_M_AXI_1_RREADY = FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 24:14:@153277.4]
  assign io_M_AXI_1_BREADY = FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 24:14:@153272.4]
  assign io_M_AXI_2_AWID = FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 24:14:@153353.4]
  assign io_M_AXI_2_AWUSER = 32'h0; // @[Zynq.scala 24:14:@153352.4]
  assign io_M_AXI_2_AWADDR = FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 24:14:@153351.4]
  assign io_M_AXI_2_AWLEN = FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 24:14:@153350.4]
  assign io_M_AXI_2_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@153349.4]
  assign io_M_AXI_2_AWBURST = 2'h1; // @[Zynq.scala 24:14:@153348.4]
  assign io_M_AXI_2_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@153347.4]
  assign io_M_AXI_2_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@153346.4]
  assign io_M_AXI_2_AWPROT = 3'h0; // @[Zynq.scala 24:14:@153345.4]
  assign io_M_AXI_2_AWQOS = 4'h0; // @[Zynq.scala 24:14:@153344.4]
  assign io_M_AXI_2_AWVALID = FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 24:14:@153343.4]
  assign io_M_AXI_2_ARID = FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 24:14:@153341.4]
  assign io_M_AXI_2_ARUSER = 32'h0; // @[Zynq.scala 24:14:@153340.4]
  assign io_M_AXI_2_ARADDR = FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 24:14:@153339.4]
  assign io_M_AXI_2_ARLEN = FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 24:14:@153338.4]
  assign io_M_AXI_2_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@153337.4]
  assign io_M_AXI_2_ARBURST = 2'h1; // @[Zynq.scala 24:14:@153336.4]
  assign io_M_AXI_2_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@153335.4]
  assign io_M_AXI_2_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@153334.4]
  assign io_M_AXI_2_ARPROT = 3'h0; // @[Zynq.scala 24:14:@153333.4]
  assign io_M_AXI_2_ARQOS = 4'h0; // @[Zynq.scala 24:14:@153332.4]
  assign io_M_AXI_2_ARVALID = FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 24:14:@153331.4]
  assign io_M_AXI_2_WDATA = FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 24:14:@153329.4]
  assign io_M_AXI_2_WSTRB = FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 24:14:@153328.4]
  assign io_M_AXI_2_WLAST = FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 24:14:@153327.4]
  assign io_M_AXI_2_WVALID = FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 24:14:@153326.4]
  assign io_M_AXI_2_RREADY = FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 24:14:@153318.4]
  assign io_M_AXI_2_BREADY = FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 24:14:@153313.4]
  assign io_M_AXI_3_AWID = FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 24:14:@153394.4]
  assign io_M_AXI_3_AWUSER = 32'h0; // @[Zynq.scala 24:14:@153393.4]
  assign io_M_AXI_3_AWADDR = FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 24:14:@153392.4]
  assign io_M_AXI_3_AWLEN = FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 24:14:@153391.4]
  assign io_M_AXI_3_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@153390.4]
  assign io_M_AXI_3_AWBURST = 2'h1; // @[Zynq.scala 24:14:@153389.4]
  assign io_M_AXI_3_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@153388.4]
  assign io_M_AXI_3_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@153387.4]
  assign io_M_AXI_3_AWPROT = 3'h0; // @[Zynq.scala 24:14:@153386.4]
  assign io_M_AXI_3_AWQOS = 4'h0; // @[Zynq.scala 24:14:@153385.4]
  assign io_M_AXI_3_AWVALID = FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 24:14:@153384.4]
  assign io_M_AXI_3_ARID = FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 24:14:@153382.4]
  assign io_M_AXI_3_ARUSER = 32'h0; // @[Zynq.scala 24:14:@153381.4]
  assign io_M_AXI_3_ARADDR = FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 24:14:@153380.4]
  assign io_M_AXI_3_ARLEN = FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 24:14:@153379.4]
  assign io_M_AXI_3_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@153378.4]
  assign io_M_AXI_3_ARBURST = 2'h1; // @[Zynq.scala 24:14:@153377.4]
  assign io_M_AXI_3_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@153376.4]
  assign io_M_AXI_3_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@153375.4]
  assign io_M_AXI_3_ARPROT = 3'h0; // @[Zynq.scala 24:14:@153374.4]
  assign io_M_AXI_3_ARQOS = 4'h0; // @[Zynq.scala 24:14:@153373.4]
  assign io_M_AXI_3_ARVALID = FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 24:14:@153372.4]
  assign io_M_AXI_3_WDATA = FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 24:14:@153370.4]
  assign io_M_AXI_3_WSTRB = FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 24:14:@153369.4]
  assign io_M_AXI_3_WLAST = FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 24:14:@153368.4]
  assign io_M_AXI_3_WVALID = FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 24:14:@153367.4]
  assign io_M_AXI_3_RREADY = FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 24:14:@153359.4]
  assign io_M_AXI_3_BREADY = FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 24:14:@153354.4]
  assign accel_clock = clock; // @[:@153068.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@153069.4 Zynq.scala 54:17:@153683.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[Zynq.scala 51:21:@153678.4]
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@153671.4]
  assign accel_io_memStreams_loads_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@153666.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0; // @[Zynq.scala 49:26:@153650.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0; // @[Zynq.scala 49:26:@153651.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0; // @[Zynq.scala 49:26:@153652.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0; // @[Zynq.scala 49:26:@153653.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0; // @[Zynq.scala 49:26:@153654.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0; // @[Zynq.scala 49:26:@153655.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0; // @[Zynq.scala 49:26:@153656.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0; // @[Zynq.scala 49:26:@153657.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0; // @[Zynq.scala 49:26:@153658.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0; // @[Zynq.scala 49:26:@153659.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0; // @[Zynq.scala 49:26:@153660.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0; // @[Zynq.scala 49:26:@153661.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0; // @[Zynq.scala 49:26:@153662.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0; // @[Zynq.scala 49:26:@153663.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0; // @[Zynq.scala 49:26:@153664.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0; // @[Zynq.scala 49:26:@153665.4]
  assign accel_io_memStreams_stores_0_cmd_ready = FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 49:26:@153649.4]
  assign accel_io_memStreams_stores_0_data_ready = FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 49:26:@153645.4]
  assign accel_io_memStreams_stores_0_wresp_valid = FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 49:26:@153640.4]
  assign accel_io_memStreams_stores_0_wresp_bits = FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 49:26:@153639.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@153638.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@153619.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0; // @[Zynq.scala 49:26:@153603.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0; // @[Zynq.scala 49:26:@153604.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0; // @[Zynq.scala 49:26:@153605.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0; // @[Zynq.scala 49:26:@153606.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0; // @[Zynq.scala 49:26:@153607.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0; // @[Zynq.scala 49:26:@153608.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0; // @[Zynq.scala 49:26:@153609.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0; // @[Zynq.scala 49:26:@153610.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0; // @[Zynq.scala 49:26:@153611.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0; // @[Zynq.scala 49:26:@153612.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0; // @[Zynq.scala 49:26:@153613.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0; // @[Zynq.scala 49:26:@153614.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0; // @[Zynq.scala 49:26:@153615.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0; // @[Zynq.scala 49:26:@153616.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0; // @[Zynq.scala 49:26:@153617.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0; // @[Zynq.scala 49:26:@153618.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@153602.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[Zynq.scala 49:26:@153567.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[Zynq.scala 49:26:@153566.4]
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 50:20:@153674.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 50:20:@153673.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 50:20:@153672.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[Zynq.scala 34:21:@153560.4]
  assign accel_io_argIns_1 = FringeZynq_io_argIns_1; // @[Zynq.scala 34:21:@153561.4]
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0; // @[Zynq.scala 40:24:@153564.4]
  assign FringeZynq_clock = clock; // @[:@153210.4]
  assign FringeZynq_reset = reset == 1'h0; // @[:@153211.4 Zynq.scala 53:18:@153682.4]
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[Zynq.scala 21:21:@153230.4]
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[Zynq.scala 21:21:@153229.4]
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[Zynq.scala 21:21:@153228.4]
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[Zynq.scala 21:21:@153226.4]
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[Zynq.scala 21:21:@153225.4]
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[Zynq.scala 21:21:@153224.4]
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[Zynq.scala 21:21:@153222.4]
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[Zynq.scala 21:21:@153221.4]
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[Zynq.scala 21:21:@153220.4]
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[Zynq.scala 21:21:@153215.4]
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[Zynq.scala 21:21:@153212.4]
  assign FringeZynq_io_M_AXI_0_AWREADY = io_M_AXI_0_AWREADY; // @[Zynq.scala 24:14:@153260.4]
  assign FringeZynq_io_M_AXI_0_ARREADY = io_M_AXI_0_ARREADY; // @[Zynq.scala 24:14:@153248.4]
  assign FringeZynq_io_M_AXI_0_WREADY = io_M_AXI_0_WREADY; // @[Zynq.scala 24:14:@153243.4]
  assign FringeZynq_io_M_AXI_0_BID = io_M_AXI_0_BID; // @[Zynq.scala 24:14:@153235.4]
  assign FringeZynq_io_M_AXI_0_BVALID = io_M_AXI_0_BVALID; // @[Zynq.scala 24:14:@153232.4]
  assign FringeZynq_io_M_AXI_1_AWREADY = io_M_AXI_1_AWREADY; // @[Zynq.scala 24:14:@153301.4]
  assign FringeZynq_io_M_AXI_1_ARREADY = io_M_AXI_1_ARREADY; // @[Zynq.scala 24:14:@153289.4]
  assign FringeZynq_io_M_AXI_1_WREADY = io_M_AXI_1_WREADY; // @[Zynq.scala 24:14:@153284.4]
  assign FringeZynq_io_M_AXI_1_BID = io_M_AXI_1_BID; // @[Zynq.scala 24:14:@153276.4]
  assign FringeZynq_io_M_AXI_1_BVALID = io_M_AXI_1_BVALID; // @[Zynq.scala 24:14:@153273.4]
  assign FringeZynq_io_M_AXI_2_AWREADY = io_M_AXI_2_AWREADY; // @[Zynq.scala 24:14:@153342.4]
  assign FringeZynq_io_M_AXI_2_ARREADY = io_M_AXI_2_ARREADY; // @[Zynq.scala 24:14:@153330.4]
  assign FringeZynq_io_M_AXI_2_WREADY = io_M_AXI_2_WREADY; // @[Zynq.scala 24:14:@153325.4]
  assign FringeZynq_io_M_AXI_2_BID = io_M_AXI_2_BID; // @[Zynq.scala 24:14:@153317.4]
  assign FringeZynq_io_M_AXI_2_BVALID = io_M_AXI_2_BVALID; // @[Zynq.scala 24:14:@153314.4]
  assign FringeZynq_io_M_AXI_3_AWREADY = io_M_AXI_3_AWREADY; // @[Zynq.scala 24:14:@153383.4]
  assign FringeZynq_io_M_AXI_3_ARREADY = io_M_AXI_3_ARREADY; // @[Zynq.scala 24:14:@153371.4]
  assign FringeZynq_io_M_AXI_3_WREADY = io_M_AXI_3_WREADY; // @[Zynq.scala 24:14:@153366.4]
  assign FringeZynq_io_M_AXI_3_BID = io_M_AXI_3_BID; // @[Zynq.scala 24:14:@153358.4]
  assign FringeZynq_io_M_AXI_3_BVALID = io_M_AXI_3_BVALID; // @[Zynq.scala 24:14:@153355.4]
  assign FringeZynq_io_done = accel_io_done; // @[Zynq.scala 52:20:@153679.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[Zynq.scala 37:26:@153563.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[Zynq.scala 36:25:@153562.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_valid = accel_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 49:26:@153648.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_addr = accel_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 49:26:@153647.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_size = accel_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 49:26:@153646.4]
  assign FringeZynq_io_memStreams_stores_0_data_valid = accel_io_memStreams_stores_0_data_valid; // @[Zynq.scala 49:26:@153644.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wdata_0 = accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 49:26:@153643.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wstrb = accel_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 49:26:@153642.4]
  assign FringeZynq_io_memStreams_stores_0_wresp_ready = accel_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 49:26:@153641.4]
  assign FringeZynq_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[Zynq.scala 50:20:@153677.4]
  assign FringeZynq_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 50:20:@153676.4]
  assign FringeZynq_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 50:20:@153675.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
module SRAMVerilogDualRead
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr0,
    input [AWIDTH-1:0] raddr1,
    input [AWIDTH-1:0] waddr,
    input raddrEn0,
    input raddrEn1,
    input waddrEn,
    input wen,
    input backpressure0,
    input backpressure1,
    input [DWIDTH-1:0] wdata,
    output reg [DWIDTH-1:0] rdata0,
    output reg [DWIDTH-1:0] rdata1
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk)
    begin
            if (wen)
            begin
                mem[waddr] <= wdata;
            end
            if (backpressure0) rdata0 <= mem[raddr0];
    end


    always @(posedge clk)
    begin
        if (backpressure1) rdata1 <= mem[raddr1];
    end
endmodule




